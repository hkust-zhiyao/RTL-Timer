module b17(clock, reset, hold, na, bs16, wr, dc, mio, ast1, ast2, ready1, ready2, datai, datao, address1, address2);
  wire reset_n_DEFINE;
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire [1:0] _00402_;
  wire _00403_;
  wire [1:0] _00404_;
  wire _00405_;
  wire [1:0] _00406_;
  wire _00407_;
  wire [1:0] _00408_;
  wire _00409_;
  wire [1:0] _00410_;
  wire _00411_;
  wire [1:0] _00412_;
  wire _00413_;
  wire [1:0] _00414_;
  wire _00415_;
  wire [1:0] _00416_;
  wire _00417_;
  wire [1:0] _00418_;
  wire _00419_;
  wire [1:0] _00420_;
  wire _00421_;
  wire [1:0] _00422_;
  wire _00423_;
  wire [1:0] _00424_;
  wire _00425_;
  wire [1:0] _00426_;
  wire _00427_;
  wire [1:0] _00428_;
  wire _00429_;
  wire [1:0] _00430_;
  wire _00431_;
  wire [1:0] _00432_;
  wire _00433_;
  wire [1:0] _00434_;
  wire _00435_;
  wire [1:0] _00436_;
  wire _00437_;
  wire [1:0] _00438_;
  wire _00439_;
  wire [1:0] _00440_;
  wire _00441_;
  wire [1:0] _00442_;
  wire _00443_;
  wire [1:0] _00444_;
  wire _00445_;
  wire [1:0] _00446_;
  wire _00447_;
  wire [1:0] _00448_;
  wire _00449_;
  wire [1:0] _00450_;
  wire _00451_;
  wire [1:0] _00452_;
  wire _00453_;
  wire [1:0] _00454_;
  wire _00455_;
  wire [1:0] _00456_;
  wire _00457_;
  wire [1:0] _00458_;
  wire _00459_;
  wire [1:0] _00460_;
  wire _00461_;
  wire [1:0] _00462_;
  wire _00463_;
  wire [1:0] _00464_;
  wire _00465_;
  wire [1:0] _00466_;
  wire _00467_;
  wire [1:0] _00468_;
  wire [1:0] _00469_;
  wire [1:0] _00470_;
  wire [2:0] _00471_;
  wire [1:0] _00472_;
  wire [2:0] _00473_;
  wire [1:0] _00474_;
  wire [2:0] _00475_;
  wire [1:0] _00476_;
  wire [2:0] _00477_;
  wire [1:0] _00478_;
  wire [2:0] _00479_;
  wire [1:0] _00480_;
  wire [2:0] _00481_;
  wire [1:0] _00482_;
  wire [1:0] _00483_;
  wire [1:0] _00484_;
  wire _00485_;
  wire _00486_;
  wire [1:0] _00487_;
  wire [1:0] _00488_;
  wire [1:0] _00489_;
  wire [1:0] _00490_;
  wire [1:0] _00491_;
  wire [1:0] _00492_;
  wire [1:0] _00493_;
  wire [1:0] _00494_;
  wire [1:0] _00495_;
  wire [1:0] _00496_;
  wire [1:0] _00497_;
  wire [1:0] _00498_;
  wire [1:0] _00499_;
  wire [1:0] _00500_;
  wire [1:0] _00501_;
  wire [1:0] _00502_;
  wire [1:0] _00503_;
  wire [1:0] _00504_;
  wire [1:0] _00505_;
  wire [1:0] _00506_;
  wire [1:0] _00507_;
  wire [1:0] _00508_;
  wire [1:0] _00509_;
  wire [1:0] _00510_;
  wire [1:0] _00511_;
  wire [1:0] _00512_;
  wire [1:0] _00513_;
  wire [1:0] _00514_;
  wire [1:0] _00515_;
  wire [1:0] _00516_;
  wire [1:0] _00517_;
  wire [1:0] _00518_;
  wire [1:0] _00519_;
  wire [2:0] _00520_;
  wire [1:0] _00521_;
  wire [2:0] _00522_;
  wire [1:0] _00523_;
  wire [2:0] _00524_;
  wire [1:0] _00525_;
  wire [2:0] _00526_;
  wire [1:0] _00527_;
  wire [2:0] _00528_;
  wire [1:0] _00529_;
  wire [2:0] _00530_;
  wire [1:0] _00531_;
  wire [2:0] _00532_;
  wire [1:0] _00533_;
  wire [2:0] _00534_;
  wire [1:0] _00535_;
  wire [2:0] _00536_;
  wire [1:0] _00537_;
  wire [2:0] _00538_;
  wire [1:0] _00539_;
  wire [2:0] _00540_;
  wire [1:0] _00541_;
  wire [2:0] _00542_;
  wire [1:0] _00543_;
  wire [2:0] _00544_;
  wire [1:0] _00545_;
  wire [2:0] _00546_;
  wire [1:0] _00547_;
  wire [2:0] _00548_;
  wire [1:0] _00549_;
  wire [2:0] _00550_;
  wire [1:0] _00551_;
  wire [2:0] _00552_;
  wire [1:0] _00553_;
  wire [2:0] _00554_;
  wire [1:0] _00555_;
  wire [2:0] _00556_;
  wire [1:0] _00557_;
  wire [2:0] _00558_;
  wire [1:0] _00559_;
  wire [2:0] _00560_;
  wire [1:0] _00561_;
  wire [2:0] _00562_;
  wire [1:0] _00563_;
  wire [2:0] _00564_;
  wire [1:0] _00565_;
  wire [2:0] _00566_;
  wire [1:0] _00567_;
  wire [2:0] _00568_;
  wire [1:0] _00569_;
  wire [2:0] _00570_;
  wire [1:0] _00571_;
  wire [2:0] _00572_;
  wire [1:0] _00573_;
  wire [2:0] _00574_;
  wire [1:0] _00575_;
  wire [2:0] _00576_;
  wire [1:0] _00577_;
  wire [2:0] _00578_;
  wire [1:0] _00579_;
  wire [2:0] _00580_;
  wire [1:0] _00581_;
  wire [2:0] _00582_;
  wire [1:0] _00583_;
  wire [1:0] _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire [2:0] _00618_;
  wire _00619_;
  wire [2:0] _00620_;
  wire _00621_;
  wire [2:0] _00622_;
  wire _00623_;
  wire [1:0] _00624_;
  wire [1:0] _00625_;
  wire [1:0] _00626_;
  wire [1:0] _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire [1:0] _00726_;
  wire _00727_;
  wire [1:0] _00728_;
  wire _00729_;
  wire [1:0] _00730_;
  wire _00731_;
  wire [1:0] _00732_;
  wire _00733_;
  wire [1:0] _00734_;
  wire _00735_;
  wire [1:0] _00736_;
  wire _00737_;
  wire [1:0] _00738_;
  wire _00739_;
  wire [1:0] _00740_;
  wire _00741_;
  wire [1:0] _00742_;
  wire _00743_;
  wire [1:0] _00744_;
  wire _00745_;
  wire [1:0] _00746_;
  wire _00747_;
  wire [1:0] _00748_;
  wire _00749_;
  wire [1:0] _00750_;
  wire _00751_;
  wire [1:0] _00752_;
  wire _00753_;
  wire [1:0] _00754_;
  wire _00755_;
  wire [1:0] _00756_;
  wire _00757_;
  wire [1:0] _00758_;
  wire _00759_;
  wire [1:0] _00760_;
  wire _00761_;
  wire [1:0] _00762_;
  wire _00763_;
  wire [1:0] _00764_;
  wire _00765_;
  wire [1:0] _00766_;
  wire _00767_;
  wire [1:0] _00768_;
  wire _00769_;
  wire [1:0] _00770_;
  wire _00771_;
  wire [1:0] _00772_;
  wire _00773_;
  wire [1:0] _00774_;
  wire _00775_;
  wire [1:0] _00776_;
  wire _00777_;
  wire [1:0] _00778_;
  wire _00779_;
  wire [1:0] _00780_;
  wire _00781_;
  wire [1:0] _00782_;
  wire _00783_;
  wire [1:0] _00784_;
  wire _00785_;
  wire [1:0] _00786_;
  wire _00787_;
  wire [1:0] _00788_;
  wire _00789_;
  wire [1:0] _00790_;
  wire _00791_;
  wire [1:0] _00792_;
  wire [1:0] _00793_;
  wire [1:0] _00794_;
  wire [2:0] _00795_;
  wire [1:0] _00796_;
  wire [2:0] _00797_;
  wire [1:0] _00798_;
  wire [2:0] _00799_;
  wire [1:0] _00800_;
  wire [2:0] _00801_;
  wire [1:0] _00802_;
  wire [2:0] _00803_;
  wire [1:0] _00804_;
  wire [2:0] _00805_;
  wire [1:0] _00806_;
  wire [1:0] _00807_;
  wire [1:0] _00808_;
  wire _00809_;
  wire _00810_;
  wire [1:0] _00811_;
  wire [1:0] _00812_;
  wire [1:0] _00813_;
  wire [1:0] _00814_;
  wire [1:0] _00815_;
  wire [1:0] _00816_;
  wire [1:0] _00817_;
  wire [1:0] _00818_;
  wire [1:0] _00819_;
  wire [1:0] _00820_;
  wire [1:0] _00821_;
  wire [1:0] _00822_;
  wire [1:0] _00823_;
  wire [1:0] _00824_;
  wire [1:0] _00825_;
  wire [1:0] _00826_;
  wire [1:0] _00827_;
  wire [1:0] _00828_;
  wire [1:0] _00829_;
  wire [1:0] _00830_;
  wire [1:0] _00831_;
  wire [1:0] _00832_;
  wire [1:0] _00833_;
  wire [1:0] _00834_;
  wire [1:0] _00835_;
  wire [1:0] _00836_;
  wire [1:0] _00837_;
  wire [1:0] _00838_;
  wire [1:0] _00839_;
  wire [1:0] _00840_;
  wire [1:0] _00841_;
  wire [1:0] _00842_;
  wire [1:0] _00843_;
  wire [2:0] _00844_;
  wire [1:0] _00845_;
  wire [2:0] _00846_;
  wire [1:0] _00847_;
  wire [2:0] _00848_;
  wire [1:0] _00849_;
  wire [2:0] _00850_;
  wire [1:0] _00851_;
  wire [2:0] _00852_;
  wire [1:0] _00853_;
  wire [2:0] _00854_;
  wire [1:0] _00855_;
  wire [2:0] _00856_;
  wire [1:0] _00857_;
  wire [2:0] _00858_;
  wire [1:0] _00859_;
  wire [2:0] _00860_;
  wire [1:0] _00861_;
  wire [2:0] _00862_;
  wire [1:0] _00863_;
  wire [2:0] _00864_;
  wire [1:0] _00865_;
  wire [2:0] _00866_;
  wire [1:0] _00867_;
  wire [2:0] _00868_;
  wire [1:0] _00869_;
  wire [2:0] _00870_;
  wire [1:0] _00871_;
  wire [2:0] _00872_;
  wire [1:0] _00873_;
  wire [2:0] _00874_;
  wire [1:0] _00875_;
  wire [2:0] _00876_;
  wire [1:0] _00877_;
  wire [2:0] _00878_;
  wire [1:0] _00879_;
  wire [2:0] _00880_;
  wire [1:0] _00881_;
  wire [2:0] _00882_;
  wire [1:0] _00883_;
  wire [2:0] _00884_;
  wire [1:0] _00885_;
  wire [2:0] _00886_;
  wire [1:0] _00887_;
  wire [2:0] _00888_;
  wire [1:0] _00889_;
  wire [2:0] _00890_;
  wire [1:0] _00891_;
  wire [2:0] _00892_;
  wire [1:0] _00893_;
  wire [2:0] _00894_;
  wire [1:0] _00895_;
  wire [2:0] _00896_;
  wire [1:0] _00897_;
  wire [2:0] _00898_;
  wire [1:0] _00899_;
  wire [2:0] _00900_;
  wire [1:0] _00901_;
  wire [2:0] _00902_;
  wire [1:0] _00903_;
  wire [2:0] _00904_;
  wire [1:0] _00905_;
  wire [2:0] _00906_;
  wire [1:0] _00907_;
  wire [1:0] _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire [2:0] _00942_;
  wire _00943_;
  wire [2:0] _00944_;
  wire _00945_;
  wire [2:0] _00946_;
  wire _00947_;
  wire [1:0] _00948_;
  wire [1:0] _00949_;
  wire [1:0] _00950_;
  wire [1:0] _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire [1:0] _01050_;
  wire _01051_;
  wire [1:0] _01052_;
  wire _01053_;
  wire [1:0] _01054_;
  wire _01055_;
  wire [1:0] _01056_;
  wire _01057_;
  wire [1:0] _01058_;
  wire _01059_;
  wire [1:0] _01060_;
  wire _01061_;
  wire [1:0] _01062_;
  wire _01063_;
  wire [1:0] _01064_;
  wire _01065_;
  wire [1:0] _01066_;
  wire _01067_;
  wire [1:0] _01068_;
  wire _01069_;
  wire [1:0] _01070_;
  wire _01071_;
  wire [1:0] _01072_;
  wire _01073_;
  wire [1:0] _01074_;
  wire _01075_;
  wire [1:0] _01076_;
  wire _01077_;
  wire [1:0] _01078_;
  wire _01079_;
  wire [1:0] _01080_;
  wire _01081_;
  wire [1:0] _01082_;
  wire _01083_;
  wire [1:0] _01084_;
  wire _01085_;
  wire [1:0] _01086_;
  wire _01087_;
  wire [1:0] _01088_;
  wire _01089_;
  wire [1:0] _01090_;
  wire _01091_;
  wire [1:0] _01092_;
  wire _01093_;
  wire [1:0] _01094_;
  wire _01095_;
  wire [1:0] _01096_;
  wire _01097_;
  wire [1:0] _01098_;
  wire _01099_;
  wire [1:0] _01100_;
  wire _01101_;
  wire [1:0] _01102_;
  wire _01103_;
  wire [1:0] _01104_;
  wire _01105_;
  wire [1:0] _01106_;
  wire _01107_;
  wire [1:0] _01108_;
  wire _01109_;
  wire [1:0] _01110_;
  wire _01111_;
  wire [1:0] _01112_;
  wire _01113_;
  wire [1:0] _01114_;
  wire _01115_;
  wire [1:0] _01116_;
  wire [1:0] _01117_;
  wire [1:0] _01118_;
  wire [2:0] _01119_;
  wire [1:0] _01120_;
  wire [2:0] _01121_;
  wire [1:0] _01122_;
  wire [2:0] _01123_;
  wire [1:0] _01124_;
  wire [2:0] _01125_;
  wire [1:0] _01126_;
  wire [2:0] _01127_;
  wire [1:0] _01128_;
  wire [2:0] _01129_;
  wire [1:0] _01130_;
  wire [1:0] _01131_;
  wire [1:0] _01132_;
  wire _01133_;
  wire _01134_;
  wire [1:0] _01135_;
  wire [1:0] _01136_;
  wire [1:0] _01137_;
  wire [1:0] _01138_;
  wire [1:0] _01139_;
  wire [1:0] _01140_;
  wire [1:0] _01141_;
  wire [1:0] _01142_;
  wire [1:0] _01143_;
  wire [1:0] _01144_;
  wire [1:0] _01145_;
  wire [1:0] _01146_;
  wire [1:0] _01147_;
  wire [1:0] _01148_;
  wire [1:0] _01149_;
  wire [1:0] _01150_;
  wire [1:0] _01151_;
  wire [1:0] _01152_;
  wire [1:0] _01153_;
  wire [1:0] _01154_;
  wire [1:0] _01155_;
  wire [1:0] _01156_;
  wire [1:0] _01157_;
  wire [1:0] _01158_;
  wire [1:0] _01159_;
  wire [1:0] _01160_;
  wire [1:0] _01161_;
  wire [1:0] _01162_;
  wire [1:0] _01163_;
  wire [1:0] _01164_;
  wire [1:0] _01165_;
  wire [1:0] _01166_;
  wire [1:0] _01167_;
  wire [2:0] _01168_;
  wire [1:0] _01169_;
  wire [2:0] _01170_;
  wire [1:0] _01171_;
  wire [2:0] _01172_;
  wire [1:0] _01173_;
  wire [2:0] _01174_;
  wire [1:0] _01175_;
  wire [2:0] _01176_;
  wire [1:0] _01177_;
  wire [2:0] _01178_;
  wire [1:0] _01179_;
  wire [2:0] _01180_;
  wire [1:0] _01181_;
  wire [2:0] _01182_;
  wire [1:0] _01183_;
  wire [2:0] _01184_;
  wire [1:0] _01185_;
  wire [2:0] _01186_;
  wire [1:0] _01187_;
  wire [2:0] _01188_;
  wire [1:0] _01189_;
  wire [2:0] _01190_;
  wire [1:0] _01191_;
  wire [2:0] _01192_;
  wire [1:0] _01193_;
  wire [2:0] _01194_;
  wire [1:0] _01195_;
  wire [2:0] _01196_;
  wire [1:0] _01197_;
  wire [2:0] _01198_;
  wire [1:0] _01199_;
  wire [2:0] _01200_;
  wire [1:0] _01201_;
  wire [2:0] _01202_;
  wire [1:0] _01203_;
  wire [2:0] _01204_;
  wire [1:0] _01205_;
  wire [2:0] _01206_;
  wire [1:0] _01207_;
  wire [2:0] _01208_;
  wire [1:0] _01209_;
  wire [2:0] _01210_;
  wire [1:0] _01211_;
  wire [2:0] _01212_;
  wire [1:0] _01213_;
  wire [2:0] _01214_;
  wire [1:0] _01215_;
  wire [2:0] _01216_;
  wire [1:0] _01217_;
  wire [2:0] _01218_;
  wire [1:0] _01219_;
  wire [2:0] _01220_;
  wire [1:0] _01221_;
  wire [2:0] _01222_;
  wire [1:0] _01223_;
  wire [2:0] _01224_;
  wire [1:0] _01225_;
  wire [2:0] _01226_;
  wire [1:0] _01227_;
  wire [2:0] _01228_;
  wire [1:0] _01229_;
  wire [2:0] _01230_;
  wire [1:0] _01231_;
  wire [1:0] _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire [2:0] _01266_;
  wire _01267_;
  wire [2:0] _01268_;
  wire _01269_;
  wire [2:0] _01270_;
  wire _01271_;
  wire [1:0] _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire [1:0] _01276_;
  wire [1:0] _01277_;
  wire _01278_;
  wire [1:0] _01279_;
  wire [1:0] _01280_;
  wire [1:0] _01281_;
  wire _01282_;
  wire [1:0] _01283_;
  wire _01284_;
  wire [1:0] _01285_;
  wire _01286_;
  wire [2:0] _01287_;
  wire [1:0] _01288_;
  wire [1:0] _01289_;
  wire [2:0] _01290_;
  wire [1:0] _01291_;
  wire [1:0] _01292_;
  wire [2:0] _01293_;
  wire [1:0] _01294_;
  wire [1:0] _01295_;
  wire [2:0] _01296_;
  wire [1:0] _01297_;
  wire [1:0] _01298_;
  wire [2:0] _01299_;
  wire [1:0] _01300_;
  wire [1:0] _01301_;
  wire [2:0] _01302_;
  wire [1:0] _01303_;
  wire [1:0] _01304_;
  wire [2:0] _01305_;
  wire [1:0] _01306_;
  wire [1:0] _01307_;
  wire [2:0] _01308_;
  wire [1:0] _01309_;
  wire [1:0] _01310_;
  wire [2:0] _01311_;
  wire [1:0] _01312_;
  wire [1:0] _01313_;
  wire [2:0] _01314_;
  wire [1:0] _01315_;
  wire [1:0] _01316_;
  wire [2:0] _01317_;
  wire [1:0] _01318_;
  wire [1:0] _01319_;
  wire [2:0] _01320_;
  wire [1:0] _01321_;
  wire [1:0] _01322_;
  wire [2:0] _01323_;
  wire [1:0] _01324_;
  wire [1:0] _01325_;
  wire [2:0] _01326_;
  wire [1:0] _01327_;
  wire [1:0] _01328_;
  wire [2:0] _01329_;
  wire [1:0] _01330_;
  wire [1:0] _01331_;
  wire [2:0] _01332_;
  wire [1:0] _01333_;
  wire [2:0] _01334_;
  wire _01335_;
  wire [1:0] _01336_;
  wire _01337_;
  wire [1:0] _01338_;
  wire [1:0] _01339_;
  wire _01340_;
  wire [1:0] _01341_;
  wire _01342_;
  wire [1:0] _01343_;
  wire [1:0] _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire [1:0] _01348_;
  wire [1:0] _01349_;
  wire _01350_;
  wire [1:0] _01351_;
  wire [1:0] _01352_;
  wire [1:0] _01353_;
  wire _01354_;
  wire [1:0] _01355_;
  wire _01356_;
  wire [1:0] _01357_;
  wire _01358_;
  wire [2:0] _01359_;
  wire [1:0] _01360_;
  wire [1:0] _01361_;
  wire [2:0] _01362_;
  wire [1:0] _01363_;
  wire [1:0] _01364_;
  wire [2:0] _01365_;
  wire [1:0] _01366_;
  wire [1:0] _01367_;
  wire [2:0] _01368_;
  wire [1:0] _01369_;
  wire [1:0] _01370_;
  wire [2:0] _01371_;
  wire [1:0] _01372_;
  wire [1:0] _01373_;
  wire [2:0] _01374_;
  wire [1:0] _01375_;
  wire [1:0] _01376_;
  wire [2:0] _01377_;
  wire [1:0] _01378_;
  wire [1:0] _01379_;
  wire [2:0] _01380_;
  wire [1:0] _01381_;
  wire [1:0] _01382_;
  wire [2:0] _01383_;
  wire [1:0] _01384_;
  wire [1:0] _01385_;
  wire [2:0] _01386_;
  wire [1:0] _01387_;
  wire [1:0] _01388_;
  wire [2:0] _01389_;
  wire [1:0] _01390_;
  wire [1:0] _01391_;
  wire [2:0] _01392_;
  wire [1:0] _01393_;
  wire [1:0] _01394_;
  wire [2:0] _01395_;
  wire [1:0] _01396_;
  wire [1:0] _01397_;
  wire [2:0] _01398_;
  wire [1:0] _01399_;
  wire [1:0] _01400_;
  wire [2:0] _01401_;
  wire [1:0] _01402_;
  wire [1:0] _01403_;
  wire [2:0] _01404_;
  wire [1:0] _01405_;
  wire [2:0] _01406_;
  wire _01407_;
  wire [1:0] _01408_;
  wire _01409_;
  wire [1:0] _01410_;
  wire [1:0] _01411_;
  wire _01412_;
  wire [1:0] _01413_;
  wire _01414_;
  wire [1:0] _01415_;
  wire [1:0] _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire [1:0] _01420_;
  wire [1:0] _01421_;
  wire _01422_;
  wire [1:0] _01423_;
  wire [1:0] _01424_;
  wire [1:0] _01425_;
  wire _01426_;
  wire [1:0] _01427_;
  wire _01428_;
  wire [1:0] _01429_;
  wire _01430_;
  wire [2:0] _01431_;
  wire [1:0] _01432_;
  wire [1:0] _01433_;
  wire [2:0] _01434_;
  wire [1:0] _01435_;
  wire [1:0] _01436_;
  wire [2:0] _01437_;
  wire [1:0] _01438_;
  wire [1:0] _01439_;
  wire [2:0] _01440_;
  wire [1:0] _01441_;
  wire [1:0] _01442_;
  wire [2:0] _01443_;
  wire [1:0] _01444_;
  wire [1:0] _01445_;
  wire [2:0] _01446_;
  wire [1:0] _01447_;
  wire [1:0] _01448_;
  wire [2:0] _01449_;
  wire [1:0] _01450_;
  wire [1:0] _01451_;
  wire [2:0] _01452_;
  wire [1:0] _01453_;
  wire [1:0] _01454_;
  wire [2:0] _01455_;
  wire [1:0] _01456_;
  wire [1:0] _01457_;
  wire [2:0] _01458_;
  wire [1:0] _01459_;
  wire [1:0] _01460_;
  wire [2:0] _01461_;
  wire [1:0] _01462_;
  wire [1:0] _01463_;
  wire [2:0] _01464_;
  wire [1:0] _01465_;
  wire [1:0] _01466_;
  wire [2:0] _01467_;
  wire [1:0] _01468_;
  wire [1:0] _01469_;
  wire [2:0] _01470_;
  wire [1:0] _01471_;
  wire [1:0] _01472_;
  wire [2:0] _01473_;
  wire [1:0] _01474_;
  wire [1:0] _01475_;
  wire [2:0] _01476_;
  wire [1:0] _01477_;
  wire [2:0] _01478_;
  wire _01479_;
  wire [1:0] _01480_;
  wire _01481_;
  wire [1:0] _01482_;
  wire [1:0] _01483_;
  wire _01484_;
  wire [1:0] _01485_;
  wire _01486_;
  wire [1:0] _01487_;
  wire _01488_;
  wire [1:0] _01489_;
  wire _01490_;
  wire [1:0] _01491_;
  wire [1:0] _01492_;
  wire [1:0] _01493_;
  wire _01494_;
  wire [2:0] _01495_;
  wire [1:0] _01496_;
  wire _01497_;
  wire [1:0] _01498_;
  wire _01499_;
  wire [1:0] _01500_;
  wire [1:0] _01501_;
  wire [1:0] _01502_;
  wire _01503_;
  wire [2:0] _01504_;
  wire [1:0] _01505_;
  wire [8:0] _01506_;
  wire [3:0] _01507_;
  wire [1:0] _01508_;
  wire _01509_;
  wire [7:0] _01510_;
  wire [3:0] _01511_;
  wire _01512_;
  wire [1:0] _01513_;
  wire _01514_;
  wire [1:0] _01515_;
  wire _01516_;
  wire [3:0] _01517_;
  wire [1:0] _01518_;
  wire _01519_;
  wire [7:0] _01520_;
  wire [3:0] _01521_;
  wire [1:0] _01522_;
  wire [1:0] _01523_;
  wire _01524_;
  wire [6:0] _01525_;
  wire [3:0] _01526_;
  wire [1:0] _01527_;
  wire [1:0] _01528_;
  wire [1:0] _01529_;
  wire [7:0] _01530_;
  wire [3:0] _01531_;
  wire [1:0] _01532_;
  wire _01533_;
  wire _01534_;
  wire [2:0] _01535_;
  wire [1:0] _01536_;
  wire [6:0] _01537_;
  wire [3:0] _01538_;
  wire [1:0] _01539_;
  wire [7:0] _01540_;
  wire [3:0] _01541_;
  wire [1:0] _01542_;
  wire _01543_;
  wire [3:0] _01544_;
  wire [1:0] _01545_;
  wire _01546_;
  wire [8:0] _01547_;
  wire [3:0] _01548_;
  wire [1:0] _01549_;
  wire _01550_;
  wire [7:0] _01551_;
  wire [3:0] _01552_;
  wire [1:0] _01553_;
  wire _01554_;
  wire [7:0] _01555_;
  wire [3:0] _01556_;
  wire [1:0] _01557_;
  wire _01558_;
  wire [6:0] _01559_;
  wire [3:0] _01560_;
  wire [1:0] _01561_;
  wire [7:0] _01562_;
  wire [3:0] _01563_;
  wire [1:0] _01564_;
  wire _01565_;
  wire [6:0] _01566_;
  wire [3:0] _01567_;
  wire [1:0] _01568_;
  wire [7:0] _01569_;
  wire [3:0] _01570_;
  wire [1:0] _01571_;
  wire _01572_;
  wire _01573_;
  wire [15:0] _01574_;
  wire [7:0] _01575_;
  wire [3:0] _01576_;
  wire [1:0] _01577_;
  wire [15:0] _01578_;
  wire [7:0] _01579_;
  wire [3:0] _01580_;
  wire [1:0] _01581_;
  wire [8:0] _01582_;
  wire [3:0] _01583_;
  wire [1:0] _01584_;
  wire _01585_;
  wire [3:0] _01586_;
  wire [1:0] _01587_;
  wire [3:0] _01588_;
  wire [1:0] _01589_;
  wire [3:0] _01590_;
  wire [1:0] _01591_;
  wire [3:0] _01592_;
  wire [1:0] _01593_;
  wire [3:0] _01594_;
  wire [1:0] _01595_;
  wire [1:0] _01596_;
  wire [3:0] _01597_;
  wire [1:0] _01598_;
  wire [3:0] _01599_;
  wire [1:0] _01600_;
  wire [1:0] _01601_;
  wire [3:0] _01602_;
  wire [1:0] _01603_;
  wire [1:0] _01604_;
  wire [1:0] _01605_;
  wire [1:0] _01606_;
  wire [1:0] _01607_;
  wire _01608_;
  wire [7:0] _01609_;
  wire [3:0] _01610_;
  wire [1:0] _01611_;
  wire [11:0] _01612_;
  wire [5:0] _01613_;
  wire [2:0] _01614_;
  wire _01615_;
  wire [7:0] _01616_;
  wire [3:0] _01617_;
  wire [1:0] _01618_;
  wire _01619_;
  wire [8:0] _01620_;
  wire [3:0] _01621_;
  wire [1:0] _01622_;
  wire _01623_;
  wire [7:0] _01624_;
  wire [3:0] _01625_;
  wire [1:0] _01626_;
  wire _01627_;
  wire _01628_;
  wire [15:0] _01629_;
  wire [7:0] _01630_;
  wire [3:0] _01631_;
  wire [1:0] _01632_;
  wire [15:0] _01633_;
  wire [7:0] _01634_;
  wire [3:0] _01635_;
  wire [1:0] _01636_;
  wire [8:0] _01637_;
  wire [3:0] _01638_;
  wire [1:0] _01639_;
  wire _01640_;
  wire [3:0] _01641_;
  wire [1:0] _01642_;
  wire [3:0] _01643_;
  wire [1:0] _01644_;
  wire [3:0] _01645_;
  wire [1:0] _01646_;
  wire [3:0] _01647_;
  wire [1:0] _01648_;
  wire [3:0] _01649_;
  wire [1:0] _01650_;
  wire [1:0] _01651_;
  wire [3:0] _01652_;
  wire [1:0] _01653_;
  wire [3:0] _01654_;
  wire [1:0] _01655_;
  wire [1:0] _01656_;
  wire [3:0] _01657_;
  wire [1:0] _01658_;
  wire [1:0] _01659_;
  wire [1:0] _01660_;
  wire [1:0] _01661_;
  wire [1:0] _01662_;
  wire _01663_;
  wire [7:0] _01664_;
  wire [3:0] _01665_;
  wire [1:0] _01666_;
  wire [11:0] _01667_;
  wire [5:0] _01668_;
  wire [2:0] _01669_;
  wire _01670_;
  wire _01671_;
  wire [15:0] _01672_;
  wire [7:0] _01673_;
  wire [3:0] _01674_;
  wire [1:0] _01675_;
  wire [15:0] _01676_;
  wire [7:0] _01677_;
  wire [3:0] _01678_;
  wire [1:0] _01679_;
  wire [6:0] _01680_;
  wire [3:0] _01681_;
  wire [1:0] _01682_;
  wire [7:0] _01683_;
  wire [3:0] _01684_;
  wire [1:0] _01685_;
  wire _01686_;
  wire [8:0] _01687_;
  wire [3:0] _01688_;
  wire [1:0] _01689_;
  wire _01690_;
  wire [3:0] _01691_;
  wire [1:0] _01692_;
  wire [3:0] _01693_;
  wire [1:0] _01694_;
  wire [3:0] _01695_;
  wire [1:0] _01696_;
  wire [3:0] _01697_;
  wire [1:0] _01698_;
  wire [3:0] _01699_;
  wire [1:0] _01700_;
  wire [1:0] _01701_;
  wire [3:0] _01702_;
  wire [1:0] _01703_;
  wire [3:0] _01704_;
  wire [1:0] _01705_;
  wire [1:0] _01706_;
  wire [3:0] _01707_;
  wire [1:0] _01708_;
  wire [1:0] _01709_;
  wire [1:0] _01710_;
  wire [1:0] _01711_;
  wire [1:0] _01712_;
  wire _01713_;
  wire [7:0] _01714_;
  wire [3:0] _01715_;
  wire [1:0] _01716_;
  wire [3:0] _01717_;
  wire [1:0] _01718_;
  wire _01719_;
  wire [11:0] _01720_;
  wire [5:0] _01721_;
  wire [2:0] _01722_;
  wire _01723_;
  wire [6:0] _01724_;
  wire [3:0] _01725_;
  wire [1:0] _01726_;
  wire [7:0] _01727_;
  wire [3:0] _01728_;
  wire [1:0] _01729_;
  wire _01730_;
  wire [1:0] _01731_;
  wire [1:0] _01732_;
  wire [1:0] _01733_;
  wire [1:0] _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire [1:0] _01744_;
  wire _01745_;
  wire [1:0] _01746_;
  wire _01747_;
  wire [1:0] _01748_;
  wire _01749_;
  wire [15:0] _01750_;
  wire [7:0] _01751_;
  wire [3:0] _01752_;
  wire [1:0] _01753_;
  wire _01754_;
  wire [15:0] _01755_;
  wire [7:0] _01756_;
  wire [3:0] _01757_;
  wire [1:0] _01758_;
  wire _01759_;
  wire [15:0] _01760_;
  wire [7:0] _01761_;
  wire [3:0] _01762_;
  wire [1:0] _01763_;
  wire _01764_;
  wire [4:0] _01765_;
  wire [2:0] _01766_;
  wire [4:0] _01767_;
  wire [2:0] _01768_;
  wire [4:0] _01769_;
  wire [2:0] _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire [15:0] _01835_;
  wire [3:0] _01836_;
  wire [15:0] _01837_;
  wire [3:0] _01838_;
  wire [15:0] _01839_;
  wire [3:0] _01840_;
  wire [15:0] _01841_;
  wire [7:0] _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire [7:0] _01846_;
  wire [15:0] _01847_;
  wire [15:0] _01848_;
  wire [15:0] _01849_;
  wire [15:0] _01850_;
  wire [7:0] _01851_;
  wire [7:0] _01852_;
  wire [3:0] _01853_;
  wire [3:0] _01854_;
  wire [3:0] _01855_;
  wire _01856_;
  wire [3:0] _01857_;
  wire [3:0] _01858_;
  wire [3:0] _01859_;
  wire _01860_;
  wire [3:0] _01861_;
  wire [3:0] _01862_;
  wire [3:0] _01863_;
  wire _01864_;
  wire [2:0] _01865_;
  wire [2:0] _01866_;
  wire _01867_;
  wire [2:0] _01868_;
  wire [2:0] _01869_;
  wire [2:0] _01870_;
  wire _01871_;
  wire [1:0] _01872_;
  wire [1:0] _01873_;
  wire [1:0] _01874_;
  wire _01875_;
  wire [31:0] _01876_;
  wire [2:0] _01877_;
  wire [511:0] _01878_;
  wire [32:0] _01879_;
  wire [255:0] _01880_;
  wire [29:0] _01881_;
  wire [11:0] _01882_;
  wire [7:0] _01883_;
  wire [6:0] _01884_;
  wire [7:0] _01885_;
  wire [6:0] _01886_;
  wire [7:0] _01887_;
  wire [6:0] _01888_;
  wire [7:0] _01889_;
  wire [6:0] _01890_;
  wire [7:0] _01891_;
  wire [511:0] _01892_;
  wire [511:0] _01893_;
  wire [63:0] _01894_;
  wire [3:0] _01895_;
  wire [1023:0] _01896_;
  wire [32:0] _01897_;
  wire [127:0] _01898_;
  wire [7:0] _01899_;
  wire [127:0] _01900_;
  wire [7:0] _01901_;
  wire [127:0] _01902_;
  wire [7:0] _01903_;
  wire [127:0] _01904_;
  wire [7:0] _01905_;
  wire [127:0] _01906_;
  wire [7:0] _01907_;
  wire [127:0] _01908_;
  wire [7:0] _01909_;
  wire [127:0] _01910_;
  wire [7:0] _01911_;
  wire [127:0] _01912_;
  wire [7:0] _01913_;
  wire [127:0] _01914_;
  wire [7:0] _01915_;
  wire [127:0] _01916_;
  wire [7:0] _01917_;
  wire [127:0] _01918_;
  wire [7:0] _01919_;
  wire [127:0] _01920_;
  wire [7:0] _01921_;
  wire [127:0] _01922_;
  wire [7:0] _01923_;
  wire [127:0] _01924_;
  wire [7:0] _01925_;
  wire [127:0] _01926_;
  wire [7:0] _01927_;
  wire [127:0] _01928_;
  wire [7:0] _01929_;
  wire [127:0] _01930_;
  wire [4:0] _01931_;
  wire [127:0] _01932_;
  wire [4:0] _01933_;
  wire [511:0] _01934_;
  wire [511:0] _01935_;
  wire [255:0] _01936_;
  wire [255:0] _01937_;
  wire [1023:0] _01938_;
  wire [2:0] _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire [2:0] _01944_;
  wire [2:0] _01945_;
  wire [2:0] _01946_;
  wire [7:0] _01947_;
  wire [7:0] _01948_;
  wire [7:0] _01949_;
  wire [7:0] _01950_;
  wire [7:0] _01951_;
  wire [7:0] _01952_;
  wire [7:0] _01953_;
  wire [7:0] _01954_;
  wire [7:0] _01955_;
  wire [7:0] _01956_;
  wire [7:0] _01957_;
  wire [7:0] _01958_;
  wire [7:0] _01959_;
  wire [7:0] _01960_;
  wire [7:0] _01961_;
  wire [7:0] _01962_;
  wire [7:0] _01963_;
  wire [7:0] _01964_;
  wire [7:0] _01965_;
  wire [7:0] _01966_;
  wire [7:0] _01967_;
  wire [7:0] _01968_;
  wire [7:0] _01969_;
  wire [7:0] _01970_;
  wire [7:0] _01971_;
  wire [7:0] _01972_;
  wire [7:0] _01973_;
  wire [7:0] _01974_;
  wire [7:0] _01975_;
  wire [7:0] _01976_;
  wire [7:0] _01977_;
  wire [7:0] _01978_;
  wire _01979_;
  wire [7:0] _01980_;
  wire [7:0] _01981_;
  wire [7:0] _01982_;
  wire [7:0] _01983_;
  wire [7:0] _01984_;
  wire [7:0] _01985_;
  wire [7:0] _01986_;
  wire [7:0] _01987_;
  wire [7:0] _01988_;
  wire [7:0] _01989_;
  wire [7:0] _01990_;
  wire [7:0] _01991_;
  wire [7:0] _01992_;
  wire [7:0] _01993_;
  wire [7:0] _01994_;
  wire [7:0] _01995_;
  wire [31:0] _01996_;
  wire _01997_;
  wire [31:0] _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire [31:0] _02009_;
  wire [31:0] _02010_;
  wire _02011_;
  wire _02012_;
  wire [14:0] _02013_;
  wire [15:0] _02014_;
  wire [31:0] _02015_;
  wire [31:0] _02016_;
  wire _02017_;
  wire _02018_;
  wire [31:0] _02019_;
  wire [4:0] _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire [31:0] _02026_;
  wire [3:0] _02027_;
  wire _02028_;
  wire [31:0] _02029_;
  wire [3:0] _02030_;
  wire [31:0] _02031_;
  wire _02032_;
  wire [31:0] _02033_;
  wire [3:0] _02034_;
  wire _02035_;
  wire _02036_;
  wire [31:0] _02037_;
  wire [4:0] _02038_;
  wire [2:0] _02039_;
  wire [2:0] _02040_;
  wire [2:0] _02041_;
  wire [2:0] _02042_;
  wire [2:0] _02043_;
  wire [31:0] _02044_;
  wire [4:0] _02045_;
  wire [31:0] _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire [3:0] _02065_;
  wire [4:0] _02066_;
  wire [7:0] _02067_;
  wire [7:0] _02068_;
  wire [7:0] _02069_;
  wire [7:0] _02070_;
  wire [7:0] _02071_;
  wire [7:0] _02072_;
  wire [7:0] _02073_;
  wire [7:0] _02074_;
  wire [7:0] _02075_;
  wire [7:0] _02076_;
  wire [7:0] _02077_;
  wire [7:0] _02078_;
  wire [7:0] _02079_;
  wire [7:0] _02080_;
  wire [7:0] _02081_;
  wire [7:0] _02082_;
  wire [2:0] _02083_;
  wire [223:0] _02084_;
  wire [223:0] _02085_;
  wire [6:0] _02086_;
  wire [31:0] _02087_;
  wire [34:0] _02088_;
  wire [34:0] _02089_;
  wire [6:0] _02090_;
  wire [4:0] _02091_;
  wire [95:0] _02092_;
  wire [95:0] _02093_;
  wire [2:0] _02094_;
  wire [31:0] _02095_;
  wire [159:0] _02096_;
  wire [159:0] _02097_;
  wire [4:0] _02098_;
  wire [31:0] _02099_;
  wire [95:0] _02100_;
  wire [95:0] _02101_;
  wire [2:0] _02102_;
  wire [31:0] _02103_;
  wire [127:0] _02104_;
  wire [127:0] _02105_;
  wire [31:0] _02106_;
  wire [44:0] _02107_;
  wire [44:0] _02108_;
  wire [2:0] _02109_;
  wire [14:0] _02110_;
  wire [47:0] _02111_;
  wire [47:0] _02112_;
  wire [15:0] _02113_;
  wire [95:0] _02114_;
  wire [95:0] _02115_;
  wire [2:0] _02116_;
  wire [31:0] _02117_;
  wire [7:0] _02118_;
  wire [7:0] _02119_;
  wire [1:0] _02120_;
  wire [3:0] _02121_;
  wire [3:0] _02122_;
  wire [15:0] _02123_;
  wire [3:0] _02124_;
  wire [3:0] _02125_;
  wire [3:0] _02126_;
  wire _02127_;
  wire [15:0] _02128_;
  wire [3:0] _02129_;
  wire [15:0] _02130_;
  wire [3:0] _02131_;
  wire [15:0] _02132_;
  wire [3:0] _02133_;
  wire [15:0] _02134_;
  wire [7:0] _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire [7:0] _02139_;
  wire [15:0] _02140_;
  wire [15:0] _02141_;
  wire [15:0] _02142_;
  wire [15:0] _02143_;
  wire [7:0] _02144_;
  wire [7:0] _02145_;
  wire [3:0] _02146_;
  wire [3:0] _02147_;
  wire [3:0] _02148_;
  wire _02149_;
  wire [3:0] _02150_;
  wire [3:0] _02151_;
  wire [3:0] _02152_;
  wire _02153_;
  wire [3:0] _02154_;
  wire [3:0] _02155_;
  wire [3:0] _02156_;
  wire _02157_;
  wire [2:0] _02158_;
  wire [2:0] _02159_;
  wire _02160_;
  wire [2:0] _02161_;
  wire [2:0] _02162_;
  wire [2:0] _02163_;
  wire _02164_;
  wire [1:0] _02165_;
  wire [1:0] _02166_;
  wire [1:0] _02167_;
  wire _02168_;
  wire [31:0] _02169_;
  wire [2:0] _02170_;
  wire [32:0] _02171_;
  wire [255:0] _02172_;
  wire [29:0] _02173_;
  wire [11:0] _02174_;
  wire [7:0] _02175_;
  wire [6:0] _02176_;
  wire [7:0] _02177_;
  wire [6:0] _02178_;
  wire [7:0] _02179_;
  wire [6:0] _02180_;
  wire [7:0] _02181_;
  wire [6:0] _02182_;
  wire [7:0] _02183_;
  wire [511:0] _02184_;
  wire [511:0] _02185_;
  wire [63:0] _02186_;
  wire [3:0] _02187_;
  wire [1023:0] _02188_;
  wire [32:0] _02189_;
  wire [127:0] _02190_;
  wire [7:0] _02191_;
  wire [127:0] _02192_;
  wire [7:0] _02193_;
  wire [127:0] _02194_;
  wire [7:0] _02195_;
  wire [127:0] _02196_;
  wire [7:0] _02197_;
  wire [127:0] _02198_;
  wire [7:0] _02199_;
  wire [127:0] _02200_;
  wire [7:0] _02201_;
  wire [127:0] _02202_;
  wire [7:0] _02203_;
  wire [127:0] _02204_;
  wire [7:0] _02205_;
  wire [127:0] _02206_;
  wire [7:0] _02207_;
  wire [127:0] _02208_;
  wire [7:0] _02209_;
  wire [127:0] _02210_;
  wire [7:0] _02211_;
  wire [127:0] _02212_;
  wire [7:0] _02213_;
  wire [127:0] _02214_;
  wire [7:0] _02215_;
  wire [127:0] _02216_;
  wire [7:0] _02217_;
  wire [127:0] _02218_;
  wire [7:0] _02219_;
  wire [127:0] _02220_;
  wire [7:0] _02221_;
  wire [127:0] _02222_;
  wire [4:0] _02223_;
  wire [127:0] _02224_;
  wire [4:0] _02225_;
  wire [511:0] _02226_;
  wire [511:0] _02227_;
  wire [255:0] _02228_;
  wire [255:0] _02229_;
  wire [1023:0] _02230_;
  wire [2:0] _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire [2:0] _02236_;
  wire [2:0] _02237_;
  wire [2:0] _02238_;
  wire [7:0] _02239_;
  wire [7:0] _02240_;
  wire [7:0] _02241_;
  wire [7:0] _02242_;
  wire [7:0] _02243_;
  wire [7:0] _02244_;
  wire [7:0] _02245_;
  wire [7:0] _02246_;
  wire [7:0] _02247_;
  wire [7:0] _02248_;
  wire [7:0] _02249_;
  wire [7:0] _02250_;
  wire [7:0] _02251_;
  wire [7:0] _02252_;
  wire [7:0] _02253_;
  wire [7:0] _02254_;
  wire [7:0] _02255_;
  wire [7:0] _02256_;
  wire [7:0] _02257_;
  wire [7:0] _02258_;
  wire [7:0] _02259_;
  wire [7:0] _02260_;
  wire [7:0] _02261_;
  wire [7:0] _02262_;
  wire [7:0] _02263_;
  wire [7:0] _02264_;
  wire [7:0] _02265_;
  wire [7:0] _02266_;
  wire [7:0] _02267_;
  wire [7:0] _02268_;
  wire [7:0] _02269_;
  wire [7:0] _02270_;
  wire _02271_;
  wire [7:0] _02272_;
  wire [7:0] _02273_;
  wire [7:0] _02274_;
  wire [7:0] _02275_;
  wire [7:0] _02276_;
  wire [7:0] _02277_;
  wire [7:0] _02278_;
  wire [7:0] _02279_;
  wire [7:0] _02280_;
  wire [7:0] _02281_;
  wire [7:0] _02282_;
  wire [7:0] _02283_;
  wire [7:0] _02284_;
  wire [7:0] _02285_;
  wire [7:0] _02286_;
  wire [7:0] _02287_;
  wire [31:0] _02288_;
  wire _02289_;
  wire [31:0] _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire [31:0] _02299_;
  wire [31:0] _02300_;
  wire _02301_;
  wire _02302_;
  wire [14:0] _02303_;
  wire [15:0] _02304_;
  wire [31:0] _02305_;
  wire [31:0] _02306_;
  wire _02307_;
  wire _02308_;
  wire [31:0] _02309_;
  wire [4:0] _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire [31:0] _02316_;
  wire [3:0] _02317_;
  wire _02318_;
  wire [31:0] _02319_;
  wire [3:0] _02320_;
  wire [31:0] _02321_;
  wire _02322_;
  wire [31:0] _02323_;
  wire [3:0] _02324_;
  wire _02325_;
  wire _02326_;
  wire [31:0] _02327_;
  wire [4:0] _02328_;
  wire [2:0] _02329_;
  wire [2:0] _02330_;
  wire [2:0] _02331_;
  wire [2:0] _02332_;
  wire [2:0] _02333_;
  wire [31:0] _02334_;
  wire [4:0] _02335_;
  wire [31:0] _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire [3:0] _02354_;
  wire [4:0] _02355_;
  wire [7:0] _02356_;
  wire [7:0] _02357_;
  wire [7:0] _02358_;
  wire [7:0] _02359_;
  wire [7:0] _02360_;
  wire [7:0] _02361_;
  wire [7:0] _02362_;
  wire [7:0] _02363_;
  wire [7:0] _02364_;
  wire [7:0] _02365_;
  wire [7:0] _02366_;
  wire [7:0] _02367_;
  wire [7:0] _02368_;
  wire [7:0] _02369_;
  wire [7:0] _02370_;
  wire [7:0] _02371_;
  wire [2:0] _02372_;
  wire [223:0] _02373_;
  wire [223:0] _02374_;
  wire [6:0] _02375_;
  wire [31:0] _02376_;
  wire [34:0] _02377_;
  wire [34:0] _02378_;
  wire [6:0] _02379_;
  wire [4:0] _02380_;
  wire [95:0] _02381_;
  wire [95:0] _02382_;
  wire [2:0] _02383_;
  wire [31:0] _02384_;
  wire [159:0] _02385_;
  wire [159:0] _02386_;
  wire [4:0] _02387_;
  wire [31:0] _02388_;
  wire [95:0] _02389_;
  wire [95:0] _02390_;
  wire [2:0] _02391_;
  wire [31:0] _02392_;
  wire [127:0] _02393_;
  wire [127:0] _02394_;
  wire [31:0] _02395_;
  wire [44:0] _02396_;
  wire [44:0] _02397_;
  wire [2:0] _02398_;
  wire [14:0] _02399_;
  wire [47:0] _02400_;
  wire [47:0] _02401_;
  wire [15:0] _02402_;
  wire [95:0] _02403_;
  wire [95:0] _02404_;
  wire [2:0] _02405_;
  wire [31:0] _02406_;
  wire [7:0] _02407_;
  wire [7:0] _02408_;
  wire [1:0] _02409_;
  wire [3:0] _02410_;
  wire [3:0] _02411_;
  wire [15:0] _02412_;
  wire [3:0] _02413_;
  wire [3:0] _02414_;
  wire [3:0] _02415_;
  wire _02416_;
  wire [15:0] _02417_;
  wire [3:0] _02418_;
  wire [15:0] _02419_;
  wire [3:0] _02420_;
  wire [15:0] _02421_;
  wire [3:0] _02422_;
  wire [15:0] _02423_;
  wire [7:0] _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire [7:0] _02428_;
  wire [15:0] _02429_;
  wire [15:0] _02430_;
  wire [15:0] _02431_;
  wire [15:0] _02432_;
  wire [7:0] _02433_;
  wire [7:0] _02434_;
  wire [3:0] _02435_;
  wire [3:0] _02436_;
  wire [3:0] _02437_;
  wire _02438_;
  wire [3:0] _02439_;
  wire [3:0] _02440_;
  wire [3:0] _02441_;
  wire _02442_;
  wire [3:0] _02443_;
  wire [3:0] _02444_;
  wire [3:0] _02445_;
  wire _02446_;
  wire [2:0] _02447_;
  wire [2:0] _02448_;
  wire _02449_;
  wire [2:0] _02450_;
  wire [2:0] _02451_;
  wire [2:0] _02452_;
  wire _02453_;
  wire [1:0] _02454_;
  wire [1:0] _02455_;
  wire [1:0] _02456_;
  wire _02457_;
  wire [31:0] _02458_;
  wire [2:0] _02459_;
  wire [32:0] _02460_;
  wire [255:0] _02461_;
  wire [29:0] _02462_;
  wire [11:0] _02463_;
  wire [7:0] _02464_;
  wire [6:0] _02465_;
  wire [7:0] _02466_;
  wire [6:0] _02467_;
  wire [7:0] _02468_;
  wire [6:0] _02469_;
  wire [7:0] _02470_;
  wire [6:0] _02471_;
  wire [7:0] _02472_;
  wire [511:0] _02473_;
  wire [511:0] _02474_;
  wire [63:0] _02475_;
  wire [3:0] _02476_;
  wire [1023:0] _02477_;
  wire [32:0] _02478_;
  wire [127:0] _02479_;
  wire [7:0] _02480_;
  wire [127:0] _02481_;
  wire [7:0] _02482_;
  wire [127:0] _02483_;
  wire [7:0] _02484_;
  wire [127:0] _02485_;
  wire [7:0] _02486_;
  wire [127:0] _02487_;
  wire [7:0] _02488_;
  wire [127:0] _02489_;
  wire [7:0] _02490_;
  wire [127:0] _02491_;
  wire [7:0] _02492_;
  wire [127:0] _02493_;
  wire [7:0] _02494_;
  wire [127:0] _02495_;
  wire [7:0] _02496_;
  wire [127:0] _02497_;
  wire [7:0] _02498_;
  wire [127:0] _02499_;
  wire [7:0] _02500_;
  wire [127:0] _02501_;
  wire [7:0] _02502_;
  wire [127:0] _02503_;
  wire [7:0] _02504_;
  wire [127:0] _02505_;
  wire [7:0] _02506_;
  wire [127:0] _02507_;
  wire [7:0] _02508_;
  wire [127:0] _02509_;
  wire [7:0] _02510_;
  wire [127:0] _02511_;
  wire [4:0] _02512_;
  wire [127:0] _02513_;
  wire [4:0] _02514_;
  wire [511:0] _02515_;
  wire [511:0] _02516_;
  wire [255:0] _02517_;
  wire [255:0] _02518_;
  wire [1023:0] _02519_;
  wire [2:0] _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire [2:0] _02525_;
  wire [2:0] _02526_;
  wire [2:0] _02527_;
  wire [7:0] _02528_;
  wire [7:0] _02529_;
  wire [7:0] _02530_;
  wire [7:0] _02531_;
  wire [7:0] _02532_;
  wire [7:0] _02533_;
  wire [7:0] _02534_;
  wire [7:0] _02535_;
  wire [7:0] _02536_;
  wire [7:0] _02537_;
  wire [7:0] _02538_;
  wire [7:0] _02539_;
  wire [7:0] _02540_;
  wire [7:0] _02541_;
  wire [7:0] _02542_;
  wire [7:0] _02543_;
  wire [7:0] _02544_;
  wire [7:0] _02545_;
  wire [7:0] _02546_;
  wire [7:0] _02547_;
  wire [7:0] _02548_;
  wire [7:0] _02549_;
  wire [7:0] _02550_;
  wire [7:0] _02551_;
  wire [7:0] _02552_;
  wire [7:0] _02553_;
  wire [7:0] _02554_;
  wire [7:0] _02555_;
  wire [7:0] _02556_;
  wire [7:0] _02557_;
  wire [7:0] _02558_;
  wire [7:0] _02559_;
  wire _02560_;
  wire [7:0] _02561_;
  wire [7:0] _02562_;
  wire [7:0] _02563_;
  wire [7:0] _02564_;
  wire [7:0] _02565_;
  wire [7:0] _02566_;
  wire [7:0] _02567_;
  wire [7:0] _02568_;
  wire [7:0] _02569_;
  wire [7:0] _02570_;
  wire [7:0] _02571_;
  wire [7:0] _02572_;
  wire [7:0] _02573_;
  wire [7:0] _02574_;
  wire [7:0] _02575_;
  wire [7:0] _02576_;
  wire [31:0] _02577_;
  wire _02578_;
  wire [31:0] _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire [31:0] _02588_;
  wire [31:0] _02589_;
  wire _02590_;
  wire _02591_;
  wire [14:0] _02592_;
  wire [15:0] _02593_;
  wire [31:0] _02594_;
  wire [31:0] _02595_;
  wire _02596_;
  wire _02597_;
  wire [31:0] _02598_;
  wire [4:0] _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire [31:0] _02605_;
  wire [3:0] _02606_;
  wire _02607_;
  wire [31:0] _02608_;
  wire [3:0] _02609_;
  wire [31:0] _02610_;
  wire _02611_;
  wire [31:0] _02612_;
  wire [3:0] _02613_;
  wire _02614_;
  wire _02615_;
  wire [31:0] _02616_;
  wire [4:0] _02617_;
  wire [2:0] _02618_;
  wire [2:0] _02619_;
  wire [2:0] _02620_;
  wire [2:0] _02621_;
  wire [2:0] _02622_;
  wire [31:0] _02623_;
  wire [4:0] _02624_;
  wire [31:0] _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire [3:0] _02643_;
  wire [4:0] _02644_;
  wire [7:0] _02645_;
  wire [7:0] _02646_;
  wire [7:0] _02647_;
  wire [7:0] _02648_;
  wire [7:0] _02649_;
  wire [7:0] _02650_;
  wire [7:0] _02651_;
  wire [7:0] _02652_;
  wire [7:0] _02653_;
  wire [7:0] _02654_;
  wire [7:0] _02655_;
  wire [7:0] _02656_;
  wire [7:0] _02657_;
  wire [7:0] _02658_;
  wire [7:0] _02659_;
  wire [7:0] _02660_;
  wire [2:0] _02661_;
  wire [223:0] _02662_;
  wire [223:0] _02663_;
  wire [6:0] _02664_;
  wire [31:0] _02665_;
  wire [34:0] _02666_;
  wire [34:0] _02667_;
  wire [6:0] _02668_;
  wire [4:0] _02669_;
  wire [95:0] _02670_;
  wire [95:0] _02671_;
  wire [2:0] _02672_;
  wire [31:0] _02673_;
  wire [159:0] _02674_;
  wire [159:0] _02675_;
  wire [4:0] _02676_;
  wire [31:0] _02677_;
  wire [95:0] _02678_;
  wire [95:0] _02679_;
  wire [2:0] _02680_;
  wire [31:0] _02681_;
  wire [127:0] _02682_;
  wire [127:0] _02683_;
  wire [31:0] _02684_;
  wire [44:0] _02685_;
  wire [44:0] _02686_;
  wire [2:0] _02687_;
  wire [14:0] _02688_;
  wire [47:0] _02689_;
  wire [47:0] _02690_;
  wire [15:0] _02691_;
  wire [95:0] _02692_;
  wire [95:0] _02693_;
  wire [2:0] _02694_;
  wire [31:0] _02695_;
  wire [7:0] _02696_;
  wire [7:0] _02697_;
  wire [1:0] _02698_;
  wire [3:0] _02699_;
  wire [3:0] _02700_;
  wire [15:0] _02701_;
  wire [3:0] _02702_;
  wire [3:0] _02703_;
  wire [3:0] _02704_;
  wire [15:0] _02705_;
  wire [15:0] _02706_;
  wire [15:0] _02707_;
  wire [15:0] _02708_;
  wire [15:0] _02709_;
  wire [15:0] _02710_;
  wire [15:0] _02711_;
  wire [15:0] _02712_;
  wire [31:0] _02713_;
  wire [31:0] _02714_;
  wire [31:0] _02715_;
  wire [5:0] _02716_;
  wire [5:0] _02717_;
  wire [5:0] _02718_;
  wire [5:0] _02719_;
  wire [5:0] _02720_;
  wire _02721_;
  wire _02722_;
  wire [7:0] _02723_;
  wire [7:0] _02724_;
  wire [7:0] _02725_;
  wire [5:0] _02726_;
  wire _02727_;
  wire _02728_;
  wire [5:0] _02729_;
  wire _02730_;
  wire _02731_;
  wire [31:0] _02732_;
  wire [31:0] _02733_;
  wire [31:0] _02734_;
  wire [4:0] _02735_;
  wire [4:0] _02736_;
  wire [4:0] _02737_;
  wire [4:0] _02738_;
  wire [5:0] _02739_;
  wire [5:0] _02740_;
  wire [5:0] _02741_;
  wire [5:0] _02742_;
  wire [31:0] _02743_;
  wire [31:0] _02744_;
  wire [31:0] _02745_;
  wire [5:0] _02746_;
  wire [5:0] _02747_;
  wire [5:0] _02748_;
  wire [5:0] _02749_;
  wire [4:0] _02750_;
  wire [4:0] _02751_;
  wire _02752_;
  wire _02753_;
  wire [7:0] _02754_;
  wire [7:0] _02755_;
  wire [7:0] _02756_;
  wire [7:0] _02757_;
  wire [7:0] _02758_;
  wire [7:0] _02759_;
  wire [15:0] _02760_;
  wire [15:0] _02761_;
  wire [15:0] _02762_;
  wire [15:0] _02763_;
  wire [15:0] _02764_;
  wire [15:0] _02765_;
  wire [15:0] _02766_;
  wire [15:0] _02767_;
  wire [15:0] _02768_;
  wire [15:0] _02769_;
  wire [15:0] _02770_;
  wire [15:0] _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire [30:0] _02778_;
  wire [4:0] _02779_;
  wire [3:0] _02780_;
  wire _02781_;
  wire [15:0] _02782_;
  wire [15:0] _02783_;
  wire [15:0] _02784_;
  wire [3:0] _02785_;
  wire _02786_;
  wire [7:0] _02787_;
  wire [7:0] _02788_;
  wire [7:0] _02789_;
  wire [3:0] _02790_;
  wire [3:0] _02791_;
  wire _02792_;
  wire [29:0] _02793_;
  wire [29:0] _02794_;
  wire [29:0] _02795_;
  wire [29:0] _02796_;
  wire [30:0] _02797_;
  wire [31:0] _02798_;
  wire [5:0] _02799_;
  wire [5:0] _02800_;
  wire [30:0] _02801_;
  wire [31:0] _02802_;
  wire [31:0] _02803_;
  wire [31:0] _02804_;
  wire [31:0] _02805_;
  wire [31:0] _02806_;
  wire [31:0] _02807_;
  wire [31:0] _02808_;
  wire [31:0] _02809_;
  wire [31:0] _02810_;
  wire [31:0] _02811_;
  wire [2:0] _02812_;
  wire [4:0] _02813_;
  wire [8:0] _02814_;
  wire [8:0] _02815_;
  wire [8:0] _02816_;
  wire [3:0] _02817_;
  wire [3:0] _02818_;
  wire [4:0] _02819_;
  wire [4:0] _02820_;
  wire [30:0] _02821_;
  wire [30:0] _02822_;
  wire _02823_;
  wire [15:0] _02824_;
  wire [15:0] _02825_;
  wire [15:0] _02826_;
  wire [31:0] _02827_;
  wire [31:0] _02828_;
  wire [1:0] _02829_;
  wire [2:0] _02830_;
  wire [2:0] _02831_;
  wire [31:0] _02832_;
  wire [31:0] _02833_;
  wire [31:0] _02834_;
  wire [511:0] _02835_;
  wire [511:0] _02836_;
  wire [255:0] _02837_;
  wire [255:0] _02838_;
  wire [63:0] _02839_;
  wire [127:0] _02840_;
  wire [127:0] _02841_;
  wire [127:0] _02842_;
  wire [127:0] _02843_;
  wire [127:0] _02844_;
  wire [127:0] _02845_;
  wire [127:0] _02846_;
  wire [127:0] _02847_;
  wire [127:0] _02848_;
  wire [127:0] _02849_;
  wire [127:0] _02850_;
  wire [511:0] _02851_;
  wire [511:0] _02852_;
  wire [511:0] _02853_;
  wire [511:0] _02854_;
  wire [511:0] _02855_;
  wire [511:0] _02856_;
  wire [63:0] _02857_;
  wire [63:0] _02858_;
  wire [63:0] _02859_;
  wire [63:0] _02860_;
  wire [1023:0] _02861_;
  wire [1023:0] _02862_;
  wire [1023:0] _02863_;
  wire [127:0] _02864_;
  wire [127:0] _02865_;
  wire [127:0] _02866_;
  wire [127:0] _02867_;
  wire [127:0] _02868_;
  wire [127:0] _02869_;
  wire [127:0] _02870_;
  wire [127:0] _02871_;
  wire [127:0] _02872_;
  wire [127:0] _02873_;
  wire [127:0] _02874_;
  wire [127:0] _02875_;
  wire [127:0] _02876_;
  wire [127:0] _02877_;
  wire [127:0] _02878_;
  wire [127:0] _02879_;
  wire [127:0] _02880_;
  wire [127:0] _02881_;
  wire [127:0] _02882_;
  wire [127:0] _02883_;
  wire [127:0] _02884_;
  wire [127:0] _02885_;
  wire [127:0] _02886_;
  wire [127:0] _02887_;
  wire [127:0] _02888_;
  wire [127:0] _02889_;
  wire [127:0] _02890_;
  wire [127:0] _02891_;
  wire [127:0] _02892_;
  wire [127:0] _02893_;
  wire [127:0] _02894_;
  wire [127:0] _02895_;
  wire [127:0] _02896_;
  wire [127:0] _02897_;
  wire [127:0] _02898_;
  wire [127:0] _02899_;
  wire [127:0] _02900_;
  wire [127:0] _02901_;
  wire [127:0] _02902_;
  wire [127:0] _02903_;
  wire [127:0] _02904_;
  wire [127:0] _02905_;
  wire [127:0] _02906_;
  wire [127:0] _02907_;
  wire [127:0] _02908_;
  wire [127:0] _02909_;
  wire [127:0] _02910_;
  wire [127:0] _02911_;
  wire [127:0] _02912_;
  wire [127:0] _02913_;
  wire [127:0] _02914_;
  wire [127:0] _02915_;
  wire [127:0] _02916_;
  wire [127:0] _02917_;
  wire [1023:0] _02918_;
  wire [1023:0] _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire [5:0] _02930_;
  wire [5:0] _02931_;
  wire [5:0] _02932_;
  wire [5:0] _02933_;
  wire [8:0] _02934_;
  wire [8:0] _02935_;
  wire [32:0] _02936_;
  wire [32:0] _02937_;
  wire [32:0] _02938_;
  wire [32:0] _02939_;
  wire [32:0] _02940_;
  wire [5:0] _02941_;
  wire [5:0] _02942_;
  wire [5:0] _02943_;
  wire [5:0] _02944_;
  wire [32:0] _02945_;
  wire [32:0] _02946_;
  wire [32:0] _02947_;
  wire [32:0] _02948_;
  wire [32:0] _02949_;
  wire [15:0] _02950_;
  wire [15:0] _02951_;
  wire [15:0] _02952_;
  wire [15:0] _02953_;
  wire [15:0] _02954_;
  wire [15:0] _02955_;
  wire [15:0] _02956_;
  wire [15:0] _02957_;
  wire [31:0] _02958_;
  wire [31:0] _02959_;
  wire [31:0] _02960_;
  wire [5:0] _02961_;
  wire [5:0] _02962_;
  wire [5:0] _02963_;
  wire [5:0] _02964_;
  wire [5:0] _02965_;
  wire _02966_;
  wire _02967_;
  wire [7:0] _02968_;
  wire [7:0] _02969_;
  wire [7:0] _02970_;
  wire [5:0] _02971_;
  wire _02972_;
  wire _02973_;
  wire [5:0] _02974_;
  wire _02975_;
  wire _02976_;
  wire [31:0] _02977_;
  wire [31:0] _02978_;
  wire [31:0] _02979_;
  wire [4:0] _02980_;
  wire [4:0] _02981_;
  wire [4:0] _02982_;
  wire [4:0] _02983_;
  wire [5:0] _02984_;
  wire [5:0] _02985_;
  wire [5:0] _02986_;
  wire [5:0] _02987_;
  wire [31:0] _02988_;
  wire [31:0] _02989_;
  wire [31:0] _02990_;
  wire [5:0] _02991_;
  wire [5:0] _02992_;
  wire [5:0] _02993_;
  wire [5:0] _02994_;
  wire [4:0] _02995_;
  wire [4:0] _02996_;
  wire _02997_;
  wire _02998_;
  wire [7:0] _02999_;
  wire [7:0] _03000_;
  wire [7:0] _03001_;
  wire [7:0] _03002_;
  wire [7:0] _03003_;
  wire [7:0] _03004_;
  wire [15:0] _03005_;
  wire [15:0] _03006_;
  wire [15:0] _03007_;
  wire [15:0] _03008_;
  wire [15:0] _03009_;
  wire [15:0] _03010_;
  wire [15:0] _03011_;
  wire [15:0] _03012_;
  wire [15:0] _03013_;
  wire [15:0] _03014_;
  wire [15:0] _03015_;
  wire [15:0] _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire [30:0] _03023_;
  wire [4:0] _03024_;
  wire [3:0] _03025_;
  wire _03026_;
  wire [15:0] _03027_;
  wire [15:0] _03028_;
  wire [15:0] _03029_;
  wire [3:0] _03030_;
  wire _03031_;
  wire [7:0] _03032_;
  wire [7:0] _03033_;
  wire [7:0] _03034_;
  wire [3:0] _03035_;
  wire [3:0] _03036_;
  wire _03037_;
  wire [29:0] _03038_;
  wire [29:0] _03039_;
  wire [29:0] _03040_;
  wire [29:0] _03041_;
  wire [30:0] _03042_;
  wire [31:0] _03043_;
  wire [5:0] _03044_;
  wire [5:0] _03045_;
  wire [30:0] _03046_;
  wire [31:0] _03047_;
  wire [31:0] _03048_;
  wire [31:0] _03049_;
  wire [31:0] _03050_;
  wire [31:0] _03051_;
  wire [31:0] _03052_;
  wire [31:0] _03053_;
  wire [31:0] _03054_;
  wire [31:0] _03055_;
  wire [31:0] _03056_;
  wire [2:0] _03057_;
  wire [4:0] _03058_;
  wire [8:0] _03059_;
  wire [8:0] _03060_;
  wire [8:0] _03061_;
  wire [3:0] _03062_;
  wire [3:0] _03063_;
  wire [4:0] _03064_;
  wire [4:0] _03065_;
  wire [30:0] _03066_;
  wire [30:0] _03067_;
  wire _03068_;
  wire [15:0] _03069_;
  wire [15:0] _03070_;
  wire [15:0] _03071_;
  wire [31:0] _03072_;
  wire [31:0] _03073_;
  wire [1:0] _03074_;
  wire [2:0] _03075_;
  wire [2:0] _03076_;
  wire [31:0] _03077_;
  wire [31:0] _03078_;
  wire [31:0] _03079_;
  wire [511:0] _03080_;
  wire [511:0] _03081_;
  wire [255:0] _03082_;
  wire [255:0] _03083_;
  wire [63:0] _03084_;
  wire [127:0] _03085_;
  wire [127:0] _03086_;
  wire [127:0] _03087_;
  wire [127:0] _03088_;
  wire [127:0] _03089_;
  wire [127:0] _03090_;
  wire [127:0] _03091_;
  wire [127:0] _03092_;
  wire [127:0] _03093_;
  wire [127:0] _03094_;
  wire [127:0] _03095_;
  wire [511:0] _03096_;
  wire [511:0] _03097_;
  wire [511:0] _03098_;
  wire [511:0] _03099_;
  wire [511:0] _03100_;
  wire [511:0] _03101_;
  wire [63:0] _03102_;
  wire [63:0] _03103_;
  wire [63:0] _03104_;
  wire [63:0] _03105_;
  wire [1023:0] _03106_;
  wire [1023:0] _03107_;
  wire [1023:0] _03108_;
  wire [127:0] _03109_;
  wire [127:0] _03110_;
  wire [127:0] _03111_;
  wire [127:0] _03112_;
  wire [127:0] _03113_;
  wire [127:0] _03114_;
  wire [127:0] _03115_;
  wire [127:0] _03116_;
  wire [127:0] _03117_;
  wire [127:0] _03118_;
  wire [127:0] _03119_;
  wire [127:0] _03120_;
  wire [127:0] _03121_;
  wire [127:0] _03122_;
  wire [127:0] _03123_;
  wire [127:0] _03124_;
  wire [127:0] _03125_;
  wire [127:0] _03126_;
  wire [127:0] _03127_;
  wire [127:0] _03128_;
  wire [127:0] _03129_;
  wire [127:0] _03130_;
  wire [127:0] _03131_;
  wire [127:0] _03132_;
  wire [127:0] _03133_;
  wire [127:0] _03134_;
  wire [127:0] _03135_;
  wire [127:0] _03136_;
  wire [127:0] _03137_;
  wire [127:0] _03138_;
  wire [127:0] _03139_;
  wire [127:0] _03140_;
  wire [127:0] _03141_;
  wire [127:0] _03142_;
  wire [127:0] _03143_;
  wire [127:0] _03144_;
  wire [127:0] _03145_;
  wire [127:0] _03146_;
  wire [127:0] _03147_;
  wire [127:0] _03148_;
  wire [127:0] _03149_;
  wire [127:0] _03150_;
  wire [127:0] _03151_;
  wire [127:0] _03152_;
  wire [127:0] _03153_;
  wire [127:0] _03154_;
  wire [127:0] _03155_;
  wire [127:0] _03156_;
  wire [127:0] _03157_;
  wire [127:0] _03158_;
  wire [127:0] _03159_;
  wire [127:0] _03160_;
  wire [127:0] _03161_;
  wire [127:0] _03162_;
  wire [1023:0] _03163_;
  wire [1023:0] _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire [5:0] _03175_;
  wire [5:0] _03176_;
  wire [5:0] _03177_;
  wire [5:0] _03178_;
  wire [8:0] _03179_;
  wire [8:0] _03180_;
  wire [32:0] _03181_;
  wire [32:0] _03182_;
  wire [32:0] _03183_;
  wire [32:0] _03184_;
  wire [32:0] _03185_;
  wire [5:0] _03186_;
  wire [5:0] _03187_;
  wire [5:0] _03188_;
  wire [5:0] _03189_;
  wire [32:0] _03190_;
  wire [32:0] _03191_;
  wire [32:0] _03192_;
  wire [32:0] _03193_;
  wire [32:0] _03194_;
  wire [15:0] _03195_;
  wire [15:0] _03196_;
  wire [15:0] _03197_;
  wire [15:0] _03198_;
  wire [15:0] _03199_;
  wire [15:0] _03200_;
  wire [15:0] _03201_;
  wire [15:0] _03202_;
  wire [31:0] _03203_;
  wire [31:0] _03204_;
  wire [31:0] _03205_;
  wire [5:0] _03206_;
  wire [5:0] _03207_;
  wire [5:0] _03208_;
  wire [5:0] _03209_;
  wire [5:0] _03210_;
  wire _03211_;
  wire _03212_;
  wire [7:0] _03213_;
  wire [7:0] _03214_;
  wire [7:0] _03215_;
  wire [5:0] _03216_;
  wire _03217_;
  wire _03218_;
  wire [5:0] _03219_;
  wire _03220_;
  wire _03221_;
  wire [31:0] _03222_;
  wire [31:0] _03223_;
  wire [31:0] _03224_;
  wire [4:0] _03225_;
  wire [4:0] _03226_;
  wire [4:0] _03227_;
  wire [4:0] _03228_;
  wire [5:0] _03229_;
  wire [5:0] _03230_;
  wire [5:0] _03231_;
  wire [5:0] _03232_;
  wire [31:0] _03233_;
  wire [31:0] _03234_;
  wire [31:0] _03235_;
  wire [5:0] _03236_;
  wire [5:0] _03237_;
  wire [5:0] _03238_;
  wire [5:0] _03239_;
  wire [4:0] _03240_;
  wire [4:0] _03241_;
  wire _03242_;
  wire _03243_;
  wire [7:0] _03244_;
  wire [7:0] _03245_;
  wire [7:0] _03246_;
  wire [7:0] _03247_;
  wire [7:0] _03248_;
  wire [7:0] _03249_;
  wire [15:0] _03250_;
  wire [15:0] _03251_;
  wire [15:0] _03252_;
  wire [15:0] _03253_;
  wire [15:0] _03254_;
  wire [15:0] _03255_;
  wire [15:0] _03256_;
  wire [15:0] _03257_;
  wire [15:0] _03258_;
  wire [15:0] _03259_;
  wire [15:0] _03260_;
  wire [15:0] _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire [30:0] _03268_;
  wire [4:0] _03269_;
  wire [3:0] _03270_;
  wire _03271_;
  wire [15:0] _03272_;
  wire [15:0] _03273_;
  wire [15:0] _03274_;
  wire [3:0] _03275_;
  wire _03276_;
  wire [7:0] _03277_;
  wire [7:0] _03278_;
  wire [7:0] _03279_;
  wire [3:0] _03280_;
  wire [3:0] _03281_;
  wire _03282_;
  wire [29:0] _03283_;
  wire [29:0] _03284_;
  wire [29:0] _03285_;
  wire [29:0] _03286_;
  wire [30:0] _03287_;
  wire [31:0] _03288_;
  wire [5:0] _03289_;
  wire [5:0] _03290_;
  wire [30:0] _03291_;
  wire [31:0] _03292_;
  wire [31:0] _03293_;
  wire [31:0] _03294_;
  wire [31:0] _03295_;
  wire [31:0] _03296_;
  wire [31:0] _03297_;
  wire [31:0] _03298_;
  wire [31:0] _03299_;
  wire [31:0] _03300_;
  wire [31:0] _03301_;
  wire [2:0] _03302_;
  wire [4:0] _03303_;
  wire [8:0] _03304_;
  wire [8:0] _03305_;
  wire [8:0] _03306_;
  wire [3:0] _03307_;
  wire [3:0] _03308_;
  wire [4:0] _03309_;
  wire [4:0] _03310_;
  wire [30:0] _03311_;
  wire [30:0] _03312_;
  wire _03313_;
  wire [15:0] _03314_;
  wire [15:0] _03315_;
  wire [15:0] _03316_;
  wire [31:0] _03317_;
  wire [31:0] _03318_;
  wire [1:0] _03319_;
  wire [2:0] _03320_;
  wire [2:0] _03321_;
  wire [31:0] _03322_;
  wire [31:0] _03323_;
  wire [31:0] _03324_;
  wire [511:0] _03325_;
  wire [511:0] _03326_;
  wire [255:0] _03327_;
  wire [255:0] _03328_;
  wire [63:0] _03329_;
  wire [127:0] _03330_;
  wire [127:0] _03331_;
  wire [127:0] _03332_;
  wire [127:0] _03333_;
  wire [127:0] _03334_;
  wire [127:0] _03335_;
  wire [127:0] _03336_;
  wire [127:0] _03337_;
  wire [127:0] _03338_;
  wire [127:0] _03339_;
  wire [127:0] _03340_;
  wire [511:0] _03341_;
  wire [511:0] _03342_;
  wire [511:0] _03343_;
  wire [511:0] _03344_;
  wire [511:0] _03345_;
  wire [511:0] _03346_;
  wire [63:0] _03347_;
  wire [63:0] _03348_;
  wire [63:0] _03349_;
  wire [63:0] _03350_;
  wire [1023:0] _03351_;
  wire [1023:0] _03352_;
  wire [1023:0] _03353_;
  wire [127:0] _03354_;
  wire [127:0] _03355_;
  wire [127:0] _03356_;
  wire [127:0] _03357_;
  wire [127:0] _03358_;
  wire [127:0] _03359_;
  wire [127:0] _03360_;
  wire [127:0] _03361_;
  wire [127:0] _03362_;
  wire [127:0] _03363_;
  wire [127:0] _03364_;
  wire [127:0] _03365_;
  wire [127:0] _03366_;
  wire [127:0] _03367_;
  wire [127:0] _03368_;
  wire [127:0] _03369_;
  wire [127:0] _03370_;
  wire [127:0] _03371_;
  wire [127:0] _03372_;
  wire [127:0] _03373_;
  wire [127:0] _03374_;
  wire [127:0] _03375_;
  wire [127:0] _03376_;
  wire [127:0] _03377_;
  wire [127:0] _03378_;
  wire [127:0] _03379_;
  wire [127:0] _03380_;
  wire [127:0] _03381_;
  wire [127:0] _03382_;
  wire [127:0] _03383_;
  wire [127:0] _03384_;
  wire [127:0] _03385_;
  wire [127:0] _03386_;
  wire [127:0] _03387_;
  wire [127:0] _03388_;
  wire [127:0] _03389_;
  wire [127:0] _03390_;
  wire [127:0] _03391_;
  wire [127:0] _03392_;
  wire [127:0] _03393_;
  wire [127:0] _03394_;
  wire [127:0] _03395_;
  wire [127:0] _03396_;
  wire [127:0] _03397_;
  wire [127:0] _03398_;
  wire [127:0] _03399_;
  wire [127:0] _03400_;
  wire [127:0] _03401_;
  wire [127:0] _03402_;
  wire [127:0] _03403_;
  wire [127:0] _03404_;
  wire [127:0] _03405_;
  wire [127:0] _03406_;
  wire [127:0] _03407_;
  wire [1023:0] _03408_;
  wire [1023:0] _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire [5:0] _03420_;
  wire [5:0] _03421_;
  wire [5:0] _03422_;
  wire [5:0] _03423_;
  wire [8:0] _03424_;
  wire [8:0] _03425_;
  wire [32:0] _03426_;
  wire [32:0] _03427_;
  wire [32:0] _03428_;
  wire [32:0] _03429_;
  wire [32:0] _03430_;
  wire [5:0] _03431_;
  wire [5:0] _03432_;
  wire [5:0] _03433_;
  wire [5:0] _03434_;
  wire [32:0] _03435_;
  wire [32:0] _03436_;
  wire [32:0] _03437_;
  wire [32:0] _03438_;
  wire [32:0] _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire [29:0] _05712_;
  wire [29:0] _05713_;
  wire _05714_;
  wire [29:0] _05715_;
  wire _05716_;
  wire [29:0] _05717_;
  wire [29:0] _05718_;
  wire _05719_;
  wire [31:0] _05720_;
  wire [31:0] _05721_;
  wire [31:0] _05722_;
  wire _05723_;
  wire [31:0] _05724_;
  wire [31:0] _05725_;
  wire [31:0] _05726_;
  wire _05727_;
  wire [31:0] _05728_;
  wire [31:0] _05729_;
  wire [31:0] _05730_;
  wire _05731_;
  wire [31:0] _05732_;
  wire [31:0] _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire P1_BS16_n;
  wire P1_CLOCK;
  wire [31:0] P1_DataWidth;
  wire [31:0] P1_Datai;
  wire P1_HOLD;
  wire P1_NA_n;
  wire P1_READY_n;
  wire P1_RESET;
  wire P2_BS16_n;
  wire P2_CLOCK;
  wire [31:0] P2_DataWidth;
  wire [31:0] P2_Datai;
  wire P2_HOLD;
  wire P2_NA_n;
  wire P2_READY_n;
  wire P2_RESET;
  wire P3_BS16_n;
  wire P3_CLOCK;
  wire [31:0] P3_DataWidth;
  wire [31:0] P3_Datai;
  wire P3_HOLD;
  wire P3_NA_n;
  wire P3_READY_n;
  wire P3_RESET;
  wire [29:0] addr1;
  wire [29:0] addr2;
  wire [29:0] addr3;
  output [29:0] address1;
  output [29:0] address2;
  wire ads1;
  wire ads2;
  wire ads3;
  output ast1;
  output ast2;
  wire [3:0] be1;
  wire [3:0] be2;
  wire [3:0] be3;
  input bs16;
  input clock;
  input [31:0] datai;
  output [31:0] datao;
  output dc;
  wire dc1;
  wire dc2;
  wire dc3;
  wire [31:0] di1;
  wire [31:0] di2;
  wire [31:0] di3;
  wire [31:0] do1;
  wire [31:0] do2;
  wire [31:0] do3;
  input hold;
  output mio;
  wire mio1;
  wire mio2;
  wire mio3;
  input na;
  wire rdy1;
  wire rdy2;
  wire rdy3;
  input ready1;
  input ready2;
  input reset;
  output wr;
  wire wr1;
  wire wr2;
  wire wr3;
  INV_X1 U0 ( .A(P1_P1_State2_PTR3), .ZN(_00296_) );
  INV_X1 U1 ( .A(P1_P1_State2_PTR1), .ZN(_00297_) );
  INV_X1 U2 ( .A(P2_P1_State2_PTR1), .ZN(_00295_) );
  INV_X1 U3 ( .A(P2_P1_State2_PTR3), .ZN(_00294_) );
  INV_X1 U4 ( .A(P3_State_PTR0), .ZN(_00306_) );
  INV_X1 U5 ( .A(P2_State_PTR0), .ZN(_00305_) );
  INV_X1 U6 ( .A(P1_State_PTR0), .ZN(_00311_) );
  DFFR_X1 P3_State_PTR2 ( .D(_02459__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_State_PTR2), .QN());
  DFFR_X1 P3_StateBS16 ( .D(_02427_), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_StateBS16), .QN());
  DFFR_X1 P3_RequestPending ( .D(_03258__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_RequestPending), .QN());
  DFFR_X1 P3_ReadRequest ( .D(_03252__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_ReadRequest), .QN());
  DFFR_X1 P3_P1_uWord_PTR14 ( .D(_02517__PTR94), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR14), .QN());
  DFFR_X1 P3_P1_lWord_PTR15 ( .D(_02518__PTR95), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR15), .QN());
  DFFR_X1 P3_P1_State2_PTR3 ( .D(_02476__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_State2_PTR3), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR31 ( .D(_03343__PTR31), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR31), .QN());
  DFFR_X1 P3_P1_More ( .D(_02434__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_More), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR8_PTR7 ( .D(_02494__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR8_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR9_PTR7 ( .D(_02492__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR9_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR10_PTR7 ( .D(_02490__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR10_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR11_PTR7 ( .D(_02488__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR11_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR12_PTR7 ( .D(_02486__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR12_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR13_PTR7 ( .D(_02484__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR13_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR14_PTR7 ( .D(_02482__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR14_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR15_PTR7 ( .D(_02480__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR15_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR1_PTR7 ( .D(_02508__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR1_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR2_PTR7 ( .D(_02506__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR2_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR3_PTR7 ( .D(_02504__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR3_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR4_PTR7 ( .D(_02502__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR4_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR5_PTR7 ( .D(_02500__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR5_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR6_PTR7 ( .D(_02498__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR6_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR7_PTR7 ( .D(_02496__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR7_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR0_PTR7 ( .D(_02510__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR0_PTR7), .QN());
  DFFR_X1 P3_P1_InstQueueWr_Addr_PTR4 ( .D(_02512__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueueWr_Addr_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueueRd_Addr_PTR4 ( .D(_02514__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueueRd_Addr_PTR4), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR31 ( .D(_03346__PTR31), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR31), .QN());
  DFFR_X1 P3_P1_Flush ( .D(_02433__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_Flush), .QN());
  DFFR_X1 P3_MemoryFetch ( .D(_03255__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_MemoryFetch), .QN());
  DFFR_X1 P3_EBX_PTR31 ( .D(_02516__PTR191), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR31), .QN());
  DFFR_X1 P3_EAX_PTR31 ( .D(_02515__PTR191), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR31), .QN());
  DFFR_X1 P3_D_C_n ( .D(_02425_), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_D_C_n), .QN());
  DFFR_X1 P3_CodeFetch ( .D(_03261__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_CodeFetch), .QN());
  DFFR_X1 P3_Address_PTR29 ( .D(_02462__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR29), .QN());
  DFFR_X1 P3_ADS_n ( .D(_02426_), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_ADS_n), .QN());
  DFFR_X1 P2_State_PTR2 ( .D(_02170__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_State_PTR2), .QN());
  DFFR_X1 P2_StateBS16 ( .D(_02138_), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_StateBS16), .QN());
  DFFR_X1 P2_RequestPending ( .D(_03013__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_RequestPending), .QN());
  DFFR_X1 P2_ReadRequest ( .D(_03007__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_ReadRequest), .QN());
  DFFR_X1 P2_P1_uWord_PTR14 ( .D(_02228__PTR94), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR14), .QN());
  DFFR_X1 P2_P1_lWord_PTR15 ( .D(_02229__PTR95), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR15), .QN());
  DFFR_X1 P2_P1_State2_PTR3 ( .D(_02187__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_State2_PTR3), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR31 ( .D(_03098__PTR31), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR31), .QN());
  DFFR_X1 P2_P1_More ( .D(_02145__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_More), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR8_PTR7 ( .D(_02205__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR8_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR9_PTR7 ( .D(_02203__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR9_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR10_PTR7 ( .D(_02201__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR10_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR11_PTR7 ( .D(_02199__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR11_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR12_PTR7 ( .D(_02197__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR12_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR13_PTR7 ( .D(_02195__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR13_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR14_PTR7 ( .D(_02193__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR14_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR15_PTR7 ( .D(_02191__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR15_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR1_PTR7 ( .D(_02219__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR1_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR2_PTR7 ( .D(_02217__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR2_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR3_PTR7 ( .D(_02215__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR3_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR4_PTR7 ( .D(_02213__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR4_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR5_PTR7 ( .D(_02211__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR5_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR6_PTR7 ( .D(_02209__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR6_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR7_PTR7 ( .D(_02207__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR7_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR0_PTR7 ( .D(_02221__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR0_PTR7), .QN());
  DFFR_X1 P2_P1_InstQueueWr_Addr_PTR4 ( .D(_02223__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueueWr_Addr_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueueRd_Addr_PTR4 ( .D(_02225__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueueRd_Addr_PTR4), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR31 ( .D(_03101__PTR31), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR31), .QN());
  DFFR_X1 P2_P1_Flush ( .D(_02144__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_Flush), .QN());
  DFFR_X1 P2_MemoryFetch ( .D(_03010__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_MemoryFetch), .QN());
  DFFR_X1 P2_EBX_PTR31 ( .D(_02227__PTR191), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR31), .QN());
  DFFR_X1 P2_EAX_PTR31 ( .D(_02226__PTR191), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR31), .QN());
  DFFR_X1 P2_D_C_n ( .D(_02136_), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_D_C_n), .QN());
  DFFR_X1 P2_CodeFetch ( .D(_03016__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_CodeFetch), .QN());
  DFFR_X1 P2_Address_PTR29 ( .D(_02173__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR29), .QN());
  DFFR_X1 P2_ADS_n ( .D(_02137_), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_ADS_n), .QN());
  DFFR_X1 P1_State_PTR2 ( .D(_01877__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_State_PTR2), .QN());
  DFFR_X1 P1_StateBS16 ( .D(_01845_), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_StateBS16), .QN());
  DFFR_X1 P1_RequestPending ( .D(_02768__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_RequestPending), .QN());
  DFFR_X1 P1_ReadRequest ( .D(_02762__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_ReadRequest), .QN());
  DFFR_X1 P1_P1_uWord_PTR14 ( .D(_01936__PTR94), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR14), .QN());
  DFFR_X1 P1_P1_lWord_PTR15 ( .D(_01937__PTR95), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR15), .QN());
  DFFR_X1 P1_P1_State2_PTR3 ( .D(_01895__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_State2_PTR3), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR31 ( .D(_02853__PTR31), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR31), .QN());
  DFFR_X1 P1_P1_More ( .D(_01852__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_More), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR8_PTR7 ( .D(_01913__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR8_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR9_PTR7 ( .D(_01911__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR9_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR10_PTR7 ( .D(_01909__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR10_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR11_PTR7 ( .D(_01907__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR11_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR12_PTR7 ( .D(_01905__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR12_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR13_PTR7 ( .D(_01903__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR13_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR14_PTR7 ( .D(_01901__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR14_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR15_PTR7 ( .D(_01899__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR15_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR1_PTR7 ( .D(_01927__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR1_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR2_PTR7 ( .D(_01925__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR2_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR3_PTR7 ( .D(_01923__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR3_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR4_PTR7 ( .D(_01921__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR4_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR5_PTR7 ( .D(_01919__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR5_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR6_PTR7 ( .D(_01917__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR6_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR7_PTR7 ( .D(_01915__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR7_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR0_PTR7 ( .D(_01929__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR0_PTR7), .QN());
  DFFR_X1 P1_P1_InstQueueWr_Addr_PTR4 ( .D(_01931__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueueWr_Addr_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueueRd_Addr_PTR4 ( .D(_01933__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueueRd_Addr_PTR4), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR31 ( .D(_02856__PTR31), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR31), .QN());
  DFFR_X1 P1_P1_Flush ( .D(_01851__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_Flush), .QN());
  DFFR_X1 P1_MemoryFetch ( .D(_02765__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_MemoryFetch), .QN());
  DFFR_X1 P1_EBX_PTR31 ( .D(_01935__PTR191), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR31), .QN());
  DFFR_X1 P1_EAX_PTR31 ( .D(_01934__PTR191), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR31), .QN());
  DFFR_X1 P1_D_C_n ( .D(_01843_), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_D_C_n), .QN());
  DFFR_X1 P1_CodeFetch ( .D(_02771__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_CodeFetch), .QN());
  DFFR_X1 P1_Address_PTR29 ( .D(_01881__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR29), .QN());
  DFFR_X1 P1_ADS_n ( .D(_01844_), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_ADS_n), .QN());
  DFFR_X1 P1_rEIP_PTR0 ( .D(_01897__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR0), .QN());
  DFFR_X1 P1_rEIP_PTR1 ( .D(_01897__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR1), .QN());
  DFFR_X1 P1_rEIP_PTR2 ( .D(_01897__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR2), .QN());
  DFFR_X1 P1_rEIP_PTR3 ( .D(_01897__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR3), .QN());
  DFFR_X1 P1_rEIP_PTR4 ( .D(_01897__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR4), .QN());
  DFFR_X1 P1_rEIP_PTR5 ( .D(_01897__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR5), .QN());
  DFFR_X1 P1_rEIP_PTR6 ( .D(_01897__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR6), .QN());
  DFFR_X1 P1_rEIP_PTR7 ( .D(_01897__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR7), .QN());
  DFFR_X1 P1_rEIP_PTR8 ( .D(_01897__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR8), .QN());
  DFFR_X1 P1_rEIP_PTR9 ( .D(_01897__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR9), .QN());
  DFFR_X1 P1_rEIP_PTR10 ( .D(_01897__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR10), .QN());
  DFFR_X1 P1_rEIP_PTR11 ( .D(_01897__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR11), .QN());
  DFFR_X1 P1_rEIP_PTR12 ( .D(_01897__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR12), .QN());
  DFFR_X1 P1_rEIP_PTR13 ( .D(_01897__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR13), .QN());
  DFFR_X1 P1_rEIP_PTR14 ( .D(_01897__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR14), .QN());
  DFFR_X1 P1_rEIP_PTR15 ( .D(_01897__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR15), .QN());
  DFFR_X1 P1_rEIP_PTR16 ( .D(_01897__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR16), .QN());
  DFFR_X1 P1_rEIP_PTR17 ( .D(_01897__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR17), .QN());
  DFFR_X1 P1_rEIP_PTR18 ( .D(_01897__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR18), .QN());
  DFFR_X1 P1_rEIP_PTR19 ( .D(_01897__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR19), .QN());
  DFFR_X1 P1_rEIP_PTR20 ( .D(_01897__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR20), .QN());
  DFFR_X1 P1_rEIP_PTR21 ( .D(_01897__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR21), .QN());
  DFFR_X1 P1_rEIP_PTR22 ( .D(_01897__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR22), .QN());
  DFFR_X1 P1_rEIP_PTR23 ( .D(_01897__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR23), .QN());
  DFFR_X1 P1_rEIP_PTR24 ( .D(_01897__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR24), .QN());
  DFFR_X1 P1_rEIP_PTR25 ( .D(_01897__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR25), .QN());
  DFFR_X1 P1_rEIP_PTR26 ( .D(_01897__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR26), .QN());
  DFFR_X1 P1_rEIP_PTR27 ( .D(_01897__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR27), .QN());
  DFFR_X1 P1_rEIP_PTR28 ( .D(_01897__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR28), .QN());
  DFFR_X1 P1_rEIP_PTR29 ( .D(_01897__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR29), .QN());
  DFFR_X1 P1_rEIP_PTR30 ( .D(_01897__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR30), .QN());
  DFFR_X1 P1_EBX_PTR0 ( .D(_01935__PTR160), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR0), .QN());
  DFFR_X1 P1_EBX_PTR1 ( .D(_01935__PTR161), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR1), .QN());
  DFFR_X1 P1_EBX_PTR2 ( .D(_01935__PTR162), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR2), .QN());
  DFFR_X1 P1_EBX_PTR3 ( .D(_01935__PTR163), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR3), .QN());
  DFFR_X1 P1_EBX_PTR4 ( .D(_01935__PTR164), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR4), .QN());
  DFFR_X1 P1_EBX_PTR5 ( .D(_01935__PTR165), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR5), .QN());
  DFFR_X1 P1_EBX_PTR6 ( .D(_01935__PTR166), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR6), .QN());
  DFFR_X1 P1_EBX_PTR7 ( .D(_01935__PTR167), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR7), .QN());
  DFFR_X1 P1_EBX_PTR8 ( .D(_01935__PTR168), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR8), .QN());
  DFFR_X1 P1_EBX_PTR9 ( .D(_01935__PTR169), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR9), .QN());
  DFFR_X1 P1_EBX_PTR10 ( .D(_01935__PTR170), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR10), .QN());
  DFFR_X1 P1_EBX_PTR11 ( .D(_01935__PTR171), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR11), .QN());
  DFFR_X1 P1_EBX_PTR12 ( .D(_01935__PTR172), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR12), .QN());
  DFFR_X1 P1_EBX_PTR13 ( .D(_01935__PTR173), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR13), .QN());
  DFFR_X1 P1_EBX_PTR14 ( .D(_01935__PTR174), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR14), .QN());
  DFFR_X1 P1_EBX_PTR15 ( .D(_01935__PTR175), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR15), .QN());
  DFFR_X1 P1_EBX_PTR16 ( .D(_01935__PTR176), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR16), .QN());
  DFFR_X1 P1_EBX_PTR17 ( .D(_01935__PTR177), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR17), .QN());
  DFFR_X1 P1_EBX_PTR18 ( .D(_01935__PTR178), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR18), .QN());
  DFFR_X1 P1_EBX_PTR19 ( .D(_01935__PTR179), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR19), .QN());
  DFFR_X1 P1_EBX_PTR20 ( .D(_01935__PTR180), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR20), .QN());
  DFFR_X1 P1_EBX_PTR21 ( .D(_01935__PTR181), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR21), .QN());
  DFFR_X1 P1_EBX_PTR22 ( .D(_01935__PTR182), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR22), .QN());
  DFFR_X1 P1_EBX_PTR23 ( .D(_01935__PTR183), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR23), .QN());
  DFFR_X1 P1_EBX_PTR24 ( .D(_01935__PTR184), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR24), .QN());
  DFFR_X1 P1_EBX_PTR25 ( .D(_01935__PTR185), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR25), .QN());
  DFFR_X1 P1_EBX_PTR26 ( .D(_01935__PTR186), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR26), .QN());
  DFFR_X1 P1_EBX_PTR27 ( .D(_01935__PTR187), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR27), .QN());
  DFFR_X1 P1_EBX_PTR28 ( .D(_01935__PTR188), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR28), .QN());
  DFFR_X1 P1_EBX_PTR29 ( .D(_01935__PTR189), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR29), .QN());
  DFFR_X1 P1_EBX_PTR30 ( .D(_01935__PTR190), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EBX_PTR30), .QN());
  DFFR_X1 P1_EAX_PTR0 ( .D(_01934__PTR160), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR0), .QN());
  DFFR_X1 P1_EAX_PTR1 ( .D(_01934__PTR161), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR1), .QN());
  DFFR_X1 P1_EAX_PTR2 ( .D(_01934__PTR162), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR2), .QN());
  DFFR_X1 P1_EAX_PTR3 ( .D(_01934__PTR163), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR3), .QN());
  DFFR_X1 P1_EAX_PTR4 ( .D(_01934__PTR164), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR4), .QN());
  DFFR_X1 P1_EAX_PTR5 ( .D(_01934__PTR165), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR5), .QN());
  DFFR_X1 P1_EAX_PTR6 ( .D(_01934__PTR166), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR6), .QN());
  DFFR_X1 P1_EAX_PTR7 ( .D(_01934__PTR167), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR7), .QN());
  DFFR_X1 P1_EAX_PTR8 ( .D(_01934__PTR168), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR8), .QN());
  DFFR_X1 P1_EAX_PTR9 ( .D(_01934__PTR169), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR9), .QN());
  DFFR_X1 P1_EAX_PTR10 ( .D(_01934__PTR170), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR10), .QN());
  DFFR_X1 P1_EAX_PTR11 ( .D(_01934__PTR171), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR11), .QN());
  DFFR_X1 P1_EAX_PTR12 ( .D(_01934__PTR172), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR12), .QN());
  DFFR_X1 P1_EAX_PTR13 ( .D(_01934__PTR173), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR13), .QN());
  DFFR_X1 P1_EAX_PTR14 ( .D(_01934__PTR174), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR14), .QN());
  DFFR_X1 P1_EAX_PTR15 ( .D(_01934__PTR175), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR15), .QN());
  DFFR_X1 P1_EAX_PTR16 ( .D(_01934__PTR176), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR16), .QN());
  DFFR_X1 P1_EAX_PTR17 ( .D(_01934__PTR177), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR17), .QN());
  DFFR_X1 P1_EAX_PTR18 ( .D(_01934__PTR178), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR18), .QN());
  DFFR_X1 P1_EAX_PTR19 ( .D(_01934__PTR179), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR19), .QN());
  DFFR_X1 P1_EAX_PTR20 ( .D(_01934__PTR180), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR20), .QN());
  DFFR_X1 P1_EAX_PTR21 ( .D(_01934__PTR181), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR21), .QN());
  DFFR_X1 P1_EAX_PTR22 ( .D(_01934__PTR182), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR22), .QN());
  DFFR_X1 P1_EAX_PTR23 ( .D(_01934__PTR183), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR23), .QN());
  DFFR_X1 P1_EAX_PTR24 ( .D(_01934__PTR184), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR24), .QN());
  DFFR_X1 P1_EAX_PTR25 ( .D(_01934__PTR185), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR25), .QN());
  DFFR_X1 P1_EAX_PTR26 ( .D(_01934__PTR186), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR26), .QN());
  DFFR_X1 P1_EAX_PTR27 ( .D(_01934__PTR187), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR27), .QN());
  DFFR_X1 P1_EAX_PTR28 ( .D(_01934__PTR188), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR28), .QN());
  DFFR_X1 P1_EAX_PTR29 ( .D(_01934__PTR189), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR29), .QN());
  DFFR_X1 P1_EAX_PTR30 ( .D(_01934__PTR190), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_EAX_PTR30), .QN());
  DFFR_X1 P1_Datao_PTR0 ( .D(_02919__PTR256), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR0), .QN());
  DFFR_X1 P1_Datao_PTR1 ( .D(_02919__PTR257), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR1), .QN());
  DFFR_X1 P1_Datao_PTR2 ( .D(_02919__PTR258), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR2), .QN());
  DFFR_X1 P1_Datao_PTR3 ( .D(_02919__PTR259), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR3), .QN());
  DFFR_X1 P1_Datao_PTR4 ( .D(_02919__PTR260), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR4), .QN());
  DFFR_X1 P1_Datao_PTR5 ( .D(_02919__PTR261), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR5), .QN());
  DFFR_X1 P1_Datao_PTR6 ( .D(_02919__PTR262), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR6), .QN());
  DFFR_X1 P1_Datao_PTR7 ( .D(_02919__PTR263), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR7), .QN());
  DFFR_X1 P1_Datao_PTR8 ( .D(_02919__PTR264), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR8), .QN());
  DFFR_X1 P1_Datao_PTR9 ( .D(_02919__PTR265), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR9), .QN());
  DFFR_X1 P1_Datao_PTR10 ( .D(_02919__PTR266), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR10), .QN());
  DFFR_X1 P1_Datao_PTR11 ( .D(_02919__PTR267), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR11), .QN());
  DFFR_X1 P1_Datao_PTR12 ( .D(_02919__PTR268), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR12), .QN());
  DFFR_X1 P1_Datao_PTR13 ( .D(_02919__PTR269), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR13), .QN());
  DFFR_X1 P1_Datao_PTR14 ( .D(_02919__PTR270), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR14), .QN());
  DFFR_X1 P1_Datao_PTR15 ( .D(_02919__PTR271), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR15), .QN());
  DFFR_X1 P1_Datao_PTR16 ( .D(_02919__PTR272), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR16), .QN());
  DFFR_X1 P1_Datao_PTR17 ( .D(_02919__PTR273), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR17), .QN());
  DFFR_X1 P1_Datao_PTR18 ( .D(_02919__PTR274), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR18), .QN());
  DFFR_X1 P1_Datao_PTR19 ( .D(_02919__PTR275), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR19), .QN());
  DFFR_X1 P1_Datao_PTR20 ( .D(_02919__PTR276), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR20), .QN());
  DFFR_X1 P1_Datao_PTR21 ( .D(_02919__PTR277), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR21), .QN());
  DFFR_X1 P1_Datao_PTR22 ( .D(_02919__PTR278), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR22), .QN());
  DFFR_X1 P1_Datao_PTR23 ( .D(_02919__PTR279), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR23), .QN());
  DFFR_X1 P1_Datao_PTR24 ( .D(_02919__PTR280), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR24), .QN());
  DFFR_X1 P1_Datao_PTR25 ( .D(_02919__PTR281), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR25), .QN());
  DFFR_X1 P1_Datao_PTR26 ( .D(_02919__PTR282), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR26), .QN());
  DFFR_X1 P1_Datao_PTR27 ( .D(_02919__PTR283), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR27), .QN());
  DFFR_X1 P1_Datao_PTR28 ( .D(_02919__PTR284), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR28), .QN());
  DFFR_X1 P1_Datao_PTR29 ( .D(_02919__PTR285), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR29), .QN());
  DFFR_X1 P1_Datao_PTR30 ( .D(_02919__PTR286), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR30), .QN());
  DFFR_X1 P1_DataWidth_reg_PTR0 ( .D(_01879__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR0), .QN());
  BUF_X1 U7 ( .A(P1_DataWidth_reg_PTR0), .Z(P1_DataWidth_PTR0) );
  DFFR_X1 P1_DataWidth_reg_PTR2 ( .D(_01879__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR2), .QN());
  BUF_X1 U8 ( .A(P1_DataWidth_reg_PTR2), .Z(P1_DataWidth_PTR2) );
  DFFR_X1 P1_DataWidth_reg_PTR3 ( .D(_01879__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR3), .QN());
  BUF_X1 U9 ( .A(P1_DataWidth_reg_PTR3), .Z(P1_DataWidth_PTR3) );
  DFFR_X1 P1_DataWidth_reg_PTR4 ( .D(_01879__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR4), .QN());
  BUF_X1 U10 ( .A(P1_DataWidth_reg_PTR4), .Z(P1_DataWidth_PTR4) );
  DFFR_X1 P1_DataWidth_reg_PTR5 ( .D(_01879__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR5), .QN());
  BUF_X1 U11 ( .A(P1_DataWidth_reg_PTR5), .Z(P1_DataWidth_PTR5) );
  DFFR_X1 P1_DataWidth_reg_PTR6 ( .D(_01879__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR6), .QN());
  BUF_X1 U12 ( .A(P1_DataWidth_reg_PTR6), .Z(P1_DataWidth_PTR6) );
  DFFR_X1 P1_DataWidth_reg_PTR7 ( .D(_01879__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR7), .QN());
  BUF_X1 U13 ( .A(P1_DataWidth_reg_PTR7), .Z(P1_DataWidth_PTR7) );
  DFFR_X1 P1_DataWidth_reg_PTR8 ( .D(_01879__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR8), .QN());
  BUF_X1 U14 ( .A(P1_DataWidth_reg_PTR8), .Z(P1_DataWidth_PTR8) );
  DFFR_X1 P1_DataWidth_reg_PTR9 ( .D(_01879__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR9), .QN());
  BUF_X1 U15 ( .A(P1_DataWidth_reg_PTR9), .Z(P1_DataWidth_PTR9) );
  DFFR_X1 P1_DataWidth_reg_PTR10 ( .D(_01879__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR10), .QN());
  BUF_X1 U16 ( .A(P1_DataWidth_reg_PTR10), .Z(P1_DataWidth_PTR10) );
  DFFR_X1 P1_DataWidth_reg_PTR11 ( .D(_01879__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR11), .QN());
  BUF_X1 U17 ( .A(P1_DataWidth_reg_PTR11), .Z(P1_DataWidth_PTR11) );
  DFFR_X1 P1_DataWidth_reg_PTR12 ( .D(_01879__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR12), .QN());
  BUF_X1 U18 ( .A(P1_DataWidth_reg_PTR12), .Z(P1_DataWidth_PTR12) );
  DFFR_X1 P1_DataWidth_reg_PTR13 ( .D(_01879__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR13), .QN());
  BUF_X1 U19 ( .A(P1_DataWidth_reg_PTR13), .Z(P1_DataWidth_PTR13) );
  DFFR_X1 P1_DataWidth_reg_PTR14 ( .D(_01879__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR14), .QN());
  BUF_X1 U20 ( .A(P1_DataWidth_reg_PTR14), .Z(P1_DataWidth_PTR14) );
  DFFR_X1 P1_DataWidth_reg_PTR15 ( .D(_01879__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR15), .QN());
  BUF_X1 U21 ( .A(P1_DataWidth_reg_PTR15), .Z(P1_DataWidth_PTR15) );
  DFFR_X1 P1_DataWidth_reg_PTR16 ( .D(_01879__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR16), .QN());
  BUF_X1 U22 ( .A(P1_DataWidth_reg_PTR16), .Z(P1_DataWidth_PTR16) );
  DFFR_X1 P1_DataWidth_reg_PTR17 ( .D(_01879__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR17), .QN());
  BUF_X1 U23 ( .A(P1_DataWidth_reg_PTR17), .Z(P1_DataWidth_PTR17) );
  DFFR_X1 P1_DataWidth_reg_PTR18 ( .D(_01879__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR18), .QN());
  BUF_X1 U24 ( .A(P1_DataWidth_reg_PTR18), .Z(P1_DataWidth_PTR18) );
  DFFR_X1 P1_DataWidth_reg_PTR19 ( .D(_01879__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR19), .QN());
  BUF_X1 U25 ( .A(P1_DataWidth_reg_PTR19), .Z(P1_DataWidth_PTR19) );
  DFFR_X1 P1_DataWidth_reg_PTR20 ( .D(_01879__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR20), .QN());
  BUF_X1 U26 ( .A(P1_DataWidth_reg_PTR20), .Z(P1_DataWidth_PTR20) );
  DFFR_X1 P1_DataWidth_reg_PTR21 ( .D(_01879__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR21), .QN());
  BUF_X1 U27 ( .A(P1_DataWidth_reg_PTR21), .Z(P1_DataWidth_PTR21) );
  DFFR_X1 P1_DataWidth_reg_PTR22 ( .D(_01879__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR22), .QN());
  BUF_X1 U28 ( .A(P1_DataWidth_reg_PTR22), .Z(P1_DataWidth_PTR22) );
  DFFR_X1 P1_DataWidth_reg_PTR23 ( .D(_01879__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR23), .QN());
  BUF_X1 U29 ( .A(P1_DataWidth_reg_PTR23), .Z(P1_DataWidth_PTR23) );
  DFFR_X1 P1_DataWidth_reg_PTR24 ( .D(_01879__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR24), .QN());
  BUF_X1 U30 ( .A(P1_DataWidth_reg_PTR24), .Z(P1_DataWidth_PTR24) );
  DFFR_X1 P1_DataWidth_reg_PTR25 ( .D(_01879__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR25), .QN());
  BUF_X1 U31 ( .A(P1_DataWidth_reg_PTR25), .Z(P1_DataWidth_PTR25) );
  DFFR_X1 P1_DataWidth_reg_PTR26 ( .D(_01879__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR26), .QN());
  BUF_X1 U32 ( .A(P1_DataWidth_reg_PTR26), .Z(P1_DataWidth_PTR26) );
  DFFR_X1 P1_DataWidth_reg_PTR27 ( .D(_01879__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR27), .QN());
  BUF_X1 U33 ( .A(P1_DataWidth_reg_PTR27), .Z(P1_DataWidth_PTR27) );
  DFFR_X1 P1_DataWidth_reg_PTR28 ( .D(_01879__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR28), .QN());
  BUF_X1 U34 ( .A(P1_DataWidth_reg_PTR28), .Z(P1_DataWidth_PTR28) );
  DFFR_X1 P1_DataWidth_reg_PTR29 ( .D(_01879__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR29), .QN());
  BUF_X1 U35 ( .A(P1_DataWidth_reg_PTR29), .Z(P1_DataWidth_PTR29) );
  DFFR_X1 P1_DataWidth_reg_PTR30 ( .D(_01879__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR30), .QN());
  BUF_X1 U36 ( .A(P1_DataWidth_reg_PTR30), .Z(P1_DataWidth_PTR30) );
  DFFR_X1 P1_State_PTR0 ( .D(_01877__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_State_PTR0), .QN());
  DFFR_X1 P1_State_PTR1 ( .D(_01877__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_State_PTR1), .QN());
  DFFR_X1 P1_Address_PTR0 ( .D(_01881__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR0), .QN());
  DFFR_X1 P1_Address_PTR1 ( .D(_01881__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR1), .QN());
  DFFR_X1 P1_Address_PTR2 ( .D(_01881__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR2), .QN());
  DFFR_X1 P1_Address_PTR3 ( .D(_01881__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR3), .QN());
  DFFR_X1 P1_Address_PTR4 ( .D(_01881__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR4), .QN());
  DFFR_X1 P1_Address_PTR5 ( .D(_01881__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR5), .QN());
  DFFR_X1 P1_Address_PTR6 ( .D(_01881__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR6), .QN());
  DFFR_X1 P1_Address_PTR7 ( .D(_01881__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR7), .QN());
  DFFR_X1 P1_Address_PTR8 ( .D(_01881__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR8), .QN());
  DFFR_X1 P1_Address_PTR9 ( .D(_01881__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR9), .QN());
  DFFR_X1 P1_Address_PTR10 ( .D(_01881__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR10), .QN());
  DFFR_X1 P1_Address_PTR11 ( .D(_01881__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR11), .QN());
  DFFR_X1 P1_Address_PTR12 ( .D(_01881__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR12), .QN());
  DFFR_X1 P1_Address_PTR13 ( .D(_01881__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR13), .QN());
  DFFR_X1 P1_Address_PTR14 ( .D(_01881__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR14), .QN());
  DFFR_X1 P1_Address_PTR15 ( .D(_01881__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR15), .QN());
  DFFR_X1 P1_Address_PTR16 ( .D(_01881__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR16), .QN());
  DFFR_X1 P1_Address_PTR17 ( .D(_01881__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR17), .QN());
  DFFR_X1 P1_Address_PTR18 ( .D(_01881__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR18), .QN());
  DFFR_X1 P1_Address_PTR19 ( .D(_01881__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR19), .QN());
  DFFR_X1 P1_Address_PTR20 ( .D(_01881__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR20), .QN());
  DFFR_X1 P1_Address_PTR21 ( .D(_01881__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR21), .QN());
  DFFR_X1 P1_Address_PTR22 ( .D(_01881__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR22), .QN());
  DFFR_X1 P1_Address_PTR23 ( .D(_01881__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR23), .QN());
  DFFR_X1 P1_Address_PTR24 ( .D(_01881__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR24), .QN());
  DFFR_X1 P1_Address_PTR25 ( .D(_01881__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR25), .QN());
  DFFR_X1 P1_Address_PTR26 ( .D(_01881__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR26), .QN());
  DFFR_X1 P1_Address_PTR27 ( .D(_01881__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR27), .QN());
  DFFR_X1 P1_Address_PTR28 ( .D(_01881__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Address_PTR28), .QN());
  DFFR_X1 P1_P1_uWord_PTR0 ( .D(_01936__PTR80), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR0), .QN());
  DFFR_X1 P1_P1_uWord_PTR1 ( .D(_01936__PTR81), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR1), .QN());
  DFFR_X1 P1_P1_uWord_PTR2 ( .D(_01936__PTR82), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR2), .QN());
  DFFR_X1 P1_P1_uWord_PTR3 ( .D(_01936__PTR83), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR3), .QN());
  DFFR_X1 P1_P1_uWord_PTR4 ( .D(_01936__PTR84), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR4), .QN());
  DFFR_X1 P1_P1_uWord_PTR5 ( .D(_01936__PTR85), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR5), .QN());
  DFFR_X1 P1_P1_uWord_PTR6 ( .D(_01936__PTR86), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR6), .QN());
  DFFR_X1 P1_P1_uWord_PTR7 ( .D(_01936__PTR87), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR7), .QN());
  DFFR_X1 P1_P1_uWord_PTR8 ( .D(_01936__PTR88), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR8), .QN());
  DFFR_X1 P1_P1_uWord_PTR9 ( .D(_01936__PTR89), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR9), .QN());
  DFFR_X1 P1_P1_uWord_PTR10 ( .D(_01936__PTR90), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR10), .QN());
  DFFR_X1 P1_P1_uWord_PTR11 ( .D(_01936__PTR91), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR11), .QN());
  DFFR_X1 P1_P1_uWord_PTR12 ( .D(_01936__PTR92), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR12), .QN());
  DFFR_X1 P1_P1_uWord_PTR13 ( .D(_01936__PTR93), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_uWord_PTR13), .QN());
  DFFR_X1 P1_P1_lWord_PTR0 ( .D(_01937__PTR80), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR0), .QN());
  DFFR_X1 P1_P1_lWord_PTR1 ( .D(_01937__PTR81), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR1), .QN());
  DFFR_X1 P1_P1_lWord_PTR2 ( .D(_01937__PTR82), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR2), .QN());
  DFFR_X1 P1_P1_lWord_PTR3 ( .D(_01937__PTR83), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR3), .QN());
  DFFR_X1 P1_P1_lWord_PTR4 ( .D(_01937__PTR84), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR4), .QN());
  DFFR_X1 P1_P1_lWord_PTR5 ( .D(_01937__PTR85), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR5), .QN());
  DFFR_X1 P1_P1_lWord_PTR6 ( .D(_01937__PTR86), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR6), .QN());
  DFFR_X1 P1_P1_lWord_PTR7 ( .D(_01937__PTR87), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR7), .QN());
  DFFR_X1 P1_P1_lWord_PTR8 ( .D(_01937__PTR88), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR8), .QN());
  DFFR_X1 P1_P1_lWord_PTR9 ( .D(_01937__PTR89), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR9), .QN());
  DFFR_X1 P1_P1_lWord_PTR10 ( .D(_01937__PTR90), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR10), .QN());
  DFFR_X1 P1_P1_lWord_PTR11 ( .D(_01937__PTR91), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR11), .QN());
  DFFR_X1 P1_P1_lWord_PTR12 ( .D(_01937__PTR92), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR12), .QN());
  DFFR_X1 P1_P1_lWord_PTR13 ( .D(_01937__PTR93), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR13), .QN());
  DFFR_X1 P1_P1_lWord_PTR14 ( .D(_01937__PTR94), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_lWord_PTR14), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR0 ( .D(_02853__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR0), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR1 ( .D(_02853__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR1), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR2 ( .D(_02853__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR2), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR3 ( .D(_02853__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR3), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR4 ( .D(_02853__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR4), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR5 ( .D(_02853__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR5), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR6 ( .D(_02853__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR6), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR7 ( .D(_02853__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR7), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR8 ( .D(_02853__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR8), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR9 ( .D(_02853__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR9), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR10 ( .D(_02853__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR10), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR11 ( .D(_02853__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR11), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR12 ( .D(_02853__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR12), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR13 ( .D(_02853__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR13), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR14 ( .D(_02853__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR14), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR15 ( .D(_02853__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR15), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR16 ( .D(_02853__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR16), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR17 ( .D(_02853__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR17), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR18 ( .D(_02853__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR18), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR19 ( .D(_02853__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR19), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR20 ( .D(_02853__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR20), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR21 ( .D(_02853__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR21), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR22 ( .D(_02853__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR22), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR23 ( .D(_02853__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR23), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR24 ( .D(_02853__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR24), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR25 ( .D(_02853__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR25), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR26 ( .D(_02853__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR26), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR27 ( .D(_02853__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR27), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR28 ( .D(_02853__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR28), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR29 ( .D(_02853__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR29), .QN());
  DFFR_X1 P1_P1_PhyAddrPointer_PTR30 ( .D(_02853__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_PhyAddrPointer_PTR30), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR0 ( .D(_02856__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR0), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR1 ( .D(_02856__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR1), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR2 ( .D(_02856__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR2), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR3 ( .D(_02856__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR3), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR4 ( .D(_02856__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR4), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR5 ( .D(_02856__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR5), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR6 ( .D(_02856__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR6), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR7 ( .D(_02856__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR7), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR8 ( .D(_02856__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR8), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR9 ( .D(_02856__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR9), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR10 ( .D(_02856__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR10), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR11 ( .D(_02856__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR11), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR12 ( .D(_02856__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR12), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR13 ( .D(_02856__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR13), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR14 ( .D(_02856__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR14), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR15 ( .D(_02856__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR15), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR16 ( .D(_02856__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR16), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR17 ( .D(_02856__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR17), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR18 ( .D(_02856__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR18), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR19 ( .D(_02856__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR19), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR20 ( .D(_02856__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR20), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR21 ( .D(_02856__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR21), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR22 ( .D(_02856__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR22), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR23 ( .D(_02856__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR23), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR24 ( .D(_02856__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR24), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR25 ( .D(_02856__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR25), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR26 ( .D(_02856__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR26), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR27 ( .D(_02856__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR27), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR28 ( .D(_02856__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR28), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR29 ( .D(_02856__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR29), .QN());
  DFFR_X1 P1_P1_InstAddrPointer_PTR30 ( .D(_02856__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstAddrPointer_PTR30), .QN());
  DFFR_X1 P1_P1_InstQueueWr_Addr_PTR0 ( .D(_01931__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueueWr_Addr_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueueWr_Addr_PTR1 ( .D(_01931__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueueWr_Addr_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueueWr_Addr_PTR2 ( .D(_01931__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueueWr_Addr_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueueWr_Addr_PTR3 ( .D(_01931__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueueWr_Addr_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueueRd_Addr_PTR0 ( .D(_01933__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueueRd_Addr_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueueRd_Addr_PTR1 ( .D(_01933__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueueRd_Addr_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueueRd_Addr_PTR2 ( .D(_01933__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueueRd_Addr_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueueRd_Addr_PTR3 ( .D(_01933__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueueRd_Addr_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR0_PTR0 ( .D(_01929__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR0_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR0_PTR1 ( .D(_01929__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR0_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR0_PTR2 ( .D(_01929__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR0_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR0_PTR3 ( .D(_01929__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR0_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR0_PTR4 ( .D(_01929__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR0_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR0_PTR5 ( .D(_01929__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR0_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR0_PTR6 ( .D(_01929__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR0_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR1_PTR0 ( .D(_01927__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR1_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR1_PTR1 ( .D(_01927__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR1_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR1_PTR2 ( .D(_01927__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR1_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR1_PTR3 ( .D(_01927__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR1_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR1_PTR4 ( .D(_01927__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR1_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR1_PTR5 ( .D(_01927__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR1_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR1_PTR6 ( .D(_01927__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR1_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR2_PTR0 ( .D(_01925__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR2_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR2_PTR1 ( .D(_01925__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR2_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR2_PTR2 ( .D(_01925__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR2_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR2_PTR3 ( .D(_01925__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR2_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR2_PTR4 ( .D(_01925__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR2_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR2_PTR5 ( .D(_01925__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR2_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR2_PTR6 ( .D(_01925__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR2_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR3_PTR0 ( .D(_01923__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR3_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR3_PTR1 ( .D(_01923__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR3_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR3_PTR2 ( .D(_01923__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR3_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR3_PTR3 ( .D(_01923__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR3_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR3_PTR4 ( .D(_01923__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR3_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR3_PTR5 ( .D(_01923__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR3_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR3_PTR6 ( .D(_01923__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR3_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR4_PTR0 ( .D(_01921__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR4_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR4_PTR1 ( .D(_01921__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR4_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR4_PTR2 ( .D(_01921__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR4_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR4_PTR3 ( .D(_01921__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR4_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR4_PTR4 ( .D(_01921__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR4_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR4_PTR5 ( .D(_01921__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR4_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR4_PTR6 ( .D(_01921__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR4_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR5_PTR0 ( .D(_01919__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR5_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR5_PTR1 ( .D(_01919__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR5_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR5_PTR2 ( .D(_01919__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR5_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR5_PTR3 ( .D(_01919__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR5_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR5_PTR4 ( .D(_01919__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR5_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR5_PTR5 ( .D(_01919__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR5_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR5_PTR6 ( .D(_01919__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR5_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR6_PTR0 ( .D(_01917__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR6_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR6_PTR1 ( .D(_01917__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR6_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR6_PTR2 ( .D(_01917__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR6_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR6_PTR3 ( .D(_01917__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR6_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR6_PTR4 ( .D(_01917__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR6_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR6_PTR5 ( .D(_01917__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR6_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR6_PTR6 ( .D(_01917__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR6_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR7_PTR0 ( .D(_01915__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR7_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR7_PTR1 ( .D(_01915__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR7_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR7_PTR2 ( .D(_01915__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR7_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR7_PTR3 ( .D(_01915__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR7_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR7_PTR4 ( .D(_01915__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR7_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR7_PTR5 ( .D(_01915__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR7_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR7_PTR6 ( .D(_01915__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR7_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR8_PTR0 ( .D(_01913__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR8_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR8_PTR1 ( .D(_01913__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR8_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR8_PTR2 ( .D(_01913__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR8_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR8_PTR3 ( .D(_01913__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR8_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR8_PTR4 ( .D(_01913__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR8_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR8_PTR5 ( .D(_01913__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR8_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR8_PTR6 ( .D(_01913__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR8_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR9_PTR0 ( .D(_01911__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR9_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR9_PTR1 ( .D(_01911__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR9_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR9_PTR2 ( .D(_01911__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR9_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR9_PTR3 ( .D(_01911__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR9_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR9_PTR4 ( .D(_01911__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR9_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR9_PTR5 ( .D(_01911__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR9_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR9_PTR6 ( .D(_01911__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR9_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR10_PTR0 ( .D(_01909__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR10_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR10_PTR1 ( .D(_01909__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR10_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR10_PTR2 ( .D(_01909__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR10_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR10_PTR3 ( .D(_01909__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR10_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR10_PTR4 ( .D(_01909__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR10_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR10_PTR5 ( .D(_01909__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR10_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR10_PTR6 ( .D(_01909__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR10_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR11_PTR0 ( .D(_01907__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR11_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR11_PTR1 ( .D(_01907__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR11_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR11_PTR2 ( .D(_01907__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR11_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR11_PTR3 ( .D(_01907__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR11_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR11_PTR4 ( .D(_01907__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR11_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR11_PTR5 ( .D(_01907__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR11_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR11_PTR6 ( .D(_01907__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR11_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR12_PTR0 ( .D(_01905__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR12_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR12_PTR1 ( .D(_01905__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR12_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR12_PTR2 ( .D(_01905__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR12_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR12_PTR3 ( .D(_01905__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR12_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR12_PTR4 ( .D(_01905__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR12_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR12_PTR5 ( .D(_01905__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR12_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR12_PTR6 ( .D(_01905__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR12_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR13_PTR0 ( .D(_01903__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR13_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR13_PTR1 ( .D(_01903__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR13_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR13_PTR2 ( .D(_01903__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR13_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR13_PTR3 ( .D(_01903__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR13_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR13_PTR4 ( .D(_01903__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR13_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR13_PTR5 ( .D(_01903__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR13_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR13_PTR6 ( .D(_01903__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR13_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR14_PTR0 ( .D(_01901__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR14_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR14_PTR1 ( .D(_01901__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR14_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR14_PTR2 ( .D(_01901__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR14_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR14_PTR3 ( .D(_01901__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR14_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR14_PTR4 ( .D(_01901__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR14_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR14_PTR5 ( .D(_01901__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR14_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR14_PTR6 ( .D(_01901__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR14_PTR6), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR15_PTR0 ( .D(_01899__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR15_PTR0), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR15_PTR1 ( .D(_01899__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR15_PTR1), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR15_PTR2 ( .D(_01899__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR15_PTR2), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR15_PTR3 ( .D(_01899__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR15_PTR3), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR15_PTR4 ( .D(_01899__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR15_PTR4), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR15_PTR5 ( .D(_01899__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR15_PTR5), .QN());
  DFFR_X1 P1_P1_InstQueue_PTR15_PTR6 ( .D(_01899__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_InstQueue_PTR15_PTR6), .QN());
  DFFR_X1 P1_P1_State2_PTR0 ( .D(_01895__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_State2_PTR0), .QN());
  DFFR_X1 P1_P1_State2_PTR1 ( .D(_01895__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_State2_PTR1), .QN());
  DFFR_X1 P1_P1_State2_PTR2 ( .D(_01895__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_P1_State2_PTR2), .QN());
  DFFR_X1 P2_rEIP_PTR0 ( .D(_02189__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR0), .QN());
  DFFR_X1 P2_rEIP_PTR1 ( .D(_02189__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR1), .QN());
  DFFR_X1 P2_rEIP_PTR2 ( .D(_02189__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR2), .QN());
  DFFR_X1 P2_rEIP_PTR3 ( .D(_02189__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR3), .QN());
  DFFR_X1 P2_rEIP_PTR4 ( .D(_02189__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR4), .QN());
  DFFR_X1 P2_rEIP_PTR5 ( .D(_02189__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR5), .QN());
  DFFR_X1 P2_rEIP_PTR6 ( .D(_02189__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR6), .QN());
  DFFR_X1 P2_rEIP_PTR7 ( .D(_02189__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR7), .QN());
  DFFR_X1 P2_rEIP_PTR8 ( .D(_02189__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR8), .QN());
  DFFR_X1 P2_rEIP_PTR9 ( .D(_02189__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR9), .QN());
  DFFR_X1 P2_rEIP_PTR10 ( .D(_02189__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR10), .QN());
  DFFR_X1 P2_rEIP_PTR11 ( .D(_02189__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR11), .QN());
  DFFR_X1 P2_rEIP_PTR12 ( .D(_02189__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR12), .QN());
  DFFR_X1 P2_rEIP_PTR13 ( .D(_02189__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR13), .QN());
  DFFR_X1 P2_rEIP_PTR14 ( .D(_02189__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR14), .QN());
  DFFR_X1 P2_rEIP_PTR15 ( .D(_02189__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR15), .QN());
  DFFR_X1 P2_rEIP_PTR16 ( .D(_02189__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR16), .QN());
  DFFR_X1 P2_rEIP_PTR17 ( .D(_02189__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR17), .QN());
  DFFR_X1 P2_rEIP_PTR18 ( .D(_02189__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR18), .QN());
  DFFR_X1 P2_rEIP_PTR19 ( .D(_02189__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR19), .QN());
  DFFR_X1 P2_rEIP_PTR20 ( .D(_02189__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR20), .QN());
  DFFR_X1 P2_rEIP_PTR21 ( .D(_02189__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR21), .QN());
  DFFR_X1 P2_rEIP_PTR22 ( .D(_02189__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR22), .QN());
  DFFR_X1 P2_rEIP_PTR23 ( .D(_02189__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR23), .QN());
  DFFR_X1 P2_rEIP_PTR24 ( .D(_02189__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR24), .QN());
  DFFR_X1 P2_rEIP_PTR25 ( .D(_02189__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR25), .QN());
  DFFR_X1 P2_rEIP_PTR26 ( .D(_02189__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR26), .QN());
  DFFR_X1 P2_rEIP_PTR27 ( .D(_02189__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR27), .QN());
  DFFR_X1 P2_rEIP_PTR28 ( .D(_02189__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR28), .QN());
  DFFR_X1 P2_rEIP_PTR29 ( .D(_02189__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR29), .QN());
  DFFR_X1 P2_rEIP_PTR30 ( .D(_02189__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR30), .QN());
  DFFR_X1 P2_EBX_PTR0 ( .D(_02227__PTR160), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR0), .QN());
  DFFR_X1 P2_EBX_PTR1 ( .D(_02227__PTR161), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR1), .QN());
  DFFR_X1 P2_EBX_PTR2 ( .D(_02227__PTR162), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR2), .QN());
  DFFR_X1 P2_EBX_PTR3 ( .D(_02227__PTR163), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR3), .QN());
  DFFR_X1 P2_EBX_PTR4 ( .D(_02227__PTR164), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR4), .QN());
  DFFR_X1 P2_EBX_PTR5 ( .D(_02227__PTR165), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR5), .QN());
  DFFR_X1 P2_EBX_PTR6 ( .D(_02227__PTR166), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR6), .QN());
  DFFR_X1 P2_EBX_PTR7 ( .D(_02227__PTR167), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR7), .QN());
  DFFR_X1 P2_EBX_PTR8 ( .D(_02227__PTR168), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR8), .QN());
  DFFR_X1 P2_EBX_PTR9 ( .D(_02227__PTR169), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR9), .QN());
  DFFR_X1 P2_EBX_PTR10 ( .D(_02227__PTR170), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR10), .QN());
  DFFR_X1 P2_EBX_PTR11 ( .D(_02227__PTR171), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR11), .QN());
  DFFR_X1 P2_EBX_PTR12 ( .D(_02227__PTR172), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR12), .QN());
  DFFR_X1 P2_EBX_PTR13 ( .D(_02227__PTR173), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR13), .QN());
  DFFR_X1 P2_EBX_PTR14 ( .D(_02227__PTR174), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR14), .QN());
  DFFR_X1 P2_EBX_PTR15 ( .D(_02227__PTR175), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR15), .QN());
  DFFR_X1 P2_EBX_PTR16 ( .D(_02227__PTR176), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR16), .QN());
  DFFR_X1 P2_EBX_PTR17 ( .D(_02227__PTR177), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR17), .QN());
  DFFR_X1 P2_EBX_PTR18 ( .D(_02227__PTR178), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR18), .QN());
  DFFR_X1 P2_EBX_PTR19 ( .D(_02227__PTR179), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR19), .QN());
  DFFR_X1 P2_EBX_PTR20 ( .D(_02227__PTR180), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR20), .QN());
  DFFR_X1 P2_EBX_PTR21 ( .D(_02227__PTR181), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR21), .QN());
  DFFR_X1 P2_EBX_PTR22 ( .D(_02227__PTR182), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR22), .QN());
  DFFR_X1 P2_EBX_PTR23 ( .D(_02227__PTR183), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR23), .QN());
  DFFR_X1 P2_EBX_PTR24 ( .D(_02227__PTR184), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR24), .QN());
  DFFR_X1 P2_EBX_PTR25 ( .D(_02227__PTR185), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR25), .QN());
  DFFR_X1 P2_EBX_PTR26 ( .D(_02227__PTR186), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR26), .QN());
  DFFR_X1 P2_EBX_PTR27 ( .D(_02227__PTR187), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR27), .QN());
  DFFR_X1 P2_EBX_PTR28 ( .D(_02227__PTR188), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR28), .QN());
  DFFR_X1 P2_EBX_PTR29 ( .D(_02227__PTR189), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR29), .QN());
  DFFR_X1 P2_EBX_PTR30 ( .D(_02227__PTR190), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EBX_PTR30), .QN());
  DFFR_X1 P2_EAX_PTR0 ( .D(_02226__PTR160), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR0), .QN());
  DFFR_X1 P2_EAX_PTR1 ( .D(_02226__PTR161), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR1), .QN());
  DFFR_X1 P2_EAX_PTR2 ( .D(_02226__PTR162), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR2), .QN());
  DFFR_X1 P2_EAX_PTR3 ( .D(_02226__PTR163), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR3), .QN());
  DFFR_X1 P2_EAX_PTR4 ( .D(_02226__PTR164), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR4), .QN());
  DFFR_X1 P2_EAX_PTR5 ( .D(_02226__PTR165), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR5), .QN());
  DFFR_X1 P2_EAX_PTR6 ( .D(_02226__PTR166), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR6), .QN());
  DFFR_X1 P2_EAX_PTR7 ( .D(_02226__PTR167), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR7), .QN());
  DFFR_X1 P2_EAX_PTR8 ( .D(_02226__PTR168), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR8), .QN());
  DFFR_X1 P2_EAX_PTR9 ( .D(_02226__PTR169), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR9), .QN());
  DFFR_X1 P2_EAX_PTR10 ( .D(_02226__PTR170), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR10), .QN());
  DFFR_X1 P2_EAX_PTR11 ( .D(_02226__PTR171), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR11), .QN());
  DFFR_X1 P2_EAX_PTR12 ( .D(_02226__PTR172), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR12), .QN());
  DFFR_X1 P2_EAX_PTR13 ( .D(_02226__PTR173), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR13), .QN());
  DFFR_X1 P2_EAX_PTR14 ( .D(_02226__PTR174), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR14), .QN());
  DFFR_X1 P2_EAX_PTR15 ( .D(_02226__PTR175), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR15), .QN());
  DFFR_X1 P2_EAX_PTR16 ( .D(_02226__PTR176), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR16), .QN());
  DFFR_X1 P2_EAX_PTR17 ( .D(_02226__PTR177), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR17), .QN());
  DFFR_X1 P2_EAX_PTR18 ( .D(_02226__PTR178), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR18), .QN());
  DFFR_X1 P2_EAX_PTR19 ( .D(_02226__PTR179), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR19), .QN());
  DFFR_X1 P2_EAX_PTR20 ( .D(_02226__PTR180), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR20), .QN());
  DFFR_X1 P2_EAX_PTR21 ( .D(_02226__PTR181), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR21), .QN());
  DFFR_X1 P2_EAX_PTR22 ( .D(_02226__PTR182), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR22), .QN());
  DFFR_X1 P2_EAX_PTR23 ( .D(_02226__PTR183), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR23), .QN());
  DFFR_X1 P2_EAX_PTR24 ( .D(_02226__PTR184), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR24), .QN());
  DFFR_X1 P2_EAX_PTR25 ( .D(_02226__PTR185), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR25), .QN());
  DFFR_X1 P2_EAX_PTR26 ( .D(_02226__PTR186), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR26), .QN());
  DFFR_X1 P2_EAX_PTR27 ( .D(_02226__PTR187), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR27), .QN());
  DFFR_X1 P2_EAX_PTR28 ( .D(_02226__PTR188), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR28), .QN());
  DFFR_X1 P2_EAX_PTR29 ( .D(_02226__PTR189), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR29), .QN());
  DFFR_X1 P2_EAX_PTR30 ( .D(_02226__PTR190), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_EAX_PTR30), .QN());
  DFFR_X1 P2_Datao_PTR0 ( .D(_03164__PTR256), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR0), .QN());
  DFFR_X1 P2_Datao_PTR1 ( .D(_03164__PTR257), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR1), .QN());
  DFFR_X1 P2_Datao_PTR2 ( .D(_03164__PTR258), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR2), .QN());
  DFFR_X1 P2_Datao_PTR3 ( .D(_03164__PTR259), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR3), .QN());
  DFFR_X1 P2_Datao_PTR4 ( .D(_03164__PTR260), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR4), .QN());
  DFFR_X1 P2_Datao_PTR5 ( .D(_03164__PTR261), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR5), .QN());
  DFFR_X1 P2_Datao_PTR6 ( .D(_03164__PTR262), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR6), .QN());
  DFFR_X1 P2_Datao_PTR7 ( .D(_03164__PTR263), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR7), .QN());
  DFFR_X1 P2_Datao_PTR8 ( .D(_03164__PTR264), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR8), .QN());
  DFFR_X1 P2_Datao_PTR9 ( .D(_03164__PTR265), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR9), .QN());
  DFFR_X1 P2_Datao_PTR10 ( .D(_03164__PTR266), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR10), .QN());
  DFFR_X1 P2_Datao_PTR11 ( .D(_03164__PTR267), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR11), .QN());
  DFFR_X1 P2_Datao_PTR12 ( .D(_03164__PTR268), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR12), .QN());
  DFFR_X1 P2_Datao_PTR13 ( .D(_03164__PTR269), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR13), .QN());
  DFFR_X1 P2_Datao_PTR14 ( .D(_03164__PTR270), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR14), .QN());
  DFFR_X1 P2_Datao_PTR15 ( .D(_03164__PTR271), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR15), .QN());
  DFFR_X1 P2_Datao_PTR16 ( .D(_03164__PTR272), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR16), .QN());
  DFFR_X1 P2_Datao_PTR17 ( .D(_03164__PTR273), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR17), .QN());
  DFFR_X1 P2_Datao_PTR18 ( .D(_03164__PTR274), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR18), .QN());
  DFFR_X1 P2_Datao_PTR19 ( .D(_03164__PTR275), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR19), .QN());
  DFFR_X1 P2_Datao_PTR20 ( .D(_03164__PTR276), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR20), .QN());
  DFFR_X1 P2_Datao_PTR21 ( .D(_03164__PTR277), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR21), .QN());
  DFFR_X1 P2_Datao_PTR22 ( .D(_03164__PTR278), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR22), .QN());
  DFFR_X1 P2_Datao_PTR23 ( .D(_03164__PTR279), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR23), .QN());
  DFFR_X1 P2_Datao_PTR24 ( .D(_03164__PTR280), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR24), .QN());
  DFFR_X1 P2_Datao_PTR25 ( .D(_03164__PTR281), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR25), .QN());
  DFFR_X1 P2_Datao_PTR26 ( .D(_03164__PTR282), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR26), .QN());
  DFFR_X1 P2_Datao_PTR27 ( .D(_03164__PTR283), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR27), .QN());
  DFFR_X1 P2_Datao_PTR28 ( .D(_03164__PTR284), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR28), .QN());
  DFFR_X1 P2_Datao_PTR29 ( .D(_03164__PTR285), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR29), .QN());
  DFFR_X1 P2_Datao_PTR30 ( .D(_03164__PTR286), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR30), .QN());
  DFFR_X1 P2_DataWidth_reg_PTR0 ( .D(_02171__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR0), .QN());
  BUF_X1 U37 ( .A(P2_DataWidth_reg_PTR0), .Z(P2_DataWidth_PTR0) );
  DFFR_X1 P2_DataWidth_reg_PTR2 ( .D(_02171__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR2), .QN());
  BUF_X1 U38 ( .A(P2_DataWidth_reg_PTR2), .Z(P2_DataWidth_PTR2) );
  DFFR_X1 P2_DataWidth_reg_PTR3 ( .D(_02171__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR3), .QN());
  BUF_X1 U39 ( .A(P2_DataWidth_reg_PTR3), .Z(P2_DataWidth_PTR3) );
  DFFR_X1 P2_DataWidth_reg_PTR4 ( .D(_02171__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR4), .QN());
  BUF_X1 U40 ( .A(P2_DataWidth_reg_PTR4), .Z(P2_DataWidth_PTR4) );
  DFFR_X1 P2_DataWidth_reg_PTR5 ( .D(_02171__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR5), .QN());
  BUF_X1 U41 ( .A(P2_DataWidth_reg_PTR5), .Z(P2_DataWidth_PTR5) );
  DFFR_X1 P2_DataWidth_reg_PTR6 ( .D(_02171__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR6), .QN());
  BUF_X1 U42 ( .A(P2_DataWidth_reg_PTR6), .Z(P2_DataWidth_PTR6) );
  DFFR_X1 P2_DataWidth_reg_PTR7 ( .D(_02171__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR7), .QN());
  BUF_X1 U43 ( .A(P2_DataWidth_reg_PTR7), .Z(P2_DataWidth_PTR7) );
  DFFR_X1 P2_DataWidth_reg_PTR8 ( .D(_02171__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR8), .QN());
  BUF_X1 U44 ( .A(P2_DataWidth_reg_PTR8), .Z(P2_DataWidth_PTR8) );
  DFFR_X1 P2_DataWidth_reg_PTR9 ( .D(_02171__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR9), .QN());
  BUF_X1 U45 ( .A(P2_DataWidth_reg_PTR9), .Z(P2_DataWidth_PTR9) );
  DFFR_X1 P2_DataWidth_reg_PTR10 ( .D(_02171__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR10), .QN());
  BUF_X1 U46 ( .A(P2_DataWidth_reg_PTR10), .Z(P2_DataWidth_PTR10) );
  DFFR_X1 P2_DataWidth_reg_PTR11 ( .D(_02171__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR11), .QN());
  BUF_X1 U47 ( .A(P2_DataWidth_reg_PTR11), .Z(P2_DataWidth_PTR11) );
  DFFR_X1 P2_DataWidth_reg_PTR12 ( .D(_02171__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR12), .QN());
  BUF_X1 U48 ( .A(P2_DataWidth_reg_PTR12), .Z(P2_DataWidth_PTR12) );
  DFFR_X1 P2_DataWidth_reg_PTR13 ( .D(_02171__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR13), .QN());
  BUF_X1 U49 ( .A(P2_DataWidth_reg_PTR13), .Z(P2_DataWidth_PTR13) );
  DFFR_X1 P2_DataWidth_reg_PTR14 ( .D(_02171__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR14), .QN());
  BUF_X1 U50 ( .A(P2_DataWidth_reg_PTR14), .Z(P2_DataWidth_PTR14) );
  DFFR_X1 P2_DataWidth_reg_PTR15 ( .D(_02171__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR15), .QN());
  BUF_X1 U51 ( .A(P2_DataWidth_reg_PTR15), .Z(P2_DataWidth_PTR15) );
  DFFR_X1 P2_DataWidth_reg_PTR16 ( .D(_02171__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR16), .QN());
  BUF_X1 U52 ( .A(P2_DataWidth_reg_PTR16), .Z(P2_DataWidth_PTR16) );
  DFFR_X1 P2_DataWidth_reg_PTR17 ( .D(_02171__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR17), .QN());
  BUF_X1 U53 ( .A(P2_DataWidth_reg_PTR17), .Z(P2_DataWidth_PTR17) );
  DFFR_X1 P2_DataWidth_reg_PTR18 ( .D(_02171__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR18), .QN());
  BUF_X1 U54 ( .A(P2_DataWidth_reg_PTR18), .Z(P2_DataWidth_PTR18) );
  DFFR_X1 P2_DataWidth_reg_PTR19 ( .D(_02171__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR19), .QN());
  BUF_X1 U55 ( .A(P2_DataWidth_reg_PTR19), .Z(P2_DataWidth_PTR19) );
  DFFR_X1 P2_DataWidth_reg_PTR20 ( .D(_02171__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR20), .QN());
  BUF_X1 U56 ( .A(P2_DataWidth_reg_PTR20), .Z(P2_DataWidth_PTR20) );
  DFFR_X1 P2_DataWidth_reg_PTR21 ( .D(_02171__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR21), .QN());
  BUF_X1 U57 ( .A(P2_DataWidth_reg_PTR21), .Z(P2_DataWidth_PTR21) );
  DFFR_X1 P2_DataWidth_reg_PTR22 ( .D(_02171__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR22), .QN());
  BUF_X1 U58 ( .A(P2_DataWidth_reg_PTR22), .Z(P2_DataWidth_PTR22) );
  DFFR_X1 P2_DataWidth_reg_PTR23 ( .D(_02171__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR23), .QN());
  BUF_X1 U59 ( .A(P2_DataWidth_reg_PTR23), .Z(P2_DataWidth_PTR23) );
  DFFR_X1 P2_DataWidth_reg_PTR24 ( .D(_02171__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR24), .QN());
  BUF_X1 U60 ( .A(P2_DataWidth_reg_PTR24), .Z(P2_DataWidth_PTR24) );
  DFFR_X1 P2_DataWidth_reg_PTR25 ( .D(_02171__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR25), .QN());
  BUF_X1 U61 ( .A(P2_DataWidth_reg_PTR25), .Z(P2_DataWidth_PTR25) );
  DFFR_X1 P2_DataWidth_reg_PTR26 ( .D(_02171__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR26), .QN());
  BUF_X1 U62 ( .A(P2_DataWidth_reg_PTR26), .Z(P2_DataWidth_PTR26) );
  DFFR_X1 P2_DataWidth_reg_PTR27 ( .D(_02171__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR27), .QN());
  BUF_X1 U63 ( .A(P2_DataWidth_reg_PTR27), .Z(P2_DataWidth_PTR27) );
  DFFR_X1 P2_DataWidth_reg_PTR28 ( .D(_02171__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR28), .QN());
  BUF_X1 U64 ( .A(P2_DataWidth_reg_PTR28), .Z(P2_DataWidth_PTR28) );
  DFFR_X1 P2_DataWidth_reg_PTR29 ( .D(_02171__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR29), .QN());
  BUF_X1 U65 ( .A(P2_DataWidth_reg_PTR29), .Z(P2_DataWidth_PTR29) );
  DFFR_X1 P2_DataWidth_reg_PTR30 ( .D(_02171__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR30), .QN());
  BUF_X1 U66 ( .A(P2_DataWidth_reg_PTR30), .Z(P2_DataWidth_PTR30) );
  DFFR_X1 P2_State_PTR0 ( .D(_02170__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_State_PTR0), .QN());
  DFFR_X1 P2_State_PTR1 ( .D(_02170__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_State_PTR1), .QN());
  DFFR_X1 P2_Address_PTR0 ( .D(_02173__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR0), .QN());
  DFFR_X1 P2_Address_PTR1 ( .D(_02173__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR1), .QN());
  DFFR_X1 P2_Address_PTR2 ( .D(_02173__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR2), .QN());
  DFFR_X1 P2_Address_PTR3 ( .D(_02173__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR3), .QN());
  DFFR_X1 P2_Address_PTR4 ( .D(_02173__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR4), .QN());
  DFFR_X1 P2_Address_PTR5 ( .D(_02173__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR5), .QN());
  DFFR_X1 P2_Address_PTR6 ( .D(_02173__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR6), .QN());
  DFFR_X1 P2_Address_PTR7 ( .D(_02173__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR7), .QN());
  DFFR_X1 P2_Address_PTR8 ( .D(_02173__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR8), .QN());
  DFFR_X1 P2_Address_PTR9 ( .D(_02173__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR9), .QN());
  DFFR_X1 P2_Address_PTR10 ( .D(_02173__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR10), .QN());
  DFFR_X1 P2_Address_PTR11 ( .D(_02173__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR11), .QN());
  DFFR_X1 P2_Address_PTR12 ( .D(_02173__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR12), .QN());
  DFFR_X1 P2_Address_PTR13 ( .D(_02173__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR13), .QN());
  DFFR_X1 P2_Address_PTR14 ( .D(_02173__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR14), .QN());
  DFFR_X1 P2_Address_PTR15 ( .D(_02173__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR15), .QN());
  DFFR_X1 P2_Address_PTR16 ( .D(_02173__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR16), .QN());
  DFFR_X1 P2_Address_PTR17 ( .D(_02173__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR17), .QN());
  DFFR_X1 P2_Address_PTR18 ( .D(_02173__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR18), .QN());
  DFFR_X1 P2_Address_PTR19 ( .D(_02173__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR19), .QN());
  DFFR_X1 P2_Address_PTR20 ( .D(_02173__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR20), .QN());
  DFFR_X1 P2_Address_PTR21 ( .D(_02173__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR21), .QN());
  DFFR_X1 P2_Address_PTR22 ( .D(_02173__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR22), .QN());
  DFFR_X1 P2_Address_PTR23 ( .D(_02173__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR23), .QN());
  DFFR_X1 P2_Address_PTR24 ( .D(_02173__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR24), .QN());
  DFFR_X1 P2_Address_PTR25 ( .D(_02173__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR25), .QN());
  DFFR_X1 P2_Address_PTR26 ( .D(_02173__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR26), .QN());
  DFFR_X1 P2_Address_PTR27 ( .D(_02173__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR27), .QN());
  DFFR_X1 P2_Address_PTR28 ( .D(_02173__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Address_PTR28), .QN());
  DFFR_X1 P2_P1_uWord_PTR0 ( .D(_02228__PTR80), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR0), .QN());
  DFFR_X1 P2_P1_uWord_PTR1 ( .D(_02228__PTR81), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR1), .QN());
  DFFR_X1 P2_P1_uWord_PTR2 ( .D(_02228__PTR82), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR2), .QN());
  DFFR_X1 P2_P1_uWord_PTR3 ( .D(_02228__PTR83), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR3), .QN());
  DFFR_X1 P2_P1_uWord_PTR4 ( .D(_02228__PTR84), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR4), .QN());
  DFFR_X1 P2_P1_uWord_PTR5 ( .D(_02228__PTR85), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR5), .QN());
  DFFR_X1 P2_P1_uWord_PTR6 ( .D(_02228__PTR86), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR6), .QN());
  DFFR_X1 P2_P1_uWord_PTR7 ( .D(_02228__PTR87), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR7), .QN());
  DFFR_X1 P2_P1_uWord_PTR8 ( .D(_02228__PTR88), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR8), .QN());
  DFFR_X1 P2_P1_uWord_PTR9 ( .D(_02228__PTR89), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR9), .QN());
  DFFR_X1 P2_P1_uWord_PTR10 ( .D(_02228__PTR90), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR10), .QN());
  DFFR_X1 P2_P1_uWord_PTR11 ( .D(_02228__PTR91), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR11), .QN());
  DFFR_X1 P2_P1_uWord_PTR12 ( .D(_02228__PTR92), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR12), .QN());
  DFFR_X1 P2_P1_uWord_PTR13 ( .D(_02228__PTR93), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_uWord_PTR13), .QN());
  DFFR_X1 P2_P1_lWord_PTR0 ( .D(_02229__PTR80), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR0), .QN());
  DFFR_X1 P2_P1_lWord_PTR1 ( .D(_02229__PTR81), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR1), .QN());
  DFFR_X1 P2_P1_lWord_PTR2 ( .D(_02229__PTR82), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR2), .QN());
  DFFR_X1 P2_P1_lWord_PTR3 ( .D(_02229__PTR83), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR3), .QN());
  DFFR_X1 P2_P1_lWord_PTR4 ( .D(_02229__PTR84), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR4), .QN());
  DFFR_X1 P2_P1_lWord_PTR5 ( .D(_02229__PTR85), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR5), .QN());
  DFFR_X1 P2_P1_lWord_PTR6 ( .D(_02229__PTR86), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR6), .QN());
  DFFR_X1 P2_P1_lWord_PTR7 ( .D(_02229__PTR87), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR7), .QN());
  DFFR_X1 P2_P1_lWord_PTR8 ( .D(_02229__PTR88), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR8), .QN());
  DFFR_X1 P2_P1_lWord_PTR9 ( .D(_02229__PTR89), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR9), .QN());
  DFFR_X1 P2_P1_lWord_PTR10 ( .D(_02229__PTR90), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR10), .QN());
  DFFR_X1 P2_P1_lWord_PTR11 ( .D(_02229__PTR91), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR11), .QN());
  DFFR_X1 P2_P1_lWord_PTR12 ( .D(_02229__PTR92), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR12), .QN());
  DFFR_X1 P2_P1_lWord_PTR13 ( .D(_02229__PTR93), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR13), .QN());
  DFFR_X1 P2_P1_lWord_PTR14 ( .D(_02229__PTR94), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_lWord_PTR14), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR0 ( .D(_03098__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR0), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR1 ( .D(_03098__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR1), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR2 ( .D(_03098__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR2), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR3 ( .D(_03098__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR3), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR4 ( .D(_03098__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR4), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR5 ( .D(_03098__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR5), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR6 ( .D(_03098__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR6), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR7 ( .D(_03098__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR7), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR8 ( .D(_03098__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR8), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR9 ( .D(_03098__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR9), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR10 ( .D(_03098__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR10), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR11 ( .D(_03098__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR11), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR12 ( .D(_03098__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR12), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR13 ( .D(_03098__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR13), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR14 ( .D(_03098__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR14), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR15 ( .D(_03098__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR15), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR16 ( .D(_03098__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR16), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR17 ( .D(_03098__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR17), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR18 ( .D(_03098__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR18), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR19 ( .D(_03098__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR19), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR20 ( .D(_03098__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR20), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR21 ( .D(_03098__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR21), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR22 ( .D(_03098__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR22), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR23 ( .D(_03098__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR23), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR24 ( .D(_03098__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR24), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR25 ( .D(_03098__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR25), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR26 ( .D(_03098__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR26), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR27 ( .D(_03098__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR27), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR28 ( .D(_03098__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR28), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR29 ( .D(_03098__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR29), .QN());
  DFFR_X1 P2_P1_PhyAddrPointer_PTR30 ( .D(_03098__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_PhyAddrPointer_PTR30), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR0 ( .D(_03101__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR0), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR1 ( .D(_03101__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR1), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR2 ( .D(_03101__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR2), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR3 ( .D(_03101__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR3), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR4 ( .D(_03101__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR4), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR5 ( .D(_03101__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR5), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR6 ( .D(_03101__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR6), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR7 ( .D(_03101__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR7), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR8 ( .D(_03101__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR8), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR9 ( .D(_03101__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR9), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR10 ( .D(_03101__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR10), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR11 ( .D(_03101__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR11), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR12 ( .D(_03101__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR12), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR13 ( .D(_03101__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR13), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR14 ( .D(_03101__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR14), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR15 ( .D(_03101__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR15), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR16 ( .D(_03101__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR16), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR17 ( .D(_03101__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR17), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR18 ( .D(_03101__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR18), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR19 ( .D(_03101__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR19), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR20 ( .D(_03101__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR20), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR21 ( .D(_03101__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR21), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR22 ( .D(_03101__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR22), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR23 ( .D(_03101__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR23), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR24 ( .D(_03101__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR24), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR25 ( .D(_03101__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR25), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR26 ( .D(_03101__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR26), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR27 ( .D(_03101__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR27), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR28 ( .D(_03101__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR28), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR29 ( .D(_03101__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR29), .QN());
  DFFR_X1 P2_P1_InstAddrPointer_PTR30 ( .D(_03101__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstAddrPointer_PTR30), .QN());
  DFFR_X1 P2_P1_InstQueueWr_Addr_PTR0 ( .D(_02223__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueueWr_Addr_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueueWr_Addr_PTR1 ( .D(_02223__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueueWr_Addr_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueueWr_Addr_PTR2 ( .D(_02223__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueueWr_Addr_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueueWr_Addr_PTR3 ( .D(_02223__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueueWr_Addr_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueueRd_Addr_PTR0 ( .D(_02225__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueueRd_Addr_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueueRd_Addr_PTR1 ( .D(_02225__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueueRd_Addr_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueueRd_Addr_PTR2 ( .D(_02225__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueueRd_Addr_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueueRd_Addr_PTR3 ( .D(_02225__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueueRd_Addr_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR0_PTR0 ( .D(_02221__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR0_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR0_PTR1 ( .D(_02221__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR0_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR0_PTR2 ( .D(_02221__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR0_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR0_PTR3 ( .D(_02221__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR0_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR0_PTR4 ( .D(_02221__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR0_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR0_PTR5 ( .D(_02221__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR0_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR0_PTR6 ( .D(_02221__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR0_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR1_PTR0 ( .D(_02219__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR1_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR1_PTR1 ( .D(_02219__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR1_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR1_PTR2 ( .D(_02219__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR1_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR1_PTR3 ( .D(_02219__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR1_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR1_PTR4 ( .D(_02219__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR1_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR1_PTR5 ( .D(_02219__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR1_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR1_PTR6 ( .D(_02219__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR1_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR2_PTR0 ( .D(_02217__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR2_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR2_PTR1 ( .D(_02217__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR2_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR2_PTR2 ( .D(_02217__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR2_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR2_PTR3 ( .D(_02217__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR2_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR2_PTR4 ( .D(_02217__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR2_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR2_PTR5 ( .D(_02217__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR2_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR2_PTR6 ( .D(_02217__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR2_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR3_PTR0 ( .D(_02215__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR3_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR3_PTR1 ( .D(_02215__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR3_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR3_PTR2 ( .D(_02215__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR3_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR3_PTR3 ( .D(_02215__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR3_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR3_PTR4 ( .D(_02215__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR3_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR3_PTR5 ( .D(_02215__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR3_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR3_PTR6 ( .D(_02215__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR3_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR4_PTR0 ( .D(_02213__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR4_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR4_PTR1 ( .D(_02213__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR4_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR4_PTR2 ( .D(_02213__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR4_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR4_PTR3 ( .D(_02213__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR4_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR4_PTR4 ( .D(_02213__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR4_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR4_PTR5 ( .D(_02213__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR4_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR4_PTR6 ( .D(_02213__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR4_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR5_PTR0 ( .D(_02211__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR5_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR5_PTR1 ( .D(_02211__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR5_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR5_PTR2 ( .D(_02211__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR5_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR5_PTR3 ( .D(_02211__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR5_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR5_PTR4 ( .D(_02211__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR5_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR5_PTR5 ( .D(_02211__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR5_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR5_PTR6 ( .D(_02211__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR5_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR6_PTR0 ( .D(_02209__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR6_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR6_PTR1 ( .D(_02209__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR6_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR6_PTR2 ( .D(_02209__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR6_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR6_PTR3 ( .D(_02209__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR6_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR6_PTR4 ( .D(_02209__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR6_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR6_PTR5 ( .D(_02209__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR6_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR6_PTR6 ( .D(_02209__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR6_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR7_PTR0 ( .D(_02207__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR7_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR7_PTR1 ( .D(_02207__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR7_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR7_PTR2 ( .D(_02207__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR7_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR7_PTR3 ( .D(_02207__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR7_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR7_PTR4 ( .D(_02207__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR7_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR7_PTR5 ( .D(_02207__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR7_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR7_PTR6 ( .D(_02207__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR7_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR8_PTR0 ( .D(_02205__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR8_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR8_PTR1 ( .D(_02205__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR8_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR8_PTR2 ( .D(_02205__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR8_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR8_PTR3 ( .D(_02205__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR8_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR8_PTR4 ( .D(_02205__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR8_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR8_PTR5 ( .D(_02205__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR8_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR8_PTR6 ( .D(_02205__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR8_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR9_PTR0 ( .D(_02203__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR9_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR9_PTR1 ( .D(_02203__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR9_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR9_PTR2 ( .D(_02203__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR9_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR9_PTR3 ( .D(_02203__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR9_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR9_PTR4 ( .D(_02203__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR9_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR9_PTR5 ( .D(_02203__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR9_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR9_PTR6 ( .D(_02203__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR9_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR10_PTR0 ( .D(_02201__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR10_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR10_PTR1 ( .D(_02201__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR10_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR10_PTR2 ( .D(_02201__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR10_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR10_PTR3 ( .D(_02201__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR10_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR10_PTR4 ( .D(_02201__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR10_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR10_PTR5 ( .D(_02201__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR10_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR10_PTR6 ( .D(_02201__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR10_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR11_PTR0 ( .D(_02199__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR11_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR11_PTR1 ( .D(_02199__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR11_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR11_PTR2 ( .D(_02199__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR11_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR11_PTR3 ( .D(_02199__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR11_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR11_PTR4 ( .D(_02199__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR11_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR11_PTR5 ( .D(_02199__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR11_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR11_PTR6 ( .D(_02199__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR11_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR12_PTR0 ( .D(_02197__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR12_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR12_PTR1 ( .D(_02197__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR12_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR12_PTR2 ( .D(_02197__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR12_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR12_PTR3 ( .D(_02197__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR12_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR12_PTR4 ( .D(_02197__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR12_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR12_PTR5 ( .D(_02197__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR12_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR12_PTR6 ( .D(_02197__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR12_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR13_PTR0 ( .D(_02195__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR13_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR13_PTR1 ( .D(_02195__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR13_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR13_PTR2 ( .D(_02195__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR13_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR13_PTR3 ( .D(_02195__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR13_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR13_PTR4 ( .D(_02195__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR13_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR13_PTR5 ( .D(_02195__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR13_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR13_PTR6 ( .D(_02195__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR13_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR14_PTR0 ( .D(_02193__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR14_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR14_PTR1 ( .D(_02193__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR14_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR14_PTR2 ( .D(_02193__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR14_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR14_PTR3 ( .D(_02193__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR14_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR14_PTR4 ( .D(_02193__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR14_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR14_PTR5 ( .D(_02193__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR14_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR14_PTR6 ( .D(_02193__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR14_PTR6), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR15_PTR0 ( .D(_02191__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR15_PTR0), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR15_PTR1 ( .D(_02191__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR15_PTR1), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR15_PTR2 ( .D(_02191__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR15_PTR2), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR15_PTR3 ( .D(_02191__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR15_PTR3), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR15_PTR4 ( .D(_02191__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR15_PTR4), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR15_PTR5 ( .D(_02191__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR15_PTR5), .QN());
  DFFR_X1 P2_P1_InstQueue_PTR15_PTR6 ( .D(_02191__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_InstQueue_PTR15_PTR6), .QN());
  DFFR_X1 P2_P1_State2_PTR0 ( .D(_02187__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_State2_PTR0), .QN());
  DFFR_X1 P2_P1_State2_PTR1 ( .D(_02187__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_State2_PTR1), .QN());
  DFFR_X1 P2_P1_State2_PTR2 ( .D(_02187__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_P1_State2_PTR2), .QN());
  DFFR_X1 P3_rEIP_PTR0 ( .D(_02478__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR0), .QN());
  DFFR_X1 P3_rEIP_PTR1 ( .D(_02478__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR1), .QN());
  DFFR_X1 P3_rEIP_PTR2 ( .D(_02478__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR2), .QN());
  DFFR_X1 P3_rEIP_PTR3 ( .D(_02478__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR3), .QN());
  DFFR_X1 P3_rEIP_PTR4 ( .D(_02478__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR4), .QN());
  DFFR_X1 P3_rEIP_PTR5 ( .D(_02478__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR5), .QN());
  DFFR_X1 P3_rEIP_PTR6 ( .D(_02478__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR6), .QN());
  DFFR_X1 P3_rEIP_PTR7 ( .D(_02478__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR7), .QN());
  DFFR_X1 P3_rEIP_PTR8 ( .D(_02478__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR8), .QN());
  DFFR_X1 P3_rEIP_PTR9 ( .D(_02478__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR9), .QN());
  DFFR_X1 P3_rEIP_PTR10 ( .D(_02478__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR10), .QN());
  DFFR_X1 P3_rEIP_PTR11 ( .D(_02478__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR11), .QN());
  DFFR_X1 P3_rEIP_PTR12 ( .D(_02478__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR12), .QN());
  DFFR_X1 P3_rEIP_PTR13 ( .D(_02478__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR13), .QN());
  DFFR_X1 P3_rEIP_PTR14 ( .D(_02478__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR14), .QN());
  DFFR_X1 P3_rEIP_PTR15 ( .D(_02478__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR15), .QN());
  DFFR_X1 P3_rEIP_PTR16 ( .D(_02478__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR16), .QN());
  DFFR_X1 P3_rEIP_PTR17 ( .D(_02478__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR17), .QN());
  DFFR_X1 P3_rEIP_PTR18 ( .D(_02478__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR18), .QN());
  DFFR_X1 P3_rEIP_PTR19 ( .D(_02478__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR19), .QN());
  DFFR_X1 P3_rEIP_PTR20 ( .D(_02478__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR20), .QN());
  DFFR_X1 P3_rEIP_PTR21 ( .D(_02478__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR21), .QN());
  DFFR_X1 P3_rEIP_PTR22 ( .D(_02478__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR22), .QN());
  DFFR_X1 P3_rEIP_PTR23 ( .D(_02478__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR23), .QN());
  DFFR_X1 P3_rEIP_PTR24 ( .D(_02478__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR24), .QN());
  DFFR_X1 P3_rEIP_PTR25 ( .D(_02478__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR25), .QN());
  DFFR_X1 P3_rEIP_PTR26 ( .D(_02478__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR26), .QN());
  DFFR_X1 P3_rEIP_PTR27 ( .D(_02478__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR27), .QN());
  DFFR_X1 P3_rEIP_PTR28 ( .D(_02478__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR28), .QN());
  DFFR_X1 P3_rEIP_PTR29 ( .D(_02478__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR29), .QN());
  DFFR_X1 P3_rEIP_PTR30 ( .D(_02478__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR30), .QN());
  DFFR_X1 P3_EBX_PTR0 ( .D(_02516__PTR160), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR0), .QN());
  DFFR_X1 P3_EBX_PTR1 ( .D(_02516__PTR161), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR1), .QN());
  DFFR_X1 P3_EBX_PTR2 ( .D(_02516__PTR162), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR2), .QN());
  DFFR_X1 P3_EBX_PTR3 ( .D(_02516__PTR163), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR3), .QN());
  DFFR_X1 P3_EBX_PTR4 ( .D(_02516__PTR164), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR4), .QN());
  DFFR_X1 P3_EBX_PTR5 ( .D(_02516__PTR165), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR5), .QN());
  DFFR_X1 P3_EBX_PTR6 ( .D(_02516__PTR166), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR6), .QN());
  DFFR_X1 P3_EBX_PTR7 ( .D(_02516__PTR167), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR7), .QN());
  DFFR_X1 P3_EBX_PTR8 ( .D(_02516__PTR168), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR8), .QN());
  DFFR_X1 P3_EBX_PTR9 ( .D(_02516__PTR169), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR9), .QN());
  DFFR_X1 P3_EBX_PTR10 ( .D(_02516__PTR170), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR10), .QN());
  DFFR_X1 P3_EBX_PTR11 ( .D(_02516__PTR171), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR11), .QN());
  DFFR_X1 P3_EBX_PTR12 ( .D(_02516__PTR172), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR12), .QN());
  DFFR_X1 P3_EBX_PTR13 ( .D(_02516__PTR173), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR13), .QN());
  DFFR_X1 P3_EBX_PTR14 ( .D(_02516__PTR174), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR14), .QN());
  DFFR_X1 P3_EBX_PTR15 ( .D(_02516__PTR175), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR15), .QN());
  DFFR_X1 P3_EBX_PTR16 ( .D(_02516__PTR176), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR16), .QN());
  DFFR_X1 P3_EBX_PTR17 ( .D(_02516__PTR177), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR17), .QN());
  DFFR_X1 P3_EBX_PTR18 ( .D(_02516__PTR178), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR18), .QN());
  DFFR_X1 P3_EBX_PTR19 ( .D(_02516__PTR179), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR19), .QN());
  DFFR_X1 P3_EBX_PTR20 ( .D(_02516__PTR180), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR20), .QN());
  DFFR_X1 P3_EBX_PTR21 ( .D(_02516__PTR181), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR21), .QN());
  DFFR_X1 P3_EBX_PTR22 ( .D(_02516__PTR182), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR22), .QN());
  DFFR_X1 P3_EBX_PTR23 ( .D(_02516__PTR183), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR23), .QN());
  DFFR_X1 P3_EBX_PTR24 ( .D(_02516__PTR184), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR24), .QN());
  DFFR_X1 P3_EBX_PTR25 ( .D(_02516__PTR185), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR25), .QN());
  DFFR_X1 P3_EBX_PTR26 ( .D(_02516__PTR186), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR26), .QN());
  DFFR_X1 P3_EBX_PTR27 ( .D(_02516__PTR187), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR27), .QN());
  DFFR_X1 P3_EBX_PTR28 ( .D(_02516__PTR188), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR28), .QN());
  DFFR_X1 P3_EBX_PTR29 ( .D(_02516__PTR189), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR29), .QN());
  DFFR_X1 P3_EBX_PTR30 ( .D(_02516__PTR190), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EBX_PTR30), .QN());
  DFFR_X1 P3_EAX_PTR0 ( .D(_02515__PTR160), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR0), .QN());
  DFFR_X1 P3_EAX_PTR1 ( .D(_02515__PTR161), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR1), .QN());
  DFFR_X1 P3_EAX_PTR2 ( .D(_02515__PTR162), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR2), .QN());
  DFFR_X1 P3_EAX_PTR3 ( .D(_02515__PTR163), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR3), .QN());
  DFFR_X1 P3_EAX_PTR4 ( .D(_02515__PTR164), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR4), .QN());
  DFFR_X1 P3_EAX_PTR5 ( .D(_02515__PTR165), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR5), .QN());
  DFFR_X1 P3_EAX_PTR6 ( .D(_02515__PTR166), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR6), .QN());
  DFFR_X1 P3_EAX_PTR7 ( .D(_02515__PTR167), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR7), .QN());
  DFFR_X1 P3_EAX_PTR8 ( .D(_02515__PTR168), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR8), .QN());
  DFFR_X1 P3_EAX_PTR9 ( .D(_02515__PTR169), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR9), .QN());
  DFFR_X1 P3_EAX_PTR10 ( .D(_02515__PTR170), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR10), .QN());
  DFFR_X1 P3_EAX_PTR11 ( .D(_02515__PTR171), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR11), .QN());
  DFFR_X1 P3_EAX_PTR12 ( .D(_02515__PTR172), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR12), .QN());
  DFFR_X1 P3_EAX_PTR13 ( .D(_02515__PTR173), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR13), .QN());
  DFFR_X1 P3_EAX_PTR14 ( .D(_02515__PTR174), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR14), .QN());
  DFFR_X1 P3_EAX_PTR15 ( .D(_02515__PTR175), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR15), .QN());
  DFFR_X1 P3_EAX_PTR16 ( .D(_02515__PTR176), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR16), .QN());
  DFFR_X1 P3_EAX_PTR17 ( .D(_02515__PTR177), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR17), .QN());
  DFFR_X1 P3_EAX_PTR18 ( .D(_02515__PTR178), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR18), .QN());
  DFFR_X1 P3_EAX_PTR19 ( .D(_02515__PTR179), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR19), .QN());
  DFFR_X1 P3_EAX_PTR20 ( .D(_02515__PTR180), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR20), .QN());
  DFFR_X1 P3_EAX_PTR21 ( .D(_02515__PTR181), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR21), .QN());
  DFFR_X1 P3_EAX_PTR22 ( .D(_02515__PTR182), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR22), .QN());
  DFFR_X1 P3_EAX_PTR23 ( .D(_02515__PTR183), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR23), .QN());
  DFFR_X1 P3_EAX_PTR24 ( .D(_02515__PTR184), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR24), .QN());
  DFFR_X1 P3_EAX_PTR25 ( .D(_02515__PTR185), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR25), .QN());
  DFFR_X1 P3_EAX_PTR26 ( .D(_02515__PTR186), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR26), .QN());
  DFFR_X1 P3_EAX_PTR27 ( .D(_02515__PTR187), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR27), .QN());
  DFFR_X1 P3_EAX_PTR28 ( .D(_02515__PTR188), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR28), .QN());
  DFFR_X1 P3_EAX_PTR29 ( .D(_02515__PTR189), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR29), .QN());
  DFFR_X1 P3_EAX_PTR30 ( .D(_02515__PTR190), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_EAX_PTR30), .QN());
  DFFR_X1 P3_Datao_PTR0 ( .D(_03409__PTR256), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR0), .QN());
  DFFR_X1 P3_Datao_PTR1 ( .D(_03409__PTR257), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR1), .QN());
  DFFR_X1 P3_Datao_PTR2 ( .D(_03409__PTR258), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR2), .QN());
  DFFR_X1 P3_Datao_PTR3 ( .D(_03409__PTR259), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR3), .QN());
  DFFR_X1 P3_Datao_PTR4 ( .D(_03409__PTR260), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR4), .QN());
  DFFR_X1 P3_Datao_PTR5 ( .D(_03409__PTR261), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR5), .QN());
  DFFR_X1 P3_Datao_PTR6 ( .D(_03409__PTR262), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR6), .QN());
  DFFR_X1 P3_Datao_PTR7 ( .D(_03409__PTR263), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR7), .QN());
  DFFR_X1 P3_Datao_PTR8 ( .D(_03409__PTR264), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR8), .QN());
  DFFR_X1 P3_Datao_PTR9 ( .D(_03409__PTR265), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR9), .QN());
  DFFR_X1 P3_Datao_PTR10 ( .D(_03409__PTR266), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR10), .QN());
  DFFR_X1 P3_Datao_PTR11 ( .D(_03409__PTR267), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR11), .QN());
  DFFR_X1 P3_Datao_PTR12 ( .D(_03409__PTR268), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR12), .QN());
  DFFR_X1 P3_Datao_PTR13 ( .D(_03409__PTR269), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR13), .QN());
  DFFR_X1 P3_Datao_PTR14 ( .D(_03409__PTR270), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR14), .QN());
  DFFR_X1 P3_Datao_PTR15 ( .D(_03409__PTR271), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR15), .QN());
  DFFR_X1 P3_Datao_PTR16 ( .D(_03409__PTR272), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR16), .QN());
  DFFR_X1 P3_Datao_PTR17 ( .D(_03409__PTR273), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR17), .QN());
  DFFR_X1 P3_Datao_PTR18 ( .D(_03409__PTR274), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR18), .QN());
  DFFR_X1 P3_Datao_PTR19 ( .D(_03409__PTR275), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR19), .QN());
  DFFR_X1 P3_Datao_PTR20 ( .D(_03409__PTR276), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR20), .QN());
  DFFR_X1 P3_Datao_PTR21 ( .D(_03409__PTR277), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR21), .QN());
  DFFR_X1 P3_Datao_PTR22 ( .D(_03409__PTR278), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR22), .QN());
  DFFR_X1 P3_Datao_PTR23 ( .D(_03409__PTR279), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR23), .QN());
  DFFR_X1 P3_Datao_PTR24 ( .D(_03409__PTR280), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR24), .QN());
  DFFR_X1 P3_Datao_PTR25 ( .D(_03409__PTR281), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR25), .QN());
  DFFR_X1 P3_Datao_PTR26 ( .D(_03409__PTR282), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR26), .QN());
  DFFR_X1 P3_Datao_PTR27 ( .D(_03409__PTR283), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR27), .QN());
  DFFR_X1 P3_Datao_PTR28 ( .D(_03409__PTR284), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR28), .QN());
  DFFR_X1 P3_Datao_PTR29 ( .D(_03409__PTR285), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR29), .QN());
  DFFR_X1 P3_Datao_PTR30 ( .D(_03409__PTR286), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR30), .QN());
  DFFR_X1 P3_DataWidth_reg_PTR0 ( .D(_02460__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR0), .QN());
  BUF_X1 U67 ( .A(P3_DataWidth_reg_PTR0), .Z(P3_DataWidth_PTR0) );
  DFFR_X1 P3_DataWidth_reg_PTR2 ( .D(_02460__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR2), .QN());
  BUF_X1 U68 ( .A(P3_DataWidth_reg_PTR2), .Z(P3_DataWidth_PTR2) );
  DFFR_X1 P3_DataWidth_reg_PTR3 ( .D(_02460__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR3), .QN());
  BUF_X1 U69 ( .A(P3_DataWidth_reg_PTR3), .Z(P3_DataWidth_PTR3) );
  DFFR_X1 P3_DataWidth_reg_PTR4 ( .D(_02460__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR4), .QN());
  BUF_X1 U70 ( .A(P3_DataWidth_reg_PTR4), .Z(P3_DataWidth_PTR4) );
  DFFR_X1 P3_DataWidth_reg_PTR5 ( .D(_02460__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR5), .QN());
  BUF_X1 U71 ( .A(P3_DataWidth_reg_PTR5), .Z(P3_DataWidth_PTR5) );
  DFFR_X1 P3_DataWidth_reg_PTR6 ( .D(_02460__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR6), .QN());
  BUF_X1 U72 ( .A(P3_DataWidth_reg_PTR6), .Z(P3_DataWidth_PTR6) );
  DFFR_X1 P3_DataWidth_reg_PTR7 ( .D(_02460__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR7), .QN());
  BUF_X1 U73 ( .A(P3_DataWidth_reg_PTR7), .Z(P3_DataWidth_PTR7) );
  DFFR_X1 P3_DataWidth_reg_PTR8 ( .D(_02460__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR8), .QN());
  BUF_X1 U74 ( .A(P3_DataWidth_reg_PTR8), .Z(P3_DataWidth_PTR8) );
  DFFR_X1 P3_DataWidth_reg_PTR9 ( .D(_02460__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR9), .QN());
  BUF_X1 U75 ( .A(P3_DataWidth_reg_PTR9), .Z(P3_DataWidth_PTR9) );
  DFFR_X1 P3_DataWidth_reg_PTR10 ( .D(_02460__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR10), .QN());
  BUF_X1 U76 ( .A(P3_DataWidth_reg_PTR10), .Z(P3_DataWidth_PTR10) );
  DFFR_X1 P3_DataWidth_reg_PTR11 ( .D(_02460__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR11), .QN());
  BUF_X1 U77 ( .A(P3_DataWidth_reg_PTR11), .Z(P3_DataWidth_PTR11) );
  DFFR_X1 P3_DataWidth_reg_PTR12 ( .D(_02460__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR12), .QN());
  BUF_X1 U78 ( .A(P3_DataWidth_reg_PTR12), .Z(P3_DataWidth_PTR12) );
  DFFR_X1 P3_DataWidth_reg_PTR13 ( .D(_02460__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR13), .QN());
  BUF_X1 U79 ( .A(P3_DataWidth_reg_PTR13), .Z(P3_DataWidth_PTR13) );
  DFFR_X1 P3_DataWidth_reg_PTR14 ( .D(_02460__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR14), .QN());
  BUF_X1 U80 ( .A(P3_DataWidth_reg_PTR14), .Z(P3_DataWidth_PTR14) );
  DFFR_X1 P3_DataWidth_reg_PTR15 ( .D(_02460__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR15), .QN());
  BUF_X1 U81 ( .A(P3_DataWidth_reg_PTR15), .Z(P3_DataWidth_PTR15) );
  DFFR_X1 P3_DataWidth_reg_PTR16 ( .D(_02460__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR16), .QN());
  BUF_X1 U82 ( .A(P3_DataWidth_reg_PTR16), .Z(P3_DataWidth_PTR16) );
  DFFR_X1 P3_DataWidth_reg_PTR17 ( .D(_02460__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR17), .QN());
  BUF_X1 U83 ( .A(P3_DataWidth_reg_PTR17), .Z(P3_DataWidth_PTR17) );
  DFFR_X1 P3_DataWidth_reg_PTR18 ( .D(_02460__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR18), .QN());
  BUF_X1 U84 ( .A(P3_DataWidth_reg_PTR18), .Z(P3_DataWidth_PTR18) );
  DFFR_X1 P3_DataWidth_reg_PTR19 ( .D(_02460__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR19), .QN());
  BUF_X1 U85 ( .A(P3_DataWidth_reg_PTR19), .Z(P3_DataWidth_PTR19) );
  DFFR_X1 P3_DataWidth_reg_PTR20 ( .D(_02460__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR20), .QN());
  BUF_X1 U86 ( .A(P3_DataWidth_reg_PTR20), .Z(P3_DataWidth_PTR20) );
  DFFR_X1 P3_DataWidth_reg_PTR21 ( .D(_02460__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR21), .QN());
  BUF_X1 U87 ( .A(P3_DataWidth_reg_PTR21), .Z(P3_DataWidth_PTR21) );
  DFFR_X1 P3_DataWidth_reg_PTR22 ( .D(_02460__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR22), .QN());
  BUF_X1 U88 ( .A(P3_DataWidth_reg_PTR22), .Z(P3_DataWidth_PTR22) );
  DFFR_X1 P3_DataWidth_reg_PTR23 ( .D(_02460__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR23), .QN());
  BUF_X1 U89 ( .A(P3_DataWidth_reg_PTR23), .Z(P3_DataWidth_PTR23) );
  DFFR_X1 P3_DataWidth_reg_PTR24 ( .D(_02460__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR24), .QN());
  BUF_X1 U90 ( .A(P3_DataWidth_reg_PTR24), .Z(P3_DataWidth_PTR24) );
  DFFR_X1 P3_DataWidth_reg_PTR25 ( .D(_02460__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR25), .QN());
  BUF_X1 U91 ( .A(P3_DataWidth_reg_PTR25), .Z(P3_DataWidth_PTR25) );
  DFFR_X1 P3_DataWidth_reg_PTR26 ( .D(_02460__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR26), .QN());
  BUF_X1 U92 ( .A(P3_DataWidth_reg_PTR26), .Z(P3_DataWidth_PTR26) );
  DFFR_X1 P3_DataWidth_reg_PTR27 ( .D(_02460__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR27), .QN());
  BUF_X1 U93 ( .A(P3_DataWidth_reg_PTR27), .Z(P3_DataWidth_PTR27) );
  DFFR_X1 P3_DataWidth_reg_PTR28 ( .D(_02460__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR28), .QN());
  BUF_X1 U94 ( .A(P3_DataWidth_reg_PTR28), .Z(P3_DataWidth_PTR28) );
  DFFR_X1 P3_DataWidth_reg_PTR29 ( .D(_02460__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR29), .QN());
  BUF_X1 U95 ( .A(P3_DataWidth_reg_PTR29), .Z(P3_DataWidth_PTR29) );
  DFFR_X1 P3_DataWidth_reg_PTR30 ( .D(_02460__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR30), .QN());
  BUF_X1 U96 ( .A(P3_DataWidth_reg_PTR30), .Z(P3_DataWidth_PTR30) );
  DFFR_X1 P3_State_PTR0 ( .D(_02459__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_State_PTR0), .QN());
  DFFR_X1 P3_State_PTR1 ( .D(_02459__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_State_PTR1), .QN());
  DFFR_X1 P3_Address_PTR0 ( .D(_02462__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR0), .QN());
  DFFR_X1 P3_Address_PTR1 ( .D(_02462__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR1), .QN());
  DFFR_X1 P3_Address_PTR2 ( .D(_02462__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR2), .QN());
  DFFR_X1 P3_Address_PTR3 ( .D(_02462__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR3), .QN());
  DFFR_X1 P3_Address_PTR4 ( .D(_02462__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR4), .QN());
  DFFR_X1 P3_Address_PTR5 ( .D(_02462__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR5), .QN());
  DFFR_X1 P3_Address_PTR6 ( .D(_02462__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR6), .QN());
  DFFR_X1 P3_Address_PTR7 ( .D(_02462__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR7), .QN());
  DFFR_X1 P3_Address_PTR8 ( .D(_02462__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR8), .QN());
  DFFR_X1 P3_Address_PTR9 ( .D(_02462__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR9), .QN());
  DFFR_X1 P3_Address_PTR10 ( .D(_02462__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR10), .QN());
  DFFR_X1 P3_Address_PTR11 ( .D(_02462__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR11), .QN());
  DFFR_X1 P3_Address_PTR12 ( .D(_02462__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR12), .QN());
  DFFR_X1 P3_Address_PTR13 ( .D(_02462__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR13), .QN());
  DFFR_X1 P3_Address_PTR14 ( .D(_02462__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR14), .QN());
  DFFR_X1 P3_Address_PTR15 ( .D(_02462__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR15), .QN());
  DFFR_X1 P3_Address_PTR16 ( .D(_02462__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR16), .QN());
  DFFR_X1 P3_Address_PTR17 ( .D(_02462__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR17), .QN());
  DFFR_X1 P3_Address_PTR18 ( .D(_02462__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR18), .QN());
  DFFR_X1 P3_Address_PTR19 ( .D(_02462__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR19), .QN());
  DFFR_X1 P3_Address_PTR20 ( .D(_02462__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR20), .QN());
  DFFR_X1 P3_Address_PTR21 ( .D(_02462__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR21), .QN());
  DFFR_X1 P3_Address_PTR22 ( .D(_02462__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR22), .QN());
  DFFR_X1 P3_Address_PTR23 ( .D(_02462__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR23), .QN());
  DFFR_X1 P3_Address_PTR24 ( .D(_02462__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR24), .QN());
  DFFR_X1 P3_Address_PTR25 ( .D(_02462__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR25), .QN());
  DFFR_X1 P3_Address_PTR26 ( .D(_02462__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR26), .QN());
  DFFR_X1 P3_Address_PTR27 ( .D(_02462__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR27), .QN());
  DFFR_X1 P3_Address_PTR28 ( .D(_02462__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Address_PTR28), .QN());
  DFFR_X1 P3_P1_uWord_PTR0 ( .D(_02517__PTR80), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR0), .QN());
  DFFR_X1 P3_P1_uWord_PTR1 ( .D(_02517__PTR81), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR1), .QN());
  DFFR_X1 P3_P1_uWord_PTR2 ( .D(_02517__PTR82), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR2), .QN());
  DFFR_X1 P3_P1_uWord_PTR3 ( .D(_02517__PTR83), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR3), .QN());
  DFFR_X1 P3_P1_uWord_PTR4 ( .D(_02517__PTR84), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR4), .QN());
  DFFR_X1 P3_P1_uWord_PTR5 ( .D(_02517__PTR85), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR5), .QN());
  DFFR_X1 P3_P1_uWord_PTR6 ( .D(_02517__PTR86), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR6), .QN());
  DFFR_X1 P3_P1_uWord_PTR7 ( .D(_02517__PTR87), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR7), .QN());
  DFFR_X1 P3_P1_uWord_PTR8 ( .D(_02517__PTR88), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR8), .QN());
  DFFR_X1 P3_P1_uWord_PTR9 ( .D(_02517__PTR89), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR9), .QN());
  DFFR_X1 P3_P1_uWord_PTR10 ( .D(_02517__PTR90), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR10), .QN());
  DFFR_X1 P3_P1_uWord_PTR11 ( .D(_02517__PTR91), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR11), .QN());
  DFFR_X1 P3_P1_uWord_PTR12 ( .D(_02517__PTR92), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR12), .QN());
  DFFR_X1 P3_P1_uWord_PTR13 ( .D(_02517__PTR93), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_uWord_PTR13), .QN());
  DFFR_X1 P3_P1_lWord_PTR0 ( .D(_02518__PTR80), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR0), .QN());
  DFFR_X1 P3_P1_lWord_PTR1 ( .D(_02518__PTR81), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR1), .QN());
  DFFR_X1 P3_P1_lWord_PTR2 ( .D(_02518__PTR82), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR2), .QN());
  DFFR_X1 P3_P1_lWord_PTR3 ( .D(_02518__PTR83), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR3), .QN());
  DFFR_X1 P3_P1_lWord_PTR4 ( .D(_02518__PTR84), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR4), .QN());
  DFFR_X1 P3_P1_lWord_PTR5 ( .D(_02518__PTR85), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR5), .QN());
  DFFR_X1 P3_P1_lWord_PTR6 ( .D(_02518__PTR86), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR6), .QN());
  DFFR_X1 P3_P1_lWord_PTR7 ( .D(_02518__PTR87), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR7), .QN());
  DFFR_X1 P3_P1_lWord_PTR8 ( .D(_02518__PTR88), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR8), .QN());
  DFFR_X1 P3_P1_lWord_PTR9 ( .D(_02518__PTR89), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR9), .QN());
  DFFR_X1 P3_P1_lWord_PTR10 ( .D(_02518__PTR90), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR10), .QN());
  DFFR_X1 P3_P1_lWord_PTR11 ( .D(_02518__PTR91), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR11), .QN());
  DFFR_X1 P3_P1_lWord_PTR12 ( .D(_02518__PTR92), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR12), .QN());
  DFFR_X1 P3_P1_lWord_PTR13 ( .D(_02518__PTR93), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR13), .QN());
  DFFR_X1 P3_P1_lWord_PTR14 ( .D(_02518__PTR94), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_lWord_PTR14), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR0 ( .D(_03343__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR0), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR1 ( .D(_03343__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR1), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR2 ( .D(_03343__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR2), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR3 ( .D(_03343__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR3), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR4 ( .D(_03343__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR4), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR5 ( .D(_03343__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR5), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR6 ( .D(_03343__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR6), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR7 ( .D(_03343__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR7), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR8 ( .D(_03343__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR8), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR9 ( .D(_03343__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR9), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR10 ( .D(_03343__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR10), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR11 ( .D(_03343__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR11), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR12 ( .D(_03343__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR12), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR13 ( .D(_03343__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR13), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR14 ( .D(_03343__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR14), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR15 ( .D(_03343__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR15), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR16 ( .D(_03343__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR16), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR17 ( .D(_03343__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR17), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR18 ( .D(_03343__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR18), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR19 ( .D(_03343__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR19), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR20 ( .D(_03343__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR20), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR21 ( .D(_03343__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR21), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR22 ( .D(_03343__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR22), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR23 ( .D(_03343__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR23), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR24 ( .D(_03343__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR24), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR25 ( .D(_03343__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR25), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR26 ( .D(_03343__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR26), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR27 ( .D(_03343__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR27), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR28 ( .D(_03343__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR28), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR29 ( .D(_03343__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR29), .QN());
  DFFR_X1 P3_P1_PhyAddrPointer_PTR30 ( .D(_03343__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_PhyAddrPointer_PTR30), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR0 ( .D(_03346__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR0), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR1 ( .D(_03346__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR1), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR2 ( .D(_03346__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR2), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR3 ( .D(_03346__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR3), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR4 ( .D(_03346__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR4), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR5 ( .D(_03346__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR5), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR6 ( .D(_03346__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR6), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR7 ( .D(_03346__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR7), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR8 ( .D(_03346__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR8), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR9 ( .D(_03346__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR9), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR10 ( .D(_03346__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR10), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR11 ( .D(_03346__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR11), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR12 ( .D(_03346__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR12), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR13 ( .D(_03346__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR13), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR14 ( .D(_03346__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR14), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR15 ( .D(_03346__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR15), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR16 ( .D(_03346__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR16), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR17 ( .D(_03346__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR17), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR18 ( .D(_03346__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR18), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR19 ( .D(_03346__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR19), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR20 ( .D(_03346__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR20), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR21 ( .D(_03346__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR21), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR22 ( .D(_03346__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR22), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR23 ( .D(_03346__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR23), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR24 ( .D(_03346__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR24), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR25 ( .D(_03346__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR25), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR26 ( .D(_03346__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR26), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR27 ( .D(_03346__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR27), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR28 ( .D(_03346__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR28), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR29 ( .D(_03346__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR29), .QN());
  DFFR_X1 P3_P1_InstAddrPointer_PTR30 ( .D(_03346__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstAddrPointer_PTR30), .QN());
  DFFR_X1 P3_P1_InstQueueWr_Addr_PTR0 ( .D(_02512__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueueWr_Addr_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueueWr_Addr_PTR1 ( .D(_02512__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueueWr_Addr_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueueWr_Addr_PTR2 ( .D(_02512__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueueWr_Addr_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueueWr_Addr_PTR3 ( .D(_02512__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueueWr_Addr_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueueRd_Addr_PTR0 ( .D(_02514__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueueRd_Addr_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueueRd_Addr_PTR1 ( .D(_02514__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueueRd_Addr_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueueRd_Addr_PTR2 ( .D(_02514__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueueRd_Addr_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueueRd_Addr_PTR3 ( .D(_02514__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueueRd_Addr_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR0_PTR0 ( .D(_02510__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR0_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR0_PTR1 ( .D(_02510__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR0_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR0_PTR2 ( .D(_02510__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR0_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR0_PTR3 ( .D(_02510__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR0_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR0_PTR4 ( .D(_02510__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR0_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR0_PTR5 ( .D(_02510__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR0_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR0_PTR6 ( .D(_02510__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR0_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR1_PTR0 ( .D(_02508__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR1_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR1_PTR1 ( .D(_02508__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR1_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR1_PTR2 ( .D(_02508__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR1_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR1_PTR3 ( .D(_02508__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR1_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR1_PTR4 ( .D(_02508__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR1_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR1_PTR5 ( .D(_02508__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR1_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR1_PTR6 ( .D(_02508__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR1_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR2_PTR0 ( .D(_02506__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR2_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR2_PTR1 ( .D(_02506__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR2_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR2_PTR2 ( .D(_02506__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR2_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR2_PTR3 ( .D(_02506__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR2_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR2_PTR4 ( .D(_02506__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR2_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR2_PTR5 ( .D(_02506__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR2_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR2_PTR6 ( .D(_02506__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR2_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR3_PTR0 ( .D(_02504__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR3_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR3_PTR1 ( .D(_02504__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR3_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR3_PTR2 ( .D(_02504__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR3_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR3_PTR3 ( .D(_02504__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR3_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR3_PTR4 ( .D(_02504__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR3_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR3_PTR5 ( .D(_02504__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR3_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR3_PTR6 ( .D(_02504__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR3_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR4_PTR0 ( .D(_02502__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR4_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR4_PTR1 ( .D(_02502__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR4_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR4_PTR2 ( .D(_02502__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR4_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR4_PTR3 ( .D(_02502__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR4_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR4_PTR4 ( .D(_02502__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR4_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR4_PTR5 ( .D(_02502__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR4_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR4_PTR6 ( .D(_02502__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR4_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR5_PTR0 ( .D(_02500__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR5_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR5_PTR1 ( .D(_02500__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR5_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR5_PTR2 ( .D(_02500__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR5_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR5_PTR3 ( .D(_02500__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR5_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR5_PTR4 ( .D(_02500__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR5_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR5_PTR5 ( .D(_02500__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR5_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR5_PTR6 ( .D(_02500__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR5_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR6_PTR0 ( .D(_02498__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR6_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR6_PTR1 ( .D(_02498__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR6_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR6_PTR2 ( .D(_02498__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR6_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR6_PTR3 ( .D(_02498__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR6_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR6_PTR4 ( .D(_02498__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR6_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR6_PTR5 ( .D(_02498__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR6_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR6_PTR6 ( .D(_02498__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR6_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR7_PTR0 ( .D(_02496__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR7_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR7_PTR1 ( .D(_02496__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR7_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR7_PTR2 ( .D(_02496__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR7_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR7_PTR3 ( .D(_02496__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR7_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR7_PTR4 ( .D(_02496__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR7_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR7_PTR5 ( .D(_02496__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR7_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR7_PTR6 ( .D(_02496__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR7_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR8_PTR0 ( .D(_02494__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR8_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR8_PTR1 ( .D(_02494__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR8_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR8_PTR2 ( .D(_02494__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR8_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR8_PTR3 ( .D(_02494__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR8_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR8_PTR4 ( .D(_02494__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR8_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR8_PTR5 ( .D(_02494__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR8_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR8_PTR6 ( .D(_02494__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR8_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR9_PTR0 ( .D(_02492__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR9_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR9_PTR1 ( .D(_02492__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR9_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR9_PTR2 ( .D(_02492__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR9_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR9_PTR3 ( .D(_02492__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR9_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR9_PTR4 ( .D(_02492__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR9_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR9_PTR5 ( .D(_02492__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR9_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR9_PTR6 ( .D(_02492__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR9_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR10_PTR0 ( .D(_02490__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR10_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR10_PTR1 ( .D(_02490__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR10_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR10_PTR2 ( .D(_02490__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR10_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR10_PTR3 ( .D(_02490__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR10_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR10_PTR4 ( .D(_02490__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR10_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR10_PTR5 ( .D(_02490__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR10_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR10_PTR6 ( .D(_02490__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR10_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR11_PTR0 ( .D(_02488__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR11_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR11_PTR1 ( .D(_02488__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR11_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR11_PTR2 ( .D(_02488__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR11_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR11_PTR3 ( .D(_02488__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR11_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR11_PTR4 ( .D(_02488__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR11_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR11_PTR5 ( .D(_02488__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR11_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR11_PTR6 ( .D(_02488__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR11_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR12_PTR0 ( .D(_02486__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR12_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR12_PTR1 ( .D(_02486__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR12_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR12_PTR2 ( .D(_02486__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR12_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR12_PTR3 ( .D(_02486__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR12_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR12_PTR4 ( .D(_02486__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR12_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR12_PTR5 ( .D(_02486__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR12_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR12_PTR6 ( .D(_02486__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR12_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR13_PTR0 ( .D(_02484__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR13_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR13_PTR1 ( .D(_02484__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR13_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR13_PTR2 ( .D(_02484__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR13_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR13_PTR3 ( .D(_02484__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR13_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR13_PTR4 ( .D(_02484__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR13_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR13_PTR5 ( .D(_02484__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR13_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR13_PTR6 ( .D(_02484__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR13_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR14_PTR0 ( .D(_02482__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR14_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR14_PTR1 ( .D(_02482__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR14_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR14_PTR2 ( .D(_02482__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR14_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR14_PTR3 ( .D(_02482__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR14_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR14_PTR4 ( .D(_02482__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR14_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR14_PTR5 ( .D(_02482__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR14_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR14_PTR6 ( .D(_02482__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR14_PTR6), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR15_PTR0 ( .D(_02480__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR15_PTR0), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR15_PTR1 ( .D(_02480__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR15_PTR1), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR15_PTR2 ( .D(_02480__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR15_PTR2), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR15_PTR3 ( .D(_02480__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR15_PTR3), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR15_PTR4 ( .D(_02480__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR15_PTR4), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR15_PTR5 ( .D(_02480__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR15_PTR5), .QN());
  DFFR_X1 P3_P1_InstQueue_PTR15_PTR6 ( .D(_02480__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_InstQueue_PTR15_PTR6), .QN());
  DFFR_X1 P3_P1_State2_PTR0 ( .D(_02476__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_State2_PTR0), .QN());
  DFFR_X1 P3_P1_State2_PTR1 ( .D(_02476__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_State2_PTR1), .QN());
  DFFR_X1 P3_P1_State2_PTR2 ( .D(_02476__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_P1_State2_PTR2), .QN());
  DFFR_X1 P3_DataWidth_reg_PTR31 ( .D(_02460__PTR32), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_DataWidth_reg_PTR31), .QN());
  BUF_X1 U97 ( .A(P3_DataWidth_reg_PTR31), .Z(P3_DataWidth_PTR31) );
  DFFR_X1 P3_Datao_PTR31 ( .D(_03409__PTR288), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_Datao_PTR31), .QN());
  DFFR_X1 P3_rEIP_PTR31 ( .D(_02478__PTR32), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_rEIP_PTR31), .QN());
  DFFR_X1 P2_DataWidth_reg_PTR31 ( .D(_02171__PTR32), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_DataWidth_reg_PTR31), .QN());
  BUF_X1 U98 ( .A(P2_DataWidth_reg_PTR31), .Z(P2_DataWidth_PTR31) );
  DFFR_X1 P2_Datao_PTR31 ( .D(_03164__PTR288), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_Datao_PTR31), .QN());
  DFFR_X1 P2_rEIP_PTR31 ( .D(_02189__PTR32), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_rEIP_PTR31), .QN());
  DFFR_X1 P1_DataWidth_reg_PTR31 ( .D(_01879__PTR32), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_DataWidth_reg_PTR31), .QN());
  BUF_X1 U99 ( .A(P1_DataWidth_reg_PTR31), .Z(P1_DataWidth_PTR31) );
  DFFR_X1 P1_Datao_PTR31 ( .D(_02919__PTR288), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_Datao_PTR31), .QN());
  DFFR_X1 P1_rEIP_PTR31 ( .D(_01897__PTR32), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_rEIP_PTR31), .QN());
  DFFR_X1 P3_BE_n_PTR3 ( .D(P3_ByteEnable_PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_BE_n_PTR3), .QN());
  DFFR_X1 P3_BE_n_PTR2 ( .D(P3_ByteEnable_PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_BE_n_PTR2), .QN());
  DFFR_X1 P3_BE_n_PTR1 ( .D(P3_ByteEnable_PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_BE_n_PTR1), .QN());
  DFFR_X1 P3_BE_n_PTR0 ( .D(P3_ByteEnable_PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_BE_n_PTR0), .QN());
  DFFR_X1 P3_W_R_n ( .D(_02428__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_W_R_n), .QN());
  DFFR_X1 P3_M_IO_n ( .D(P3_MemoryFetch), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_M_IO_n), .QN());
  DFFR_X1 P2_BE_n_PTR3 ( .D(P2_ByteEnable_PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_BE_n_PTR3), .QN());
  DFFR_X1 P2_BE_n_PTR2 ( .D(P2_ByteEnable_PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_BE_n_PTR2), .QN());
  DFFR_X1 P2_BE_n_PTR1 ( .D(P2_ByteEnable_PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_BE_n_PTR1), .QN());
  DFFR_X1 P2_BE_n_PTR0 ( .D(P2_ByteEnable_PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_BE_n_PTR0), .QN());
  DFFR_X1 P2_W_R_n ( .D(_02139__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_W_R_n), .QN());
  DFFR_X1 P2_M_IO_n ( .D(P2_MemoryFetch), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_M_IO_n), .QN());
  DFFR_X1 P1_BE_n_PTR3 ( .D(P1_ByteEnable_PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_BE_n_PTR3), .QN());
  DFFR_X1 P1_BE_n_PTR2 ( .D(P1_ByteEnable_PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_BE_n_PTR2), .QN());
  DFFR_X1 P1_BE_n_PTR1 ( .D(P1_ByteEnable_PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_BE_n_PTR1), .QN());
  DFFR_X1 P1_BE_n_PTR0 ( .D(P1_ByteEnable_PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_BE_n_PTR0), .QN());
  DFFR_X1 P1_W_R_n ( .D(_01846__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_W_R_n), .QN());
  DFFR_X1 P1_M_IO_n ( .D(P1_MemoryFetch), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_M_IO_n), .QN());
  INV_X1 U100 ( .A(_01883__PTR0), .ZN(_00267_) );
  INV_X1 U101 ( .A(_01883__PTR3), .ZN(_00268_) );
  INV_X1 U102 ( .A(_01883__PTR1), .ZN(_00262_) );
  INV_X1 U103 ( .A(_01883__PTR2), .ZN(_00263_) );
  INV_X1 U104 ( .A(_01883__PTR5), .ZN(_00264_) );
  INV_X1 U105 ( .A(_01883__PTR6), .ZN(_00265_) );
  INV_X1 U106 ( .A(_01883__PTR4), .ZN(_00269_) );
  INV_X1 U107 ( .A(_01883__PTR7), .ZN(_00266_) );
  INV_X1 U108 ( .A(P2_Datao_PTR16), .ZN(_05726__PTR16) );
  INV_X1 U109 ( .A(P2_Datao_PTR17), .ZN(_05726__PTR17) );
  INV_X1 U110 ( .A(P2_Datao_PTR18), .ZN(_05726__PTR18) );
  INV_X1 U111 ( .A(P2_Datao_PTR19), .ZN(_05726__PTR19) );
  INV_X1 U112 ( .A(P2_Datao_PTR20), .ZN(_05726__PTR20) );
  INV_X1 U113 ( .A(P2_Datao_PTR21), .ZN(_05726__PTR21) );
  INV_X1 U114 ( .A(P2_Datao_PTR22), .ZN(_05726__PTR22) );
  INV_X1 U115 ( .A(P2_Datao_PTR23), .ZN(_05726__PTR23) );
  INV_X1 U116 ( .A(P2_Datao_PTR24), .ZN(_05726__PTR24) );
  INV_X1 U117 ( .A(P2_Datao_PTR25), .ZN(_05726__PTR25) );
  INV_X1 U118 ( .A(P2_Datao_PTR26), .ZN(_05726__PTR26) );
  INV_X1 U119 ( .A(P2_Datao_PTR27), .ZN(_05726__PTR27) );
  INV_X1 U120 ( .A(P2_Datao_PTR28), .ZN(_05726__PTR28) );
  INV_X1 U121 ( .A(P2_Datao_PTR29), .ZN(_05726__PTR29) );
  INV_X1 U122 ( .A(P2_Datao_PTR8), .ZN(_05726__PTR8) );
  INV_X1 U123 ( .A(P2_Datao_PTR9), .ZN(_05726__PTR9) );
  INV_X1 U124 ( .A(P2_Datao_PTR10), .ZN(_05726__PTR10) );
  INV_X1 U125 ( .A(P2_Datao_PTR11), .ZN(_05726__PTR11) );
  INV_X1 U126 ( .A(P2_Datao_PTR12), .ZN(_05726__PTR12) );
  INV_X1 U127 ( .A(P2_Datao_PTR13), .ZN(_05726__PTR13) );
  INV_X1 U128 ( .A(P2_Datao_PTR14), .ZN(_05726__PTR14) );
  INV_X1 U129 ( .A(P2_Datao_PTR15), .ZN(_05726__PTR15) );
  INV_X1 U130 ( .A(P2_Datao_PTR4), .ZN(_05726__PTR4) );
  INV_X1 U131 ( .A(P2_Datao_PTR5), .ZN(_05726__PTR5) );
  INV_X1 U132 ( .A(P2_Datao_PTR6), .ZN(_05726__PTR6) );
  INV_X1 U133 ( .A(P2_Datao_PTR7), .ZN(_05726__PTR7) );
  INV_X1 U134 ( .A(P2_Datao_PTR2), .ZN(_05726__PTR2) );
  INV_X1 U135 ( .A(P2_Datao_PTR3), .ZN(_05726__PTR3) );
  INV_X1 U136 ( .A(P1_Datao_PTR16), .ZN(_05722__PTR16) );
  INV_X1 U137 ( .A(P1_Datao_PTR17), .ZN(_05722__PTR17) );
  INV_X1 U138 ( .A(P1_Datao_PTR18), .ZN(_05722__PTR18) );
  INV_X1 U139 ( .A(P1_Datao_PTR19), .ZN(_05722__PTR19) );
  INV_X1 U140 ( .A(P1_Datao_PTR20), .ZN(_05722__PTR20) );
  INV_X1 U141 ( .A(P1_Datao_PTR21), .ZN(_05722__PTR21) );
  INV_X1 U142 ( .A(P1_Datao_PTR22), .ZN(_05722__PTR22) );
  INV_X1 U143 ( .A(P1_Datao_PTR23), .ZN(_05722__PTR23) );
  INV_X1 U144 ( .A(P1_Datao_PTR24), .ZN(_05722__PTR24) );
  INV_X1 U145 ( .A(P1_Datao_PTR25), .ZN(_05722__PTR25) );
  INV_X1 U146 ( .A(P1_Datao_PTR26), .ZN(_05722__PTR26) );
  INV_X1 U147 ( .A(P1_Datao_PTR27), .ZN(_05722__PTR27) );
  INV_X1 U148 ( .A(P1_Datao_PTR28), .ZN(_05722__PTR28) );
  INV_X1 U149 ( .A(P1_Datao_PTR29), .ZN(_05722__PTR29) );
  INV_X1 U150 ( .A(P1_Datao_PTR8), .ZN(_05722__PTR8) );
  INV_X1 U151 ( .A(P1_Datao_PTR9), .ZN(_05722__PTR9) );
  INV_X1 U152 ( .A(P1_Datao_PTR10), .ZN(_05722__PTR10) );
  INV_X1 U153 ( .A(P1_Datao_PTR11), .ZN(_05722__PTR11) );
  INV_X1 U154 ( .A(P1_Datao_PTR12), .ZN(_05722__PTR12) );
  INV_X1 U155 ( .A(P1_Datao_PTR13), .ZN(_05722__PTR13) );
  INV_X1 U156 ( .A(P1_Datao_PTR14), .ZN(_05722__PTR14) );
  INV_X1 U157 ( .A(P1_Datao_PTR15), .ZN(_05722__PTR15) );
  INV_X1 U158 ( .A(P1_Datao_PTR4), .ZN(_05722__PTR4) );
  INV_X1 U159 ( .A(P1_Datao_PTR5), .ZN(_05722__PTR5) );
  INV_X1 U160 ( .A(P1_Datao_PTR6), .ZN(_05722__PTR6) );
  INV_X1 U161 ( .A(P1_Datao_PTR7), .ZN(_05722__PTR7) );
  INV_X1 U162 ( .A(P1_Datao_PTR2), .ZN(_05722__PTR2) );
  INV_X1 U163 ( .A(P1_Datao_PTR3), .ZN(_05722__PTR3) );
  INV_X1 U164 ( .A(P3_Datao_PTR16), .ZN(_05730__PTR16) );
  INV_X1 U165 ( .A(P3_Datao_PTR17), .ZN(_05730__PTR17) );
  INV_X1 U166 ( .A(P3_Datao_PTR18), .ZN(_05730__PTR18) );
  INV_X1 U167 ( .A(P3_Datao_PTR19), .ZN(_05730__PTR19) );
  INV_X1 U168 ( .A(P3_Datao_PTR20), .ZN(_05730__PTR20) );
  INV_X1 U169 ( .A(P3_Datao_PTR21), .ZN(_05730__PTR21) );
  INV_X1 U170 ( .A(P3_Datao_PTR22), .ZN(_05730__PTR22) );
  INV_X1 U171 ( .A(P3_Datao_PTR23), .ZN(_05730__PTR23) );
  INV_X1 U172 ( .A(P3_Datao_PTR24), .ZN(_05730__PTR24) );
  INV_X1 U173 ( .A(P3_Datao_PTR25), .ZN(_05730__PTR25) );
  INV_X1 U174 ( .A(P3_Datao_PTR26), .ZN(_05730__PTR26) );
  INV_X1 U175 ( .A(P3_Datao_PTR27), .ZN(_05730__PTR27) );
  INV_X1 U176 ( .A(P3_Datao_PTR28), .ZN(_05730__PTR28) );
  INV_X1 U177 ( .A(P3_Datao_PTR29), .ZN(_05730__PTR29) );
  INV_X1 U178 ( .A(P3_Datao_PTR8), .ZN(_05730__PTR8) );
  INV_X1 U179 ( .A(P3_Datao_PTR9), .ZN(_05730__PTR9) );
  INV_X1 U180 ( .A(P3_Datao_PTR10), .ZN(_05730__PTR10) );
  INV_X1 U181 ( .A(P3_Datao_PTR11), .ZN(_05730__PTR11) );
  INV_X1 U182 ( .A(P3_Datao_PTR12), .ZN(_05730__PTR12) );
  INV_X1 U183 ( .A(P3_Datao_PTR13), .ZN(_05730__PTR13) );
  INV_X1 U184 ( .A(P3_Datao_PTR14), .ZN(_05730__PTR14) );
  INV_X1 U185 ( .A(P3_Datao_PTR15), .ZN(_05730__PTR15) );
  INV_X1 U186 ( .A(P3_Datao_PTR4), .ZN(_05730__PTR4) );
  INV_X1 U187 ( .A(P3_Datao_PTR5), .ZN(_05730__PTR5) );
  INV_X1 U188 ( .A(P3_Datao_PTR6), .ZN(_05730__PTR6) );
  INV_X1 U189 ( .A(P3_Datao_PTR7), .ZN(_05730__PTR7) );
  INV_X1 U190 ( .A(P3_Datao_PTR2), .ZN(_05730__PTR2) );
  INV_X1 U191 ( .A(P3_Datao_PTR3), .ZN(_05730__PTR3) );
  INV_X1 U192 ( .A(_02175__PTR1), .ZN(_00270_) );
  INV_X1 U193 ( .A(_02175__PTR2), .ZN(_00273_) );
  INV_X1 U194 ( .A(_02175__PTR5), .ZN(_00272_) );
  INV_X1 U195 ( .A(_02175__PTR6), .ZN(_00259_) );
  INV_X1 U196 ( .A(_02175__PTR4), .ZN(_00261_) );
  INV_X1 U197 ( .A(_02175__PTR7), .ZN(_00260_) );
  INV_X1 U198 ( .A(_02175__PTR0), .ZN(_00274_) );
  INV_X1 U199 ( .A(_02175__PTR3), .ZN(_00271_) );
  INV_X1 U200 ( .A(P1_P1_InstQueueRd_Addr_PTR0), .ZN(_01884__PTR3) );
  INV_X1 U201 ( .A(P1_P1_InstAddrPointer_PTR16), .ZN(_02745__PTR16) );
  INV_X1 U202 ( .A(P1_P1_InstAddrPointer_PTR17), .ZN(_02745__PTR17) );
  INV_X1 U203 ( .A(P1_P1_InstAddrPointer_PTR18), .ZN(_02745__PTR18) );
  INV_X1 U204 ( .A(P1_P1_InstAddrPointer_PTR19), .ZN(_02745__PTR19) );
  INV_X1 U205 ( .A(P1_P1_InstAddrPointer_PTR20), .ZN(_02745__PTR20) );
  INV_X1 U206 ( .A(P1_P1_InstAddrPointer_PTR21), .ZN(_02745__PTR21) );
  INV_X1 U207 ( .A(P1_P1_InstAddrPointer_PTR22), .ZN(_02745__PTR22) );
  INV_X1 U208 ( .A(P1_P1_InstAddrPointer_PTR23), .ZN(_02745__PTR23) );
  INV_X1 U209 ( .A(P1_P1_InstAddrPointer_PTR24), .ZN(_02745__PTR24) );
  INV_X1 U210 ( .A(P1_P1_InstAddrPointer_PTR25), .ZN(_02745__PTR25) );
  INV_X1 U211 ( .A(P1_P1_InstAddrPointer_PTR26), .ZN(_02745__PTR26) );
  INV_X1 U212 ( .A(P1_P1_InstAddrPointer_PTR27), .ZN(_02745__PTR27) );
  INV_X1 U213 ( .A(P1_P1_InstAddrPointer_PTR28), .ZN(_02745__PTR28) );
  INV_X1 U214 ( .A(P1_P1_InstAddrPointer_PTR29), .ZN(_02745__PTR29) );
  INV_X1 U215 ( .A(P1_P1_InstAddrPointer_PTR30), .ZN(_02745__PTR30) );
  INV_X1 U216 ( .A(P1_P1_InstAddrPointer_PTR8), .ZN(_02745__PTR8) );
  INV_X1 U217 ( .A(P1_P1_InstAddrPointer_PTR9), .ZN(_02745__PTR9) );
  INV_X1 U218 ( .A(P1_P1_InstAddrPointer_PTR10), .ZN(_02745__PTR10) );
  INV_X1 U219 ( .A(P1_P1_InstAddrPointer_PTR11), .ZN(_02745__PTR11) );
  INV_X1 U220 ( .A(P1_P1_InstAddrPointer_PTR12), .ZN(_02745__PTR12) );
  INV_X1 U221 ( .A(P1_P1_InstAddrPointer_PTR13), .ZN(_02745__PTR13) );
  INV_X1 U222 ( .A(P1_P1_InstAddrPointer_PTR14), .ZN(_02745__PTR14) );
  INV_X1 U223 ( .A(P1_P1_InstAddrPointer_PTR15), .ZN(_02745__PTR15) );
  INV_X1 U224 ( .A(P1_P1_InstAddrPointer_PTR4), .ZN(_02745__PTR4) );
  INV_X1 U225 ( .A(P1_P1_InstAddrPointer_PTR5), .ZN(_02745__PTR5) );
  INV_X1 U226 ( .A(P1_P1_InstAddrPointer_PTR6), .ZN(_02745__PTR6) );
  INV_X1 U227 ( .A(P1_P1_InstAddrPointer_PTR7), .ZN(_02745__PTR7) );
  INV_X1 U228 ( .A(P1_P1_InstAddrPointer_PTR3), .ZN(_02745__PTR3) );
  INV_X1 U229 ( .A(_02746__PTR4), .ZN(_02749__PTR4) );
  INV_X1 U230 ( .A(_02720__PTR5), .ZN(_02716__PTR5) );
  INV_X1 U231 ( .A(_02739__PTR4), .ZN(_02742__PTR4) );
  INV_X1 U232 ( .A(_02718__PTR0), .ZN(_02717__PTR0) );
  INV_X1 U233 ( .A(P1_EBX_PTR16), .ZN(_02734__PTR16) );
  INV_X1 U234 ( .A(P1_EBX_PTR17), .ZN(_02734__PTR17) );
  INV_X1 U235 ( .A(P1_EBX_PTR18), .ZN(_02734__PTR18) );
  INV_X1 U236 ( .A(P1_EBX_PTR19), .ZN(_02734__PTR19) );
  INV_X1 U237 ( .A(P1_EBX_PTR20), .ZN(_02734__PTR20) );
  INV_X1 U238 ( .A(P1_EBX_PTR21), .ZN(_02734__PTR21) );
  INV_X1 U239 ( .A(P1_EBX_PTR22), .ZN(_02734__PTR22) );
  INV_X1 U240 ( .A(P1_EBX_PTR23), .ZN(_02734__PTR23) );
  INV_X1 U241 ( .A(P1_EBX_PTR24), .ZN(_02734__PTR24) );
  INV_X1 U242 ( .A(P1_EBX_PTR25), .ZN(_02734__PTR25) );
  INV_X1 U243 ( .A(P1_EBX_PTR26), .ZN(_02734__PTR26) );
  INV_X1 U244 ( .A(P1_EBX_PTR27), .ZN(_02734__PTR27) );
  INV_X1 U245 ( .A(P1_EBX_PTR28), .ZN(_02734__PTR28) );
  INV_X1 U246 ( .A(P1_EBX_PTR29), .ZN(_02734__PTR29) );
  INV_X1 U247 ( .A(P1_EBX_PTR30), .ZN(_02734__PTR30) );
  INV_X1 U248 ( .A(P1_EBX_PTR8), .ZN(_02734__PTR8) );
  INV_X1 U249 ( .A(P1_EBX_PTR9), .ZN(_02734__PTR9) );
  INV_X1 U250 ( .A(P1_EBX_PTR10), .ZN(_02734__PTR10) );
  INV_X1 U251 ( .A(P1_EBX_PTR11), .ZN(_02734__PTR11) );
  INV_X1 U252 ( .A(P1_EBX_PTR12), .ZN(_02734__PTR12) );
  INV_X1 U253 ( .A(P1_EBX_PTR13), .ZN(_02734__PTR13) );
  INV_X1 U254 ( .A(P1_EBX_PTR14), .ZN(_02734__PTR14) );
  INV_X1 U255 ( .A(P1_EBX_PTR15), .ZN(_02734__PTR15) );
  INV_X1 U256 ( .A(P1_EBX_PTR4), .ZN(_02734__PTR4) );
  INV_X1 U257 ( .A(P1_EBX_PTR5), .ZN(_02734__PTR5) );
  INV_X1 U258 ( .A(P1_EBX_PTR6), .ZN(_02734__PTR6) );
  INV_X1 U259 ( .A(P1_EBX_PTR7), .ZN(_02734__PTR7) );
  INV_X1 U260 ( .A(P1_EBX_PTR2), .ZN(_02734__PTR2) );
  INV_X1 U261 ( .A(P1_EBX_PTR3), .ZN(_02734__PTR3) );
  INV_X1 U262 ( .A(P1_EBX_PTR1), .ZN(_02734__PTR1) );
  INV_X1 U263 ( .A(P1_EBX_PTR0), .ZN(_02100__PTR32) );
  INV_X1 U264 ( .A(P1_P1_InstAddrPointer_PTR2), .ZN(_02745__PTR2) );
  INV_X1 U265 ( .A(P1_P1_InstAddrPointer_PTR1), .ZN(_02084__PTR33) );
  INV_X1 U266 ( .A(P1_P1_InstAddrPointer_PTR0), .ZN(_02084__PTR0) );
  INV_X1 U267 ( .A(_02809__PTR0), .ZN(_02939__PTR0) );
  INV_X1 U268 ( .A(_02464__PTR1), .ZN(_00277_) );
  INV_X1 U269 ( .A(_02464__PTR2), .ZN(_00278_) );
  INV_X1 U270 ( .A(_02464__PTR5), .ZN(_00279_) );
  INV_X1 U271 ( .A(_02464__PTR6), .ZN(_00280_) );
  INV_X1 U272 ( .A(_02464__PTR4), .ZN(_00281_) );
  INV_X1 U273 ( .A(_02464__PTR7), .ZN(_00282_) );
  INV_X1 U274 ( .A(_02464__PTR0), .ZN(_00283_) );
  INV_X1 U275 ( .A(_02464__PTR3), .ZN(_00284_) );
  INV_X1 U276 ( .A(_01892__PTR144), .ZN(_02715__PTR16) );
  INV_X1 U277 ( .A(_01892__PTR145), .ZN(_02715__PTR17) );
  INV_X1 U278 ( .A(_01892__PTR146), .ZN(_02715__PTR18) );
  INV_X1 U279 ( .A(_01892__PTR147), .ZN(_02715__PTR19) );
  INV_X1 U280 ( .A(_01892__PTR148), .ZN(_02715__PTR20) );
  INV_X1 U281 ( .A(_01892__PTR149), .ZN(_02715__PTR21) );
  INV_X1 U282 ( .A(_01892__PTR150), .ZN(_02715__PTR22) );
  INV_X1 U283 ( .A(_01892__PTR151), .ZN(_02715__PTR23) );
  INV_X1 U284 ( .A(_01892__PTR152), .ZN(_02715__PTR24) );
  INV_X1 U285 ( .A(_01892__PTR153), .ZN(_02715__PTR25) );
  INV_X1 U286 ( .A(_01892__PTR154), .ZN(_02715__PTR26) );
  INV_X1 U287 ( .A(_01892__PTR155), .ZN(_02715__PTR27) );
  INV_X1 U288 ( .A(_01892__PTR156), .ZN(_02715__PTR28) );
  INV_X1 U289 ( .A(_01892__PTR157), .ZN(_02715__PTR29) );
  INV_X1 U290 ( .A(_01892__PTR158), .ZN(_02715__PTR30) );
  INV_X1 U291 ( .A(_01892__PTR136), .ZN(_02715__PTR8) );
  INV_X1 U292 ( .A(_01892__PTR137), .ZN(_02715__PTR9) );
  INV_X1 U293 ( .A(_01892__PTR138), .ZN(_02715__PTR10) );
  INV_X1 U294 ( .A(_01892__PTR139), .ZN(_02715__PTR11) );
  INV_X1 U295 ( .A(_01892__PTR140), .ZN(_02715__PTR12) );
  INV_X1 U296 ( .A(_01892__PTR141), .ZN(_02715__PTR13) );
  INV_X1 U297 ( .A(_01892__PTR142), .ZN(_02715__PTR14) );
  INV_X1 U298 ( .A(_01892__PTR143), .ZN(_02715__PTR15) );
  INV_X1 U299 ( .A(_01892__PTR132), .ZN(_02715__PTR4) );
  INV_X1 U300 ( .A(_01892__PTR133), .ZN(_02715__PTR5) );
  INV_X1 U301 ( .A(_01892__PTR134), .ZN(_02715__PTR6) );
  INV_X1 U302 ( .A(_01892__PTR135), .ZN(_02715__PTR7) );
  INV_X1 U303 ( .A(_01892__PTR130), .ZN(_02715__PTR2) );
  INV_X1 U304 ( .A(_01892__PTR131), .ZN(_02715__PTR3) );
  INV_X1 U305 ( .A(P1_P1_PhyAddrPointer_PTR0), .ZN(_02715__PTR0) );
  INV_X1 U306 ( .A(P1_P1_InstQueueWr_Addr_PTR0), .ZN(_01836__PTR0) );
  INV_X1 U307 ( .A(P2_P1_InstAddrPointer_PTR16), .ZN(_02990__PTR16) );
  INV_X1 U308 ( .A(P2_P1_InstAddrPointer_PTR19), .ZN(_02990__PTR19) );
  INV_X1 U309 ( .A(P2_P1_InstAddrPointer_PTR21), .ZN(_02990__PTR21) );
  INV_X1 U310 ( .A(P2_P1_InstAddrPointer_PTR26), .ZN(_02990__PTR26) );
  INV_X1 U311 ( .A(P2_P1_InstAddrPointer_PTR8), .ZN(_02990__PTR8) );
  INV_X1 U312 ( .A(P2_P1_InstAddrPointer_PTR13), .ZN(_02990__PTR13) );
  INV_X1 U313 ( .A(P2_P1_InstAddrPointer_PTR4), .ZN(_02990__PTR4) );
  INV_X1 U314 ( .A(P2_P1_InstAddrPointer_PTR3), .ZN(_02990__PTR3) );
  INV_X1 U315 ( .A(_02991__PTR4), .ZN(_02994__PTR4) );
  INV_X1 U316 ( .A(_02965__PTR5), .ZN(_02961__PTR5) );
  INV_X1 U317 ( .A(P2_P1_InstQueueRd_Addr_PTR2), .ZN(_02178__PTR5) );
  INV_X1 U318 ( .A(_02984__PTR4), .ZN(_02987__PTR4) );
  INV_X1 U319 ( .A(P2_EBX_PTR16), .ZN(_02979__PTR16) );
  INV_X1 U320 ( .A(P2_EBX_PTR17), .ZN(_02979__PTR17) );
  INV_X1 U321 ( .A(P2_EBX_PTR19), .ZN(_02979__PTR19) );
  INV_X1 U322 ( .A(P2_EBX_PTR21), .ZN(_02979__PTR21) );
  INV_X1 U323 ( .A(P2_EBX_PTR25), .ZN(_02979__PTR25) );
  INV_X1 U324 ( .A(P2_EBX_PTR26), .ZN(_02979__PTR26) );
  INV_X1 U325 ( .A(P2_EBX_PTR30), .ZN(_02979__PTR30) );
  INV_X1 U326 ( .A(P2_EBX_PTR8), .ZN(_02979__PTR8) );
  INV_X1 U327 ( .A(P2_EBX_PTR9), .ZN(_02979__PTR9) );
  INV_X1 U328 ( .A(P2_EBX_PTR13), .ZN(_02979__PTR13) );
  INV_X1 U329 ( .A(P2_EBX_PTR15), .ZN(_02979__PTR15) );
  INV_X1 U330 ( .A(P2_EBX_PTR4), .ZN(_02979__PTR4) );
  INV_X1 U331 ( .A(P2_EBX_PTR5), .ZN(_02979__PTR5) );
  INV_X1 U332 ( .A(P2_EBX_PTR6), .ZN(_02979__PTR6) );
  INV_X1 U333 ( .A(P2_EBX_PTR3), .ZN(_02979__PTR3) );
  INV_X1 U334 ( .A(P2_EBX_PTR1), .ZN(_02979__PTR1) );
  INV_X1 U335 ( .A(P2_EBX_PTR0), .ZN(_02389__PTR32) );
  INV_X1 U336 ( .A(P2_P1_InstAddrPointer_PTR0), .ZN(_02373__PTR0) );
  INV_X1 U337 ( .A(P2_P1_InstAddrPointer_PTR2), .ZN(_02990__PTR2) );
  INV_X1 U338 ( .A(P2_P1_InstAddrPointer_PTR1), .ZN(_02373__PTR33) );
  INV_X1 U339 ( .A(_03054__PTR0), .ZN(_03184__PTR0) );
  INV_X1 U340 ( .A(P2_P1_PhyAddrPointer_PTR1), .ZN(_02184__PTR129) );
  INV_X1 U341 ( .A(_02184__PTR145), .ZN(_02960__PTR17) );
  INV_X1 U342 ( .A(_02184__PTR146), .ZN(_02960__PTR18) );
  INV_X1 U343 ( .A(_02184__PTR147), .ZN(_02960__PTR19) );
  INV_X1 U344 ( .A(_02184__PTR148), .ZN(_02960__PTR20) );
  INV_X1 U345 ( .A(_02184__PTR154), .ZN(_02960__PTR26) );
  INV_X1 U346 ( .A(_02184__PTR158), .ZN(_02960__PTR30) );
  INV_X1 U347 ( .A(_02184__PTR138), .ZN(_02960__PTR10) );
  INV_X1 U348 ( .A(_02184__PTR140), .ZN(_02960__PTR12) );
  INV_X1 U349 ( .A(_02184__PTR142), .ZN(_02960__PTR14) );
  INV_X1 U350 ( .A(_02184__PTR134), .ZN(_02960__PTR6) );
  INV_X1 U351 ( .A(_02184__PTR135), .ZN(_02960__PTR7) );
  INV_X1 U352 ( .A(_02184__PTR130), .ZN(_02960__PTR2) );
  INV_X1 U353 ( .A(_02184__PTR131), .ZN(_02960__PTR3) );
  INV_X1 U354 ( .A(P3_P1_InstAddrPointer_PTR17), .ZN(_03235__PTR17) );
  INV_X1 U355 ( .A(P3_P1_InstAddrPointer_PTR20), .ZN(_03235__PTR20) );
  INV_X1 U356 ( .A(P3_P1_InstAddrPointer_PTR21), .ZN(_03235__PTR21) );
  INV_X1 U357 ( .A(P3_P1_InstAddrPointer_PTR22), .ZN(_03235__PTR22) );
  INV_X1 U358 ( .A(P3_P1_InstAddrPointer_PTR28), .ZN(_03235__PTR28) );
  INV_X1 U359 ( .A(P3_P1_InstAddrPointer_PTR10), .ZN(_03235__PTR10) );
  INV_X1 U360 ( .A(P3_P1_InstAddrPointer_PTR11), .ZN(_03235__PTR11) );
  INV_X1 U361 ( .A(P3_P1_InstAddrPointer_PTR4), .ZN(_03235__PTR4) );
  INV_X1 U362 ( .A(P3_P1_InstAddrPointer_PTR7), .ZN(_03235__PTR7) );
  INV_X1 U363 ( .A(_03236__PTR4), .ZN(_03239__PTR4) );
  INV_X1 U364 ( .A(_03210__PTR5), .ZN(_03206__PTR5) );
  INV_X1 U365 ( .A(P3_P1_InstQueueRd_Addr_PTR0), .ZN(_02465__PTR3) );
  INV_X1 U366 ( .A(_03229__PTR4), .ZN(_03232__PTR4) );
  INV_X1 U367 ( .A(P3_EBX_PTR20), .ZN(_03224__PTR20) );
  INV_X1 U368 ( .A(P3_EBX_PTR2), .ZN(_03224__PTR2) );
  INV_X1 U369 ( .A(P3_EBX_PTR3), .ZN(_03224__PTR3) );
  INV_X1 U370 ( .A(P3_P1_InstAddrPointer_PTR0), .ZN(_02662__PTR0) );
  INV_X1 U371 ( .A(P3_P1_InstAddrPointer_PTR1), .ZN(_02662__PTR33) );
  INV_X1 U372 ( .A(_03299__PTR0), .ZN(_03429__PTR0) );
  INV_X1 U373 ( .A(_02473__PTR132), .ZN(_03205__PTR4) );
  INV_X1 U374 ( .A(_02473__PTR133), .ZN(_03205__PTR5) );
  INV_X1 U375 ( .A(_02473__PTR131), .ZN(_03205__PTR3) );
  INV_X1 U376 ( .A(P3_P1_PhyAddrPointer_PTR0), .ZN(_03205__PTR0) );
  INV_X1 U377 ( .A(P1_DataWidth_PTR0), .ZN(_00289_) );
  INV_X1 U378 ( .A(P1_P1_InstQueueRd_Addr_PTR1), .ZN(_01890__PTR4) );
  INV_X1 U379 ( .A(P1_P1_InstQueueRd_Addr_PTR2), .ZN(_01886__PTR5) );
  INV_X1 U380 ( .A(P1_EAX_PTR0), .ZN(_02096__PTR32) );
  INV_X1 U381 ( .A(P1_P1_PhyAddrPointer_PTR2), .ZN(_02795__PTR0) );
  INV_X1 U382 ( .A(P2_DataWidth_PTR0), .ZN(_00290_) );
  INV_X1 U383 ( .A(P2_P1_InstQueueRd_Addr_PTR0), .ZN(_02176__PTR3) );
  INV_X1 U384 ( .A(P2_EAX_PTR0), .ZN(_02385__PTR32) );
  INV_X1 U385 ( .A(P2_rEIP_PTR1), .ZN(_02174__PTR7) );
  INV_X1 U386 ( .A(P2_P1_PhyAddrPointer_PTR2), .ZN(_03040__PTR0) );
  INV_X1 U387 ( .A(P3_DataWidth_PTR0), .ZN(_00291_) );
  INV_X1 U388 ( .A(P3_EBX_PTR0), .ZN(_02678__PTR32) );
  INV_X1 U389 ( .A(P3_P1_InstQueueRd_Addr_PTR1), .ZN(_02471__PTR4) );
  INV_X1 U390 ( .A(P3_P1_InstQueueRd_Addr_PTR2), .ZN(_02467__PTR5) );
  INV_X1 U391 ( .A(P3_EAX_PTR0), .ZN(_02674__PTR32) );
  INV_X1 U392 ( .A(P3_rEIP_PTR1), .ZN(_02463__PTR7) );
  INV_X1 U393 ( .A(P3_P1_PhyAddrPointer_PTR2), .ZN(_03285__PTR0) );
  INV_X1 U394 ( .A(_02963__PTR0), .ZN(_02962__PTR0) );
  INV_X1 U395 ( .A(_03208__PTR0), .ZN(_03207__PTR0) );
  INV_X1 U396 ( .A(_02224__PTR57), .ZN(_02991__PTR1) );
  INV_X1 U397 ( .A(_02224__PTR59), .ZN(_02991__PTR3) );
  INV_X1 U398 ( .A(_02224__PTR58), .ZN(_02991__PTR2) );
  INV_X1 U399 ( .A(_02513__PTR59), .ZN(_03236__PTR3) );
  INV_X1 U400 ( .A(P1_P1_PhyAddrPointer_PTR1), .ZN(_01892__PTR129) );
  INV_X1 U401 ( .A(P3_P1_PhyAddrPointer_PTR1), .ZN(_02473__PTR129) );
  INV_X1 U402 ( .A(P3_P1_State2_PTR2), .ZN(_00299_) );
  INV_X1 U403 ( .A(P3_P1_State2_PTR1), .ZN(_00293_) );
  INV_X1 U404 ( .A(P3_P1_State2_PTR3), .ZN(_00292_) );
  INV_X1 U405 ( .A(P3_P1_State2_PTR0), .ZN(_00298_) );
  INV_X1 U406 ( .A(_02581_), .ZN(_00307_) );
  INV_X1 U407 ( .A(P3_State_PTR1), .ZN(_00288_) );
  INV_X1 U408 ( .A(_02475__PTR28), .ZN(_00308_) );
  INV_X1 U409 ( .A(P2_State_PTR1), .ZN(_00286_) );
  INV_X1 U410 ( .A(_02292_), .ZN(_00309_) );
  INV_X1 U411 ( .A(P2_State_PTR2), .ZN(_00285_) );
  INV_X1 U412 ( .A(P2_P1_State2_PTR2), .ZN(_00301_) );
  INV_X1 U413 ( .A(P2_P1_State2_PTR0), .ZN(_00300_) );
  INV_X1 U414 ( .A(P1_P1_State2_PTR0), .ZN(_00302_) );
  INV_X1 U415 ( .A(P1_P1_State2_PTR2), .ZN(_00303_) );
  INV_X1 U416 ( .A(_02186__PTR28), .ZN(_00304_) );
  INV_X1 U417 ( .A(_02001_), .ZN(_00312_) );
  INV_X1 U418 ( .A(P1_State_PTR1), .ZN(_00276_) );
  INV_X1 U419 ( .A(_01894__PTR28), .ZN(_00310_) );
  INV_X1 U420 ( .A(P3_State_PTR2), .ZN(_00287_) );
  INV_X1 U421 ( .A(P1_State_PTR2), .ZN(_00275_) );
  OR2_X1 U422 ( .A1(_02115__PTR23), .A2(_02115__PTR55), .ZN(_01743_) );
  OR2_X1 U423 ( .A1(_01743_), .A2(_02115__PTR87), .ZN(_02117__PTR23) );
  OR2_X1 U424 ( .A1(_02115__PTR22), .A2(_02115__PTR54), .ZN(_00313_) );
  OR2_X1 U425 ( .A1(_00313_), .A2(_02115__PTR86), .ZN(_02117__PTR22) );
  OR2_X1 U426 ( .A1(_02115__PTR21), .A2(_02115__PTR53), .ZN(_00314_) );
  OR2_X1 U427 ( .A1(_00314_), .A2(_02115__PTR85), .ZN(_02117__PTR21) );
  OR2_X1 U428 ( .A1(_02115__PTR20), .A2(_02115__PTR52), .ZN(_00315_) );
  OR2_X1 U429 ( .A1(_00315_), .A2(_02115__PTR84), .ZN(_02117__PTR20) );
  OR2_X1 U430 ( .A1(_02115__PTR19), .A2(_02115__PTR51), .ZN(_00316_) );
  OR2_X1 U431 ( .A1(_00316_), .A2(_02115__PTR83), .ZN(_02117__PTR19) );
  OR2_X1 U432 ( .A1(_02115__PTR18), .A2(_02115__PTR50), .ZN(_00317_) );
  OR2_X1 U433 ( .A1(_00317_), .A2(_02115__PTR82), .ZN(_02117__PTR18) );
  OR2_X1 U434 ( .A1(_02115__PTR17), .A2(_02115__PTR49), .ZN(_00318_) );
  OR2_X1 U435 ( .A1(_00318_), .A2(_02115__PTR81), .ZN(_02117__PTR17) );
  OR2_X1 U436 ( .A1(_02115__PTR16), .A2(_02115__PTR48), .ZN(_00319_) );
  OR2_X1 U437 ( .A1(_00319_), .A2(_02115__PTR80), .ZN(_02117__PTR16) );
  OR2_X1 U438 ( .A1(_02115__PTR15), .A2(_02115__PTR47), .ZN(_00320_) );
  OR2_X1 U439 ( .A1(_00320_), .A2(_02115__PTR79), .ZN(_02117__PTR15) );
  OR2_X1 U440 ( .A1(_02115__PTR14), .A2(_02115__PTR46), .ZN(_00321_) );
  OR2_X1 U441 ( .A1(_00321_), .A2(_02115__PTR78), .ZN(_02117__PTR14) );
  OR2_X1 U442 ( .A1(_02115__PTR13), .A2(_02115__PTR45), .ZN(_00322_) );
  OR2_X1 U443 ( .A1(_00322_), .A2(_02115__PTR77), .ZN(_02117__PTR13) );
  OR2_X1 U444 ( .A1(_02115__PTR12), .A2(_02115__PTR44), .ZN(_00323_) );
  OR2_X1 U445 ( .A1(_00323_), .A2(_02115__PTR76), .ZN(_02117__PTR12) );
  OR2_X1 U446 ( .A1(_02115__PTR11), .A2(_02115__PTR43), .ZN(_00324_) );
  OR2_X1 U447 ( .A1(_00324_), .A2(_02115__PTR75), .ZN(_02117__PTR11) );
  OR2_X1 U448 ( .A1(_02115__PTR10), .A2(_02115__PTR42), .ZN(_00325_) );
  OR2_X1 U449 ( .A1(_00325_), .A2(_02115__PTR74), .ZN(_02117__PTR10) );
  OR2_X1 U450 ( .A1(_02115__PTR9), .A2(_02115__PTR41), .ZN(_00326_) );
  OR2_X1 U451 ( .A1(_00326_), .A2(_02115__PTR73), .ZN(_02117__PTR9) );
  OR2_X1 U452 ( .A1(_02115__PTR8), .A2(_02115__PTR40), .ZN(_00327_) );
  OR2_X1 U453 ( .A1(_00327_), .A2(_02115__PTR72), .ZN(_02117__PTR8) );
  OR2_X1 U454 ( .A1(_02115__PTR7), .A2(_02115__PTR39), .ZN(_00328_) );
  OR2_X1 U455 ( .A1(_00328_), .A2(_02115__PTR71), .ZN(_02117__PTR7) );
  OR2_X1 U456 ( .A1(_02115__PTR6), .A2(_02115__PTR38), .ZN(_00329_) );
  OR2_X1 U457 ( .A1(_00329_), .A2(_02115__PTR70), .ZN(_02117__PTR6) );
  OR2_X1 U458 ( .A1(_02115__PTR5), .A2(_02115__PTR37), .ZN(_00330_) );
  OR2_X1 U459 ( .A1(_00330_), .A2(_02115__PTR69), .ZN(_02117__PTR5) );
  OR2_X1 U460 ( .A1(_02115__PTR4), .A2(_02115__PTR36), .ZN(_00331_) );
  OR2_X1 U461 ( .A1(_00331_), .A2(_02115__PTR68), .ZN(_02117__PTR4) );
  OR2_X1 U462 ( .A1(_02115__PTR3), .A2(_02115__PTR35), .ZN(_00332_) );
  OR2_X1 U463 ( .A1(_00332_), .A2(_02115__PTR67), .ZN(_02117__PTR3) );
  OR2_X1 U464 ( .A1(_02115__PTR2), .A2(_02115__PTR34), .ZN(_00333_) );
  OR2_X1 U465 ( .A1(_00333_), .A2(_02115__PTR66), .ZN(_02117__PTR2) );
  OR2_X1 U466 ( .A1(_02115__PTR1), .A2(_02115__PTR33), .ZN(_00334_) );
  OR2_X1 U467 ( .A1(_00334_), .A2(_02115__PTR65), .ZN(_02117__PTR1) );
  OR2_X1 U468 ( .A1(_02115__PTR0), .A2(_02115__PTR32), .ZN(_00335_) );
  OR2_X1 U469 ( .A1(_00335_), .A2(_02115__PTR64), .ZN(_02117__PTR0) );
  OR2_X1 U470 ( .A1(_02116__PTR0), .A2(_01863__PTR0), .ZN(_00336_) );
  OR2_X1 U471 ( .A1(_00336_), .A2(_01863__PTR2), .ZN(_02927_) );
  OR2_X1 U472 ( .A1(_02112__PTR15), .A2(_02112__PTR31), .ZN(_00337_) );
  OR2_X1 U473 ( .A1(_00337_), .A2(_02112__PTR47), .ZN(_02113__PTR15) );
  OR2_X1 U474 ( .A1(_02112__PTR14), .A2(_02112__PTR30), .ZN(_00338_) );
  OR2_X1 U475 ( .A1(_00338_), .A2(_02112__PTR46), .ZN(_02113__PTR14) );
  OR2_X1 U476 ( .A1(_02112__PTR13), .A2(_02112__PTR29), .ZN(_00339_) );
  OR2_X1 U477 ( .A1(_00339_), .A2(_02112__PTR45), .ZN(_02113__PTR13) );
  OR2_X1 U478 ( .A1(_02112__PTR12), .A2(_02112__PTR28), .ZN(_00340_) );
  OR2_X1 U479 ( .A1(_00340_), .A2(_02112__PTR44), .ZN(_02113__PTR12) );
  OR2_X1 U480 ( .A1(_02112__PTR11), .A2(_02112__PTR27), .ZN(_00341_) );
  OR2_X1 U481 ( .A1(_00341_), .A2(_02112__PTR43), .ZN(_02113__PTR11) );
  OR2_X1 U482 ( .A1(_02112__PTR10), .A2(_02112__PTR26), .ZN(_00342_) );
  OR2_X1 U483 ( .A1(_00342_), .A2(_02112__PTR42), .ZN(_02113__PTR10) );
  OR2_X1 U484 ( .A1(_02112__PTR9), .A2(_02112__PTR25), .ZN(_00343_) );
  OR2_X1 U485 ( .A1(_00343_), .A2(_02112__PTR41), .ZN(_02113__PTR9) );
  OR2_X1 U486 ( .A1(_02112__PTR8), .A2(_02112__PTR24), .ZN(_00344_) );
  OR2_X1 U487 ( .A1(_00344_), .A2(_02112__PTR40), .ZN(_02113__PTR8) );
  OR2_X1 U488 ( .A1(_02112__PTR7), .A2(_02112__PTR23), .ZN(_00345_) );
  OR2_X1 U489 ( .A1(_00345_), .A2(_02112__PTR39), .ZN(_02113__PTR7) );
  OR2_X1 U490 ( .A1(_02112__PTR6), .A2(_02112__PTR22), .ZN(_00346_) );
  OR2_X1 U491 ( .A1(_00346_), .A2(_02112__PTR38), .ZN(_02113__PTR6) );
  OR2_X1 U492 ( .A1(_02112__PTR5), .A2(_02112__PTR21), .ZN(_00347_) );
  OR2_X1 U493 ( .A1(_00347_), .A2(_02112__PTR37), .ZN(_02113__PTR5) );
  OR2_X1 U494 ( .A1(_02112__PTR4), .A2(_02112__PTR20), .ZN(_00348_) );
  OR2_X1 U495 ( .A1(_00348_), .A2(_02112__PTR36), .ZN(_02113__PTR4) );
  OR2_X1 U496 ( .A1(_02112__PTR3), .A2(_02112__PTR19), .ZN(_00349_) );
  OR2_X1 U497 ( .A1(_00349_), .A2(_02112__PTR35), .ZN(_02113__PTR3) );
  OR2_X1 U498 ( .A1(_02112__PTR2), .A2(_02112__PTR18), .ZN(_00350_) );
  OR2_X1 U499 ( .A1(_00350_), .A2(_02112__PTR34), .ZN(_02113__PTR2) );
  OR2_X1 U500 ( .A1(_02112__PTR1), .A2(_02112__PTR17), .ZN(_00351_) );
  OR2_X1 U501 ( .A1(_00351_), .A2(_02112__PTR33), .ZN(_02113__PTR1) );
  OR2_X1 U502 ( .A1(_02112__PTR0), .A2(_02112__PTR16), .ZN(_00352_) );
  OR2_X1 U503 ( .A1(_00352_), .A2(_02112__PTR32), .ZN(_02113__PTR0) );
  OR2_X1 U504 ( .A1(_02108__PTR14), .A2(_02108__PTR29), .ZN(_00354_) );
  OR2_X1 U505 ( .A1(_00354_), .A2(_02108__PTR44), .ZN(_02110__PTR14) );
  OR2_X1 U506 ( .A1(_02108__PTR13), .A2(_02108__PTR28), .ZN(_00355_) );
  OR2_X1 U507 ( .A1(_00355_), .A2(_02108__PTR43), .ZN(_02110__PTR13) );
  OR2_X1 U508 ( .A1(_02108__PTR12), .A2(_02108__PTR27), .ZN(_00356_) );
  OR2_X1 U509 ( .A1(_00356_), .A2(_02108__PTR42), .ZN(_02110__PTR12) );
  OR2_X1 U510 ( .A1(_02108__PTR11), .A2(_02108__PTR26), .ZN(_00357_) );
  OR2_X1 U511 ( .A1(_00357_), .A2(_02108__PTR41), .ZN(_02110__PTR11) );
  OR2_X1 U512 ( .A1(_02108__PTR10), .A2(_02108__PTR25), .ZN(_00358_) );
  OR2_X1 U513 ( .A1(_00358_), .A2(_02108__PTR40), .ZN(_02110__PTR10) );
  OR2_X1 U514 ( .A1(_02108__PTR9), .A2(_02108__PTR24), .ZN(_00359_) );
  OR2_X1 U515 ( .A1(_00359_), .A2(_02108__PTR39), .ZN(_02110__PTR9) );
  OR2_X1 U516 ( .A1(_02108__PTR8), .A2(_02108__PTR23), .ZN(_00360_) );
  OR2_X1 U517 ( .A1(_00360_), .A2(_02108__PTR38), .ZN(_02110__PTR8) );
  OR2_X1 U518 ( .A1(_02108__PTR7), .A2(_02108__PTR22), .ZN(_00361_) );
  OR2_X1 U519 ( .A1(_00361_), .A2(_02108__PTR37), .ZN(_02110__PTR7) );
  OR2_X1 U520 ( .A1(_02108__PTR6), .A2(_02108__PTR21), .ZN(_00362_) );
  OR2_X1 U521 ( .A1(_00362_), .A2(_02108__PTR36), .ZN(_02110__PTR6) );
  OR2_X1 U522 ( .A1(_02108__PTR5), .A2(_02108__PTR20), .ZN(_00363_) );
  OR2_X1 U523 ( .A1(_00363_), .A2(_02108__PTR35), .ZN(_02110__PTR5) );
  OR2_X1 U524 ( .A1(_02108__PTR4), .A2(_02108__PTR19), .ZN(_00364_) );
  OR2_X1 U525 ( .A1(_00364_), .A2(_02108__PTR34), .ZN(_02110__PTR4) );
  OR2_X1 U526 ( .A1(_02108__PTR3), .A2(_02108__PTR18), .ZN(_00365_) );
  OR2_X1 U527 ( .A1(_00365_), .A2(_02108__PTR33), .ZN(_02110__PTR3) );
  OR2_X1 U528 ( .A1(_02108__PTR2), .A2(_02108__PTR17), .ZN(_00366_) );
  OR2_X1 U529 ( .A1(_00366_), .A2(_02108__PTR32), .ZN(_02110__PTR2) );
  OR2_X1 U530 ( .A1(_02108__PTR1), .A2(_02108__PTR16), .ZN(_00367_) );
  OR2_X1 U531 ( .A1(_00367_), .A2(_02108__PTR31), .ZN(_02110__PTR1) );
  OR2_X1 U532 ( .A1(_02108__PTR0), .A2(_02108__PTR15), .ZN(_00368_) );
  OR2_X1 U533 ( .A1(_00368_), .A2(_02108__PTR30), .ZN(_02110__PTR0) );
  OR2_X1 U534 ( .A1(_02109__PTR0), .A2(_01863__PTR2), .ZN(_00353_) );
  OR2_X1 U535 ( .A1(_00353_), .A2(_02090__PTR4), .ZN(_02926_) );
  OR2_X1 U536 ( .A1(_02101__PTR0), .A2(_02101__PTR32), .ZN(_00369_) );
  OR2_X1 U537 ( .A1(_00369_), .A2(_02101__PTR64), .ZN(_02103__PTR0) );
  OR2_X1 U538 ( .A1(_02101__PTR1), .A2(_02101__PTR33), .ZN(_00370_) );
  OR2_X1 U539 ( .A1(_00370_), .A2(_02101__PTR65), .ZN(_02103__PTR1) );
  OR2_X1 U540 ( .A1(_02101__PTR2), .A2(_02101__PTR34), .ZN(_00371_) );
  OR2_X1 U541 ( .A1(_00371_), .A2(_02101__PTR66), .ZN(_02103__PTR2) );
  OR2_X1 U542 ( .A1(_02101__PTR3), .A2(_02101__PTR35), .ZN(_00372_) );
  OR2_X1 U543 ( .A1(_00372_), .A2(_02101__PTR67), .ZN(_02103__PTR3) );
  OR2_X1 U544 ( .A1(_02101__PTR4), .A2(_02101__PTR36), .ZN(_00373_) );
  OR2_X1 U545 ( .A1(_00373_), .A2(_02101__PTR68), .ZN(_02103__PTR4) );
  OR2_X1 U546 ( .A1(_02101__PTR5), .A2(_02101__PTR37), .ZN(_00374_) );
  OR2_X1 U547 ( .A1(_00374_), .A2(_02101__PTR69), .ZN(_02103__PTR5) );
  OR2_X1 U548 ( .A1(_02101__PTR6), .A2(_02101__PTR38), .ZN(_00375_) );
  OR2_X1 U549 ( .A1(_00375_), .A2(_02101__PTR70), .ZN(_02103__PTR6) );
  OR2_X1 U550 ( .A1(_02101__PTR7), .A2(_02101__PTR39), .ZN(_00376_) );
  OR2_X1 U551 ( .A1(_00376_), .A2(_02101__PTR71), .ZN(_02103__PTR7) );
  OR2_X1 U552 ( .A1(_02101__PTR8), .A2(_02101__PTR40), .ZN(_00377_) );
  OR2_X1 U553 ( .A1(_00377_), .A2(_02101__PTR72), .ZN(_02103__PTR8) );
  OR2_X1 U554 ( .A1(_02101__PTR9), .A2(_02101__PTR41), .ZN(_00378_) );
  OR2_X1 U555 ( .A1(_00378_), .A2(_02101__PTR73), .ZN(_02103__PTR9) );
  OR2_X1 U556 ( .A1(_02101__PTR10), .A2(_02101__PTR42), .ZN(_00379_) );
  OR2_X1 U557 ( .A1(_00379_), .A2(_02101__PTR74), .ZN(_02103__PTR10) );
  OR2_X1 U558 ( .A1(_02101__PTR11), .A2(_02101__PTR43), .ZN(_00380_) );
  OR2_X1 U559 ( .A1(_00380_), .A2(_02101__PTR75), .ZN(_02103__PTR11) );
  OR2_X1 U560 ( .A1(_02101__PTR12), .A2(_02101__PTR44), .ZN(_00381_) );
  OR2_X1 U561 ( .A1(_00381_), .A2(_02101__PTR76), .ZN(_02103__PTR12) );
  OR2_X1 U562 ( .A1(_02101__PTR13), .A2(_02101__PTR45), .ZN(_00382_) );
  OR2_X1 U563 ( .A1(_00382_), .A2(_02101__PTR77), .ZN(_02103__PTR13) );
  OR2_X1 U564 ( .A1(_02101__PTR14), .A2(_02101__PTR46), .ZN(_00383_) );
  OR2_X1 U565 ( .A1(_00383_), .A2(_02101__PTR78), .ZN(_02103__PTR14) );
  OR2_X1 U566 ( .A1(_02101__PTR15), .A2(_02101__PTR47), .ZN(_00384_) );
  OR2_X1 U567 ( .A1(_00384_), .A2(_02101__PTR79), .ZN(_02103__PTR15) );
  OR2_X1 U568 ( .A1(_02101__PTR16), .A2(_02101__PTR48), .ZN(_00385_) );
  OR2_X1 U569 ( .A1(_00385_), .A2(_02101__PTR80), .ZN(_02103__PTR16) );
  OR2_X1 U570 ( .A1(_02101__PTR17), .A2(_02101__PTR49), .ZN(_00386_) );
  OR2_X1 U571 ( .A1(_00386_), .A2(_02101__PTR81), .ZN(_02103__PTR17) );
  OR2_X1 U572 ( .A1(_02101__PTR18), .A2(_02101__PTR50), .ZN(_00387_) );
  OR2_X1 U573 ( .A1(_00387_), .A2(_02101__PTR82), .ZN(_02103__PTR18) );
  OR2_X1 U574 ( .A1(_02101__PTR19), .A2(_02101__PTR51), .ZN(_00388_) );
  OR2_X1 U575 ( .A1(_00388_), .A2(_02101__PTR83), .ZN(_02103__PTR19) );
  OR2_X1 U576 ( .A1(_02101__PTR20), .A2(_02101__PTR52), .ZN(_00389_) );
  OR2_X1 U577 ( .A1(_00389_), .A2(_02101__PTR84), .ZN(_02103__PTR20) );
  OR2_X1 U578 ( .A1(_02101__PTR21), .A2(_02101__PTR53), .ZN(_00390_) );
  OR2_X1 U579 ( .A1(_00390_), .A2(_02101__PTR85), .ZN(_02103__PTR21) );
  OR2_X1 U580 ( .A1(_02101__PTR22), .A2(_02101__PTR54), .ZN(_00391_) );
  OR2_X1 U581 ( .A1(_00391_), .A2(_02101__PTR86), .ZN(_02103__PTR22) );
  OR2_X1 U582 ( .A1(_02101__PTR23), .A2(_02101__PTR55), .ZN(_00392_) );
  OR2_X1 U583 ( .A1(_00392_), .A2(_02101__PTR87), .ZN(_02103__PTR23) );
  OR2_X1 U584 ( .A1(_02101__PTR24), .A2(_02101__PTR56), .ZN(_00393_) );
  OR2_X1 U585 ( .A1(_00393_), .A2(_02101__PTR88), .ZN(_02103__PTR24) );
  OR2_X1 U586 ( .A1(_02101__PTR25), .A2(_02101__PTR57), .ZN(_00394_) );
  OR2_X1 U587 ( .A1(_00394_), .A2(_02101__PTR89), .ZN(_02103__PTR25) );
  OR2_X1 U588 ( .A1(_02101__PTR26), .A2(_02101__PTR58), .ZN(_00395_) );
  OR2_X1 U589 ( .A1(_00395_), .A2(_02101__PTR90), .ZN(_02103__PTR26) );
  OR2_X1 U590 ( .A1(_02101__PTR27), .A2(_02101__PTR59), .ZN(_00396_) );
  OR2_X1 U591 ( .A1(_00396_), .A2(_02101__PTR91), .ZN(_02103__PTR27) );
  OR2_X1 U592 ( .A1(_02101__PTR28), .A2(_02101__PTR60), .ZN(_00397_) );
  OR2_X1 U593 ( .A1(_00397_), .A2(_02101__PTR92), .ZN(_02103__PTR28) );
  OR2_X1 U594 ( .A1(_02101__PTR29), .A2(_02101__PTR61), .ZN(_00398_) );
  OR2_X1 U595 ( .A1(_00398_), .A2(_02101__PTR93), .ZN(_02103__PTR29) );
  OR2_X1 U596 ( .A1(_02101__PTR30), .A2(_02101__PTR62), .ZN(_00399_) );
  OR2_X1 U597 ( .A1(_00399_), .A2(_02101__PTR94), .ZN(_02103__PTR30) );
  OR2_X1 U598 ( .A1(_02101__PTR31), .A2(_02101__PTR63), .ZN(_00400_) );
  OR2_X1 U599 ( .A1(_00400_), .A2(_02101__PTR95), .ZN(_02103__PTR31) );
  OR2_X1 U600 ( .A1(_02102__PTR0), .A2(_02102__PTR1), .ZN(_00401_) );
  OR2_X1 U601 ( .A1(_00401_), .A2(_02102__PTR2), .ZN(_02924_) );
  OR2_X1 U602 ( .A1(_02097__PTR31), .A2(_02097__PTR63), .ZN(_00402__PTR0) );
  OR2_X1 U603 ( .A1(_02097__PTR95), .A2(_02097__PTR127), .ZN(_00402__PTR1) );
  OR2_X1 U604 ( .A1(_00402__PTR0), .A2(_00402__PTR1), .ZN(_00403_) );
  OR2_X1 U605 ( .A1(_00403_), .A2(_02097__PTR159), .ZN(_02099__PTR31) );
  OR2_X1 U606 ( .A1(_02097__PTR30), .A2(_02097__PTR62), .ZN(_00404__PTR0) );
  OR2_X1 U607 ( .A1(_02097__PTR94), .A2(_02097__PTR126), .ZN(_00404__PTR1) );
  OR2_X1 U608 ( .A1(_00404__PTR0), .A2(_00404__PTR1), .ZN(_00405_) );
  OR2_X1 U609 ( .A1(_00405_), .A2(_02097__PTR158), .ZN(_02099__PTR30) );
  OR2_X1 U610 ( .A1(_02097__PTR29), .A2(_02097__PTR61), .ZN(_00406__PTR0) );
  OR2_X1 U611 ( .A1(_02097__PTR93), .A2(_02097__PTR125), .ZN(_00406__PTR1) );
  OR2_X1 U612 ( .A1(_00406__PTR0), .A2(_00406__PTR1), .ZN(_00407_) );
  OR2_X1 U613 ( .A1(_00407_), .A2(_02097__PTR157), .ZN(_02099__PTR29) );
  OR2_X1 U614 ( .A1(_02097__PTR28), .A2(_02097__PTR60), .ZN(_00408__PTR0) );
  OR2_X1 U615 ( .A1(_02097__PTR92), .A2(_02097__PTR124), .ZN(_00408__PTR1) );
  OR2_X1 U616 ( .A1(_00408__PTR0), .A2(_00408__PTR1), .ZN(_00409_) );
  OR2_X1 U617 ( .A1(_00409_), .A2(_02097__PTR156), .ZN(_02099__PTR28) );
  OR2_X1 U618 ( .A1(_02097__PTR27), .A2(_02097__PTR59), .ZN(_00410__PTR0) );
  OR2_X1 U619 ( .A1(_02097__PTR91), .A2(_02097__PTR123), .ZN(_00410__PTR1) );
  OR2_X1 U620 ( .A1(_00410__PTR0), .A2(_00410__PTR1), .ZN(_00411_) );
  OR2_X1 U621 ( .A1(_00411_), .A2(_02097__PTR155), .ZN(_02099__PTR27) );
  OR2_X1 U622 ( .A1(_02097__PTR26), .A2(_02097__PTR58), .ZN(_00412__PTR0) );
  OR2_X1 U623 ( .A1(_02097__PTR90), .A2(_02097__PTR122), .ZN(_00412__PTR1) );
  OR2_X1 U624 ( .A1(_00412__PTR0), .A2(_00412__PTR1), .ZN(_00413_) );
  OR2_X1 U625 ( .A1(_00413_), .A2(_02097__PTR154), .ZN(_02099__PTR26) );
  OR2_X1 U626 ( .A1(_02097__PTR25), .A2(_02097__PTR57), .ZN(_00414__PTR0) );
  OR2_X1 U627 ( .A1(_02097__PTR89), .A2(_02097__PTR121), .ZN(_00414__PTR1) );
  OR2_X1 U628 ( .A1(_00414__PTR0), .A2(_00414__PTR1), .ZN(_00415_) );
  OR2_X1 U629 ( .A1(_00415_), .A2(_02097__PTR153), .ZN(_02099__PTR25) );
  OR2_X1 U630 ( .A1(_02097__PTR24), .A2(_02097__PTR56), .ZN(_00416__PTR0) );
  OR2_X1 U631 ( .A1(_02097__PTR88), .A2(_02097__PTR120), .ZN(_00416__PTR1) );
  OR2_X1 U632 ( .A1(_00416__PTR0), .A2(_00416__PTR1), .ZN(_00417_) );
  OR2_X1 U633 ( .A1(_00417_), .A2(_02097__PTR152), .ZN(_02099__PTR24) );
  OR2_X1 U634 ( .A1(_02097__PTR23), .A2(_02097__PTR55), .ZN(_00418__PTR0) );
  OR2_X1 U635 ( .A1(_02097__PTR87), .A2(_02097__PTR119), .ZN(_00418__PTR1) );
  OR2_X1 U636 ( .A1(_00418__PTR0), .A2(_00418__PTR1), .ZN(_00419_) );
  OR2_X1 U637 ( .A1(_00419_), .A2(_02097__PTR151), .ZN(_02099__PTR23) );
  OR2_X1 U638 ( .A1(_02097__PTR22), .A2(_02097__PTR54), .ZN(_00420__PTR0) );
  OR2_X1 U639 ( .A1(_02097__PTR86), .A2(_02097__PTR118), .ZN(_00420__PTR1) );
  OR2_X1 U640 ( .A1(_00420__PTR0), .A2(_00420__PTR1), .ZN(_00421_) );
  OR2_X1 U641 ( .A1(_00421_), .A2(_02097__PTR150), .ZN(_02099__PTR22) );
  OR2_X1 U642 ( .A1(_02097__PTR21), .A2(_02097__PTR53), .ZN(_00422__PTR0) );
  OR2_X1 U643 ( .A1(_02097__PTR85), .A2(_02097__PTR117), .ZN(_00422__PTR1) );
  OR2_X1 U644 ( .A1(_00422__PTR0), .A2(_00422__PTR1), .ZN(_00423_) );
  OR2_X1 U645 ( .A1(_00423_), .A2(_02097__PTR149), .ZN(_02099__PTR21) );
  OR2_X1 U646 ( .A1(_02097__PTR20), .A2(_02097__PTR52), .ZN(_00424__PTR0) );
  OR2_X1 U647 ( .A1(_02097__PTR84), .A2(_02097__PTR116), .ZN(_00424__PTR1) );
  OR2_X1 U648 ( .A1(_00424__PTR0), .A2(_00424__PTR1), .ZN(_00425_) );
  OR2_X1 U649 ( .A1(_00425_), .A2(_02097__PTR148), .ZN(_02099__PTR20) );
  OR2_X1 U650 ( .A1(_02097__PTR19), .A2(_02097__PTR51), .ZN(_00426__PTR0) );
  OR2_X1 U651 ( .A1(_02097__PTR83), .A2(_02097__PTR115), .ZN(_00426__PTR1) );
  OR2_X1 U652 ( .A1(_00426__PTR0), .A2(_00426__PTR1), .ZN(_00427_) );
  OR2_X1 U653 ( .A1(_00427_), .A2(_02097__PTR147), .ZN(_02099__PTR19) );
  OR2_X1 U654 ( .A1(_02097__PTR18), .A2(_02097__PTR50), .ZN(_00428__PTR0) );
  OR2_X1 U655 ( .A1(_02097__PTR82), .A2(_02097__PTR114), .ZN(_00428__PTR1) );
  OR2_X1 U656 ( .A1(_00428__PTR0), .A2(_00428__PTR1), .ZN(_00429_) );
  OR2_X1 U657 ( .A1(_00429_), .A2(_02097__PTR146), .ZN(_02099__PTR18) );
  OR2_X1 U658 ( .A1(_02097__PTR17), .A2(_02097__PTR49), .ZN(_00430__PTR0) );
  OR2_X1 U659 ( .A1(_02097__PTR81), .A2(_02097__PTR113), .ZN(_00430__PTR1) );
  OR2_X1 U660 ( .A1(_00430__PTR0), .A2(_00430__PTR1), .ZN(_00431_) );
  OR2_X1 U661 ( .A1(_00431_), .A2(_02097__PTR145), .ZN(_02099__PTR17) );
  OR2_X1 U662 ( .A1(_02097__PTR16), .A2(_02097__PTR48), .ZN(_00432__PTR0) );
  OR2_X1 U663 ( .A1(_02097__PTR80), .A2(_02097__PTR112), .ZN(_00432__PTR1) );
  OR2_X1 U664 ( .A1(_00432__PTR0), .A2(_00432__PTR1), .ZN(_00433_) );
  OR2_X1 U665 ( .A1(_00433_), .A2(_02097__PTR144), .ZN(_02099__PTR16) );
  OR2_X1 U666 ( .A1(_02097__PTR15), .A2(_02097__PTR47), .ZN(_00434__PTR0) );
  OR2_X1 U667 ( .A1(_02097__PTR79), .A2(_02097__PTR111), .ZN(_00434__PTR1) );
  OR2_X1 U668 ( .A1(_00434__PTR0), .A2(_00434__PTR1), .ZN(_00435_) );
  OR2_X1 U669 ( .A1(_00435_), .A2(_02097__PTR143), .ZN(_02099__PTR15) );
  OR2_X1 U670 ( .A1(_02097__PTR14), .A2(_02097__PTR46), .ZN(_00436__PTR0) );
  OR2_X1 U671 ( .A1(_02097__PTR78), .A2(_02097__PTR110), .ZN(_00436__PTR1) );
  OR2_X1 U672 ( .A1(_00436__PTR0), .A2(_00436__PTR1), .ZN(_00437_) );
  OR2_X1 U673 ( .A1(_00437_), .A2(_02097__PTR142), .ZN(_02099__PTR14) );
  OR2_X1 U674 ( .A1(_02097__PTR13), .A2(_02097__PTR45), .ZN(_00438__PTR0) );
  OR2_X1 U675 ( .A1(_02097__PTR77), .A2(_02097__PTR109), .ZN(_00438__PTR1) );
  OR2_X1 U676 ( .A1(_00438__PTR0), .A2(_00438__PTR1), .ZN(_00439_) );
  OR2_X1 U677 ( .A1(_00439_), .A2(_02097__PTR141), .ZN(_02099__PTR13) );
  OR2_X1 U678 ( .A1(_02097__PTR12), .A2(_02097__PTR44), .ZN(_00440__PTR0) );
  OR2_X1 U679 ( .A1(_02097__PTR76), .A2(_02097__PTR108), .ZN(_00440__PTR1) );
  OR2_X1 U680 ( .A1(_00440__PTR0), .A2(_00440__PTR1), .ZN(_00441_) );
  OR2_X1 U681 ( .A1(_00441_), .A2(_02097__PTR140), .ZN(_02099__PTR12) );
  OR2_X1 U682 ( .A1(_02097__PTR11), .A2(_02097__PTR43), .ZN(_00442__PTR0) );
  OR2_X1 U683 ( .A1(_02097__PTR75), .A2(_02097__PTR107), .ZN(_00442__PTR1) );
  OR2_X1 U684 ( .A1(_00442__PTR0), .A2(_00442__PTR1), .ZN(_00443_) );
  OR2_X1 U685 ( .A1(_00443_), .A2(_02097__PTR139), .ZN(_02099__PTR11) );
  OR2_X1 U686 ( .A1(_02097__PTR10), .A2(_02097__PTR42), .ZN(_00444__PTR0) );
  OR2_X1 U687 ( .A1(_02097__PTR74), .A2(_02097__PTR106), .ZN(_00444__PTR1) );
  OR2_X1 U688 ( .A1(_00444__PTR0), .A2(_00444__PTR1), .ZN(_00445_) );
  OR2_X1 U689 ( .A1(_00445_), .A2(_02097__PTR138), .ZN(_02099__PTR10) );
  OR2_X1 U690 ( .A1(_02097__PTR9), .A2(_02097__PTR41), .ZN(_00446__PTR0) );
  OR2_X1 U691 ( .A1(_02097__PTR73), .A2(_02097__PTR105), .ZN(_00446__PTR1) );
  OR2_X1 U692 ( .A1(_00446__PTR0), .A2(_00446__PTR1), .ZN(_00447_) );
  OR2_X1 U693 ( .A1(_00447_), .A2(_02097__PTR137), .ZN(_02099__PTR9) );
  OR2_X1 U694 ( .A1(_02097__PTR8), .A2(_02097__PTR40), .ZN(_00448__PTR0) );
  OR2_X1 U695 ( .A1(_02097__PTR72), .A2(_02097__PTR104), .ZN(_00448__PTR1) );
  OR2_X1 U696 ( .A1(_00448__PTR0), .A2(_00448__PTR1), .ZN(_00449_) );
  OR2_X1 U697 ( .A1(_00449_), .A2(_02097__PTR136), .ZN(_02099__PTR8) );
  OR2_X1 U698 ( .A1(_02097__PTR7), .A2(_02097__PTR39), .ZN(_00450__PTR0) );
  OR2_X1 U699 ( .A1(_02097__PTR71), .A2(_02097__PTR103), .ZN(_00450__PTR1) );
  OR2_X1 U700 ( .A1(_00450__PTR0), .A2(_00450__PTR1), .ZN(_00451_) );
  OR2_X1 U701 ( .A1(_00451_), .A2(_02097__PTR135), .ZN(_02099__PTR7) );
  OR2_X1 U702 ( .A1(_02097__PTR6), .A2(_02097__PTR38), .ZN(_00452__PTR0) );
  OR2_X1 U703 ( .A1(_02097__PTR70), .A2(_02097__PTR102), .ZN(_00452__PTR1) );
  OR2_X1 U704 ( .A1(_00452__PTR0), .A2(_00452__PTR1), .ZN(_00453_) );
  OR2_X1 U705 ( .A1(_00453_), .A2(_02097__PTR134), .ZN(_02099__PTR6) );
  OR2_X1 U706 ( .A1(_02097__PTR5), .A2(_02097__PTR37), .ZN(_00454__PTR0) );
  OR2_X1 U707 ( .A1(_02097__PTR69), .A2(_02097__PTR101), .ZN(_00454__PTR1) );
  OR2_X1 U708 ( .A1(_00454__PTR0), .A2(_00454__PTR1), .ZN(_00455_) );
  OR2_X1 U709 ( .A1(_00455_), .A2(_02097__PTR133), .ZN(_02099__PTR5) );
  OR2_X1 U710 ( .A1(_02097__PTR4), .A2(_02097__PTR36), .ZN(_00456__PTR0) );
  OR2_X1 U711 ( .A1(_02097__PTR68), .A2(_02097__PTR100), .ZN(_00456__PTR1) );
  OR2_X1 U712 ( .A1(_00456__PTR0), .A2(_00456__PTR1), .ZN(_00457_) );
  OR2_X1 U713 ( .A1(_00457_), .A2(_02097__PTR132), .ZN(_02099__PTR4) );
  OR2_X1 U714 ( .A1(_02097__PTR3), .A2(_02097__PTR35), .ZN(_00458__PTR0) );
  OR2_X1 U715 ( .A1(_02097__PTR67), .A2(_02097__PTR99), .ZN(_00458__PTR1) );
  OR2_X1 U716 ( .A1(_00458__PTR0), .A2(_00458__PTR1), .ZN(_00459_) );
  OR2_X1 U717 ( .A1(_00459_), .A2(_02097__PTR131), .ZN(_02099__PTR3) );
  OR2_X1 U718 ( .A1(_02097__PTR2), .A2(_02097__PTR34), .ZN(_00460__PTR0) );
  OR2_X1 U719 ( .A1(_02097__PTR66), .A2(_02097__PTR98), .ZN(_00460__PTR1) );
  OR2_X1 U720 ( .A1(_00460__PTR0), .A2(_00460__PTR1), .ZN(_00461_) );
  OR2_X1 U721 ( .A1(_00461_), .A2(_02097__PTR130), .ZN(_02099__PTR2) );
  OR2_X1 U722 ( .A1(_02097__PTR1), .A2(_02097__PTR33), .ZN(_00462__PTR0) );
  OR2_X1 U723 ( .A1(_02097__PTR65), .A2(_02097__PTR97), .ZN(_00462__PTR1) );
  OR2_X1 U724 ( .A1(_00462__PTR0), .A2(_00462__PTR1), .ZN(_00463_) );
  OR2_X1 U725 ( .A1(_00463_), .A2(_02097__PTR129), .ZN(_02099__PTR1) );
  OR2_X1 U726 ( .A1(_02097__PTR0), .A2(_02097__PTR32), .ZN(_00464__PTR0) );
  OR2_X1 U727 ( .A1(_02097__PTR64), .A2(_02097__PTR96), .ZN(_00464__PTR1) );
  OR2_X1 U728 ( .A1(_00464__PTR0), .A2(_00464__PTR1), .ZN(_00465_) );
  OR2_X1 U729 ( .A1(_00465_), .A2(_02097__PTR128), .ZN(_02099__PTR0) );
  OR2_X1 U730 ( .A1(_02098__PTR0), .A2(_02098__PTR1), .ZN(_00466__PTR0) );
  OR2_X1 U731 ( .A1(_02090__PTR3), .A2(_02090__PTR4), .ZN(_01855__PTR1) );
  OR2_X1 U732 ( .A1(_00466__PTR0), .A2(_01855__PTR1), .ZN(_00467_) );
  OR2_X1 U733 ( .A1(_00467_), .A2(_02098__PTR4), .ZN(_02923_) );
  OR2_X1 U734 ( .A1(_01858__PTR0), .A2(_01858__PTR1), .ZN(_00468__PTR0) );
  OR2_X1 U735 ( .A1(_01858__PTR2), .A2(_01858__PTR3), .ZN(_00468__PTR1) );
  OR2_X1 U736 ( .A1(_00468__PTR0), .A2(_00468__PTR1), .ZN(_01860_) );
  OR2_X1 U737 ( .A1(_00469__PTR0), .A2(_00469__PTR1), .ZN(_02773_) );
  OR2_X1 U738 ( .A1(_01854__PTR0), .A2(_01854__PTR1), .ZN(_00470__PTR0) );
  OR2_X1 U739 ( .A1(_01854__PTR2), .A2(_01854__PTR3), .ZN(_00470__PTR1) );
  OR2_X1 U740 ( .A1(_00470__PTR0), .A2(_00470__PTR1), .ZN(_01856_) );
  OR2_X1 U741 ( .A1(_01855__PTR2), .A2(_01855__PTR3), .ZN(_02090__PTR6) );
  OR2_X1 U742 ( .A1(_00469__PTR0), .A2(_02090__PTR6), .ZN(_02772_) );
  OR2_X1 U743 ( .A1(_02089__PTR14), .A2(_02089__PTR19), .ZN(_00471__PTR1) );
  OR2_X1 U744 ( .A1(_02089__PTR24), .A2(_02089__PTR29), .ZN(_00471__PTR2) );
  OR2_X1 U745 ( .A1(_00471__PTR2), .A2(_02089__PTR34), .ZN(_00472__PTR1) );
  OR2_X1 U746 ( .A1(_00471__PTR1), .A2(_00472__PTR1), .ZN(_02091__PTR4) );
  OR2_X1 U747 ( .A1(_02089__PTR3), .A2(_02089__PTR8), .ZN(_00473__PTR0) );
  OR2_X1 U748 ( .A1(_02089__PTR13), .A2(_02089__PTR18), .ZN(_00473__PTR1) );
  OR2_X1 U749 ( .A1(_02089__PTR23), .A2(_02089__PTR28), .ZN(_00473__PTR2) );
  OR2_X1 U750 ( .A1(_00473__PTR0), .A2(_00473__PTR1), .ZN(_00474__PTR0) );
  OR2_X1 U751 ( .A1(_00473__PTR2), .A2(_02089__PTR33), .ZN(_00474__PTR1) );
  OR2_X1 U752 ( .A1(_00474__PTR0), .A2(_00474__PTR1), .ZN(_02091__PTR3) );
  OR2_X1 U753 ( .A1(_02089__PTR2), .A2(_02089__PTR7), .ZN(_00475__PTR0) );
  OR2_X1 U754 ( .A1(_02089__PTR12), .A2(_02089__PTR17), .ZN(_00475__PTR1) );
  OR2_X1 U755 ( .A1(_02089__PTR22), .A2(_02089__PTR27), .ZN(_00475__PTR2) );
  OR2_X1 U756 ( .A1(_00475__PTR0), .A2(_00475__PTR1), .ZN(_00476__PTR0) );
  OR2_X1 U757 ( .A1(_00475__PTR2), .A2(_02089__PTR32), .ZN(_00476__PTR1) );
  OR2_X1 U758 ( .A1(_00476__PTR0), .A2(_00476__PTR1), .ZN(_02091__PTR2) );
  OR2_X1 U759 ( .A1(_02089__PTR1), .A2(_02089__PTR6), .ZN(_00477__PTR0) );
  OR2_X1 U760 ( .A1(_02089__PTR11), .A2(_02089__PTR16), .ZN(_00477__PTR1) );
  OR2_X1 U761 ( .A1(_02089__PTR21), .A2(_02089__PTR26), .ZN(_00477__PTR2) );
  OR2_X1 U762 ( .A1(_00477__PTR0), .A2(_00477__PTR1), .ZN(_00478__PTR0) );
  OR2_X1 U763 ( .A1(_00477__PTR2), .A2(_02089__PTR31), .ZN(_00478__PTR1) );
  OR2_X1 U764 ( .A1(_00478__PTR0), .A2(_00478__PTR1), .ZN(_02091__PTR1) );
  OR2_X1 U765 ( .A1(_02089__PTR0), .A2(_02089__PTR5), .ZN(_00479__PTR0) );
  OR2_X1 U766 ( .A1(_02089__PTR10), .A2(_02089__PTR15), .ZN(_00479__PTR1) );
  OR2_X1 U767 ( .A1(_02089__PTR20), .A2(_02089__PTR25), .ZN(_00479__PTR2) );
  OR2_X1 U768 ( .A1(_00479__PTR0), .A2(_00479__PTR1), .ZN(_00480__PTR0) );
  OR2_X1 U769 ( .A1(_00479__PTR2), .A2(_02089__PTR30), .ZN(_00480__PTR1) );
  OR2_X1 U770 ( .A1(_00480__PTR0), .A2(_00480__PTR1), .ZN(_02091__PTR0) );
  OR2_X1 U771 ( .A1(_01855__PTR0), .A2(_02090__PTR3), .ZN(_00481__PTR1) );
  OR2_X1 U772 ( .A1(_02090__PTR4), .A2(_02086__PTR4), .ZN(_00481__PTR2) );
  OR2_X1 U773 ( .A1(_00481__PTR0), .A2(_00481__PTR1), .ZN(_00482__PTR0) );
  OR2_X1 U774 ( .A1(_00481__PTR2), .A2(_02090__PTR6), .ZN(_00482__PTR1) );
  OR2_X1 U775 ( .A1(_00482__PTR0), .A2(_00482__PTR1), .ZN(_02921_) );
  OR2_X1 U776 ( .A1(_01873__PTR0), .A2(_01873__PTR1), .ZN(_01875_) );
  OR2_X1 U777 ( .A1(_01862__PTR0), .A2(_01862__PTR1), .ZN(_00483__PTR0) );
  OR2_X1 U778 ( .A1(_01862__PTR2), .A2(_01862__PTR3), .ZN(_00483__PTR1) );
  OR2_X1 U779 ( .A1(_00483__PTR0), .A2(_00483__PTR1), .ZN(_01864_) );
  OR2_X1 U780 ( .A1(_01863__PTR0), .A2(_01855__PTR1), .ZN(_00484__PTR0) );
  OR2_X1 U781 ( .A1(_01863__PTR2), .A2(_01863__PTR3), .ZN(_00484__PTR1) );
  OR2_X1 U782 ( .A1(_00484__PTR0), .A2(_00484__PTR1), .ZN(_02774_) );
  OR2_X1 U783 ( .A1(_01869__PTR0), .A2(_01869__PTR1), .ZN(_00485_) );
  OR2_X1 U784 ( .A1(_00485_), .A2(_01869__PTR2), .ZN(_01871_) );
  OR2_X1 U785 ( .A1(_01870__PTR0), .A2(_01870__PTR1), .ZN(_01874__PTR0) );
  OR2_X1 U786 ( .A1(_01874__PTR0), .A2(_01863__PTR3), .ZN(_02776_) );
  OR2_X1 U787 ( .A1(_01866__PTR0), .A2(_01866__PTR1), .ZN(_00486_) );
  OR2_X1 U788 ( .A1(_00486_), .A2(_01866__PTR2), .ZN(_01867_) );
  OR2_X1 U789 ( .A1(_00469__PTR0), .A2(_01863__PTR3), .ZN(_02775_) );
  OR2_X1 U790 ( .A1(_02105__PTR31), .A2(_02105__PTR63), .ZN(_00487__PTR0) );
  OR2_X1 U791 ( .A1(_02105__PTR95), .A2(_02105__PTR127), .ZN(_00487__PTR1) );
  OR2_X1 U792 ( .A1(_00487__PTR0), .A2(_00487__PTR1), .ZN(_02106__PTR31) );
  OR2_X1 U793 ( .A1(_02105__PTR30), .A2(_02105__PTR62), .ZN(_00488__PTR0) );
  OR2_X1 U794 ( .A1(_02105__PTR94), .A2(_02105__PTR126), .ZN(_00488__PTR1) );
  OR2_X1 U795 ( .A1(_00488__PTR0), .A2(_00488__PTR1), .ZN(_02106__PTR30) );
  OR2_X1 U796 ( .A1(_02105__PTR29), .A2(_02105__PTR61), .ZN(_00489__PTR0) );
  OR2_X1 U797 ( .A1(_02105__PTR93), .A2(_02105__PTR125), .ZN(_00489__PTR1) );
  OR2_X1 U798 ( .A1(_00489__PTR0), .A2(_00489__PTR1), .ZN(_02106__PTR29) );
  OR2_X1 U799 ( .A1(_02105__PTR28), .A2(_02105__PTR60), .ZN(_00490__PTR0) );
  OR2_X1 U800 ( .A1(_02105__PTR92), .A2(_02105__PTR124), .ZN(_00490__PTR1) );
  OR2_X1 U801 ( .A1(_00490__PTR0), .A2(_00490__PTR1), .ZN(_02106__PTR28) );
  OR2_X1 U802 ( .A1(_02105__PTR27), .A2(_02105__PTR59), .ZN(_00491__PTR0) );
  OR2_X1 U803 ( .A1(_02105__PTR91), .A2(_02105__PTR123), .ZN(_00491__PTR1) );
  OR2_X1 U804 ( .A1(_00491__PTR0), .A2(_00491__PTR1), .ZN(_02106__PTR27) );
  OR2_X1 U805 ( .A1(_02105__PTR26), .A2(_02105__PTR58), .ZN(_00492__PTR0) );
  OR2_X1 U806 ( .A1(_02105__PTR90), .A2(_02105__PTR122), .ZN(_00492__PTR1) );
  OR2_X1 U807 ( .A1(_00492__PTR0), .A2(_00492__PTR1), .ZN(_02106__PTR26) );
  OR2_X1 U808 ( .A1(_02105__PTR25), .A2(_02105__PTR57), .ZN(_00493__PTR0) );
  OR2_X1 U809 ( .A1(_02105__PTR89), .A2(_02105__PTR121), .ZN(_00493__PTR1) );
  OR2_X1 U810 ( .A1(_00493__PTR0), .A2(_00493__PTR1), .ZN(_02106__PTR25) );
  OR2_X1 U811 ( .A1(_02105__PTR24), .A2(_02105__PTR56), .ZN(_00494__PTR0) );
  OR2_X1 U812 ( .A1(_02105__PTR88), .A2(_02105__PTR120), .ZN(_00494__PTR1) );
  OR2_X1 U813 ( .A1(_00494__PTR0), .A2(_00494__PTR1), .ZN(_02106__PTR24) );
  OR2_X1 U814 ( .A1(_02105__PTR23), .A2(_02105__PTR55), .ZN(_00495__PTR0) );
  OR2_X1 U815 ( .A1(_02105__PTR87), .A2(_02105__PTR119), .ZN(_00495__PTR1) );
  OR2_X1 U816 ( .A1(_00495__PTR0), .A2(_00495__PTR1), .ZN(_02106__PTR23) );
  OR2_X1 U817 ( .A1(_02105__PTR22), .A2(_02105__PTR54), .ZN(_00496__PTR0) );
  OR2_X1 U818 ( .A1(_02105__PTR86), .A2(_02105__PTR118), .ZN(_00496__PTR1) );
  OR2_X1 U819 ( .A1(_00496__PTR0), .A2(_00496__PTR1), .ZN(_02106__PTR22) );
  OR2_X1 U820 ( .A1(_02105__PTR21), .A2(_02105__PTR53), .ZN(_00497__PTR0) );
  OR2_X1 U821 ( .A1(_02105__PTR85), .A2(_02105__PTR117), .ZN(_00497__PTR1) );
  OR2_X1 U822 ( .A1(_00497__PTR0), .A2(_00497__PTR1), .ZN(_02106__PTR21) );
  OR2_X1 U823 ( .A1(_02105__PTR20), .A2(_02105__PTR52), .ZN(_00498__PTR0) );
  OR2_X1 U824 ( .A1(_02105__PTR84), .A2(_02105__PTR116), .ZN(_00498__PTR1) );
  OR2_X1 U825 ( .A1(_00498__PTR0), .A2(_00498__PTR1), .ZN(_02106__PTR20) );
  OR2_X1 U826 ( .A1(_02105__PTR19), .A2(_02105__PTR51), .ZN(_00499__PTR0) );
  OR2_X1 U827 ( .A1(_02105__PTR83), .A2(_02105__PTR115), .ZN(_00499__PTR1) );
  OR2_X1 U828 ( .A1(_00499__PTR0), .A2(_00499__PTR1), .ZN(_02106__PTR19) );
  OR2_X1 U829 ( .A1(_02105__PTR18), .A2(_02105__PTR50), .ZN(_00500__PTR0) );
  OR2_X1 U830 ( .A1(_02105__PTR82), .A2(_02105__PTR114), .ZN(_00500__PTR1) );
  OR2_X1 U831 ( .A1(_00500__PTR0), .A2(_00500__PTR1), .ZN(_02106__PTR18) );
  OR2_X1 U832 ( .A1(_02105__PTR17), .A2(_02105__PTR49), .ZN(_00501__PTR0) );
  OR2_X1 U833 ( .A1(_02105__PTR81), .A2(_02105__PTR113), .ZN(_00501__PTR1) );
  OR2_X1 U834 ( .A1(_00501__PTR0), .A2(_00501__PTR1), .ZN(_02106__PTR17) );
  OR2_X1 U835 ( .A1(_02105__PTR16), .A2(_02105__PTR48), .ZN(_00502__PTR0) );
  OR2_X1 U836 ( .A1(_02105__PTR80), .A2(_02105__PTR112), .ZN(_00502__PTR1) );
  OR2_X1 U837 ( .A1(_00502__PTR0), .A2(_00502__PTR1), .ZN(_02106__PTR16) );
  OR2_X1 U838 ( .A1(_02105__PTR15), .A2(_02105__PTR47), .ZN(_00503__PTR0) );
  OR2_X1 U839 ( .A1(_02105__PTR79), .A2(_02105__PTR111), .ZN(_00503__PTR1) );
  OR2_X1 U840 ( .A1(_00503__PTR0), .A2(_00503__PTR1), .ZN(_02106__PTR15) );
  OR2_X1 U841 ( .A1(_02105__PTR14), .A2(_02105__PTR46), .ZN(_00504__PTR0) );
  OR2_X1 U842 ( .A1(_02105__PTR78), .A2(_02105__PTR110), .ZN(_00504__PTR1) );
  OR2_X1 U843 ( .A1(_00504__PTR0), .A2(_00504__PTR1), .ZN(_02106__PTR14) );
  OR2_X1 U844 ( .A1(_02105__PTR13), .A2(_02105__PTR45), .ZN(_00505__PTR0) );
  OR2_X1 U845 ( .A1(_02105__PTR77), .A2(_02105__PTR109), .ZN(_00505__PTR1) );
  OR2_X1 U846 ( .A1(_00505__PTR0), .A2(_00505__PTR1), .ZN(_02106__PTR13) );
  OR2_X1 U847 ( .A1(_02105__PTR12), .A2(_02105__PTR44), .ZN(_00506__PTR0) );
  OR2_X1 U848 ( .A1(_02105__PTR76), .A2(_02105__PTR108), .ZN(_00506__PTR1) );
  OR2_X1 U849 ( .A1(_00506__PTR0), .A2(_00506__PTR1), .ZN(_02106__PTR12) );
  OR2_X1 U850 ( .A1(_02105__PTR11), .A2(_02105__PTR43), .ZN(_00507__PTR0) );
  OR2_X1 U851 ( .A1(_02105__PTR75), .A2(_02105__PTR107), .ZN(_00507__PTR1) );
  OR2_X1 U852 ( .A1(_00507__PTR0), .A2(_00507__PTR1), .ZN(_02106__PTR11) );
  OR2_X1 U853 ( .A1(_02105__PTR10), .A2(_02105__PTR42), .ZN(_00508__PTR0) );
  OR2_X1 U854 ( .A1(_02105__PTR74), .A2(_02105__PTR106), .ZN(_00508__PTR1) );
  OR2_X1 U855 ( .A1(_00508__PTR0), .A2(_00508__PTR1), .ZN(_02106__PTR10) );
  OR2_X1 U856 ( .A1(_02105__PTR9), .A2(_02105__PTR41), .ZN(_00509__PTR0) );
  OR2_X1 U857 ( .A1(_02105__PTR73), .A2(_02105__PTR105), .ZN(_00509__PTR1) );
  OR2_X1 U858 ( .A1(_00509__PTR0), .A2(_00509__PTR1), .ZN(_02106__PTR9) );
  OR2_X1 U859 ( .A1(_02105__PTR8), .A2(_02105__PTR40), .ZN(_00510__PTR0) );
  OR2_X1 U860 ( .A1(_02105__PTR72), .A2(_02105__PTR104), .ZN(_00510__PTR1) );
  OR2_X1 U861 ( .A1(_00510__PTR0), .A2(_00510__PTR1), .ZN(_02106__PTR8) );
  OR2_X1 U862 ( .A1(_02105__PTR7), .A2(_02105__PTR39), .ZN(_00511__PTR0) );
  OR2_X1 U863 ( .A1(_02105__PTR71), .A2(_02105__PTR103), .ZN(_00511__PTR1) );
  OR2_X1 U864 ( .A1(_00511__PTR0), .A2(_00511__PTR1), .ZN(_02106__PTR7) );
  OR2_X1 U865 ( .A1(_02105__PTR6), .A2(_02105__PTR38), .ZN(_00512__PTR0) );
  OR2_X1 U866 ( .A1(_02105__PTR70), .A2(_02105__PTR102), .ZN(_00512__PTR1) );
  OR2_X1 U867 ( .A1(_00512__PTR0), .A2(_00512__PTR1), .ZN(_02106__PTR6) );
  OR2_X1 U868 ( .A1(_02105__PTR5), .A2(_02105__PTR37), .ZN(_00513__PTR0) );
  OR2_X1 U869 ( .A1(_02105__PTR69), .A2(_02105__PTR101), .ZN(_00513__PTR1) );
  OR2_X1 U870 ( .A1(_00513__PTR0), .A2(_00513__PTR1), .ZN(_02106__PTR5) );
  OR2_X1 U871 ( .A1(_02105__PTR4), .A2(_02105__PTR36), .ZN(_00514__PTR0) );
  OR2_X1 U872 ( .A1(_02105__PTR68), .A2(_02105__PTR100), .ZN(_00514__PTR1) );
  OR2_X1 U873 ( .A1(_00514__PTR0), .A2(_00514__PTR1), .ZN(_02106__PTR4) );
  OR2_X1 U874 ( .A1(_02105__PTR3), .A2(_02105__PTR35), .ZN(_00515__PTR0) );
  OR2_X1 U875 ( .A1(_02105__PTR67), .A2(_02105__PTR99), .ZN(_00515__PTR1) );
  OR2_X1 U876 ( .A1(_00515__PTR0), .A2(_00515__PTR1), .ZN(_02106__PTR3) );
  OR2_X1 U877 ( .A1(_02105__PTR2), .A2(_02105__PTR34), .ZN(_00516__PTR0) );
  OR2_X1 U878 ( .A1(_02105__PTR66), .A2(_02105__PTR98), .ZN(_00516__PTR1) );
  OR2_X1 U879 ( .A1(_00516__PTR0), .A2(_00516__PTR1), .ZN(_02106__PTR2) );
  OR2_X1 U880 ( .A1(_02105__PTR1), .A2(_02105__PTR33), .ZN(_00517__PTR0) );
  OR2_X1 U881 ( .A1(_02105__PTR65), .A2(_02105__PTR97), .ZN(_00517__PTR1) );
  OR2_X1 U882 ( .A1(_00517__PTR0), .A2(_00517__PTR1), .ZN(_02106__PTR1) );
  OR2_X1 U883 ( .A1(_02105__PTR0), .A2(_02105__PTR32), .ZN(_00518__PTR0) );
  OR2_X1 U884 ( .A1(_02105__PTR64), .A2(_02105__PTR96), .ZN(_00518__PTR1) );
  OR2_X1 U885 ( .A1(_00518__PTR0), .A2(_00518__PTR1), .ZN(_02106__PTR0) );
  OR2_X1 U886 ( .A1(_01863__PTR3), .A2(_01870__PTR0), .ZN(_00519__PTR0) );
  OR2_X1 U887 ( .A1(_01863__PTR2), .A2(_02090__PTR4), .ZN(_01870__PTR1) );
  OR2_X1 U888 ( .A1(_00519__PTR0), .A2(_01870__PTR1), .ZN(_02925_) );
  OR2_X1 U889 ( .A1(_02085__PTR31), .A2(_02085__PTR63), .ZN(_00520__PTR0) );
  OR2_X1 U890 ( .A1(_02085__PTR95), .A2(_02085__PTR127), .ZN(_00520__PTR1) );
  OR2_X1 U891 ( .A1(_02085__PTR159), .A2(_02085__PTR191), .ZN(_00520__PTR2) );
  OR2_X1 U892 ( .A1(_00520__PTR0), .A2(_00520__PTR1), .ZN(_00521__PTR0) );
  OR2_X1 U893 ( .A1(_00520__PTR2), .A2(_02085__PTR223), .ZN(_00521__PTR1) );
  OR2_X1 U894 ( .A1(_00521__PTR0), .A2(_00521__PTR1), .ZN(_02087__PTR31) );
  OR2_X1 U895 ( .A1(_02085__PTR30), .A2(_02085__PTR62), .ZN(_00522__PTR0) );
  OR2_X1 U896 ( .A1(_02085__PTR94), .A2(_02085__PTR126), .ZN(_00522__PTR1) );
  OR2_X1 U897 ( .A1(_02085__PTR158), .A2(_02085__PTR190), .ZN(_00522__PTR2) );
  OR2_X1 U898 ( .A1(_00522__PTR0), .A2(_00522__PTR1), .ZN(_00523__PTR0) );
  OR2_X1 U899 ( .A1(_00522__PTR2), .A2(_02085__PTR222), .ZN(_00523__PTR1) );
  OR2_X1 U900 ( .A1(_00523__PTR0), .A2(_00523__PTR1), .ZN(_02087__PTR30) );
  OR2_X1 U901 ( .A1(_02085__PTR29), .A2(_02085__PTR61), .ZN(_00524__PTR0) );
  OR2_X1 U902 ( .A1(_02085__PTR93), .A2(_02085__PTR125), .ZN(_00524__PTR1) );
  OR2_X1 U903 ( .A1(_02085__PTR157), .A2(_02085__PTR189), .ZN(_00524__PTR2) );
  OR2_X1 U904 ( .A1(_00524__PTR0), .A2(_00524__PTR1), .ZN(_00525__PTR0) );
  OR2_X1 U905 ( .A1(_00524__PTR2), .A2(_02085__PTR221), .ZN(_00525__PTR1) );
  OR2_X1 U906 ( .A1(_00525__PTR0), .A2(_00525__PTR1), .ZN(_02087__PTR29) );
  OR2_X1 U907 ( .A1(_02085__PTR28), .A2(_02085__PTR60), .ZN(_00526__PTR0) );
  OR2_X1 U908 ( .A1(_02085__PTR92), .A2(_02085__PTR124), .ZN(_00526__PTR1) );
  OR2_X1 U909 ( .A1(_02085__PTR156), .A2(_02085__PTR188), .ZN(_00526__PTR2) );
  OR2_X1 U910 ( .A1(_00526__PTR0), .A2(_00526__PTR1), .ZN(_00527__PTR0) );
  OR2_X1 U911 ( .A1(_00526__PTR2), .A2(_02085__PTR220), .ZN(_00527__PTR1) );
  OR2_X1 U912 ( .A1(_00527__PTR0), .A2(_00527__PTR1), .ZN(_02087__PTR28) );
  OR2_X1 U913 ( .A1(_02085__PTR27), .A2(_02085__PTR59), .ZN(_00528__PTR0) );
  OR2_X1 U914 ( .A1(_02085__PTR91), .A2(_02085__PTR123), .ZN(_00528__PTR1) );
  OR2_X1 U915 ( .A1(_02085__PTR155), .A2(_02085__PTR187), .ZN(_00528__PTR2) );
  OR2_X1 U916 ( .A1(_00528__PTR0), .A2(_00528__PTR1), .ZN(_00529__PTR0) );
  OR2_X1 U917 ( .A1(_00528__PTR2), .A2(_02085__PTR219), .ZN(_00529__PTR1) );
  OR2_X1 U918 ( .A1(_00529__PTR0), .A2(_00529__PTR1), .ZN(_02087__PTR27) );
  OR2_X1 U919 ( .A1(_02085__PTR26), .A2(_02085__PTR58), .ZN(_00530__PTR0) );
  OR2_X1 U920 ( .A1(_02085__PTR90), .A2(_02085__PTR122), .ZN(_00530__PTR1) );
  OR2_X1 U921 ( .A1(_02085__PTR154), .A2(_02085__PTR186), .ZN(_00530__PTR2) );
  OR2_X1 U922 ( .A1(_00530__PTR0), .A2(_00530__PTR1), .ZN(_00531__PTR0) );
  OR2_X1 U923 ( .A1(_00530__PTR2), .A2(_02085__PTR218), .ZN(_00531__PTR1) );
  OR2_X1 U924 ( .A1(_00531__PTR0), .A2(_00531__PTR1), .ZN(_02087__PTR26) );
  OR2_X1 U925 ( .A1(_02085__PTR25), .A2(_02085__PTR57), .ZN(_00532__PTR0) );
  OR2_X1 U926 ( .A1(_02085__PTR89), .A2(_02085__PTR121), .ZN(_00532__PTR1) );
  OR2_X1 U927 ( .A1(_02085__PTR153), .A2(_02085__PTR185), .ZN(_00532__PTR2) );
  OR2_X1 U928 ( .A1(_00532__PTR0), .A2(_00532__PTR1), .ZN(_00533__PTR0) );
  OR2_X1 U929 ( .A1(_00532__PTR2), .A2(_02085__PTR217), .ZN(_00533__PTR1) );
  OR2_X1 U930 ( .A1(_00533__PTR0), .A2(_00533__PTR1), .ZN(_02087__PTR25) );
  OR2_X1 U931 ( .A1(_02085__PTR24), .A2(_02085__PTR56), .ZN(_00534__PTR0) );
  OR2_X1 U932 ( .A1(_02085__PTR88), .A2(_02085__PTR120), .ZN(_00534__PTR1) );
  OR2_X1 U933 ( .A1(_02085__PTR152), .A2(_02085__PTR184), .ZN(_00534__PTR2) );
  OR2_X1 U934 ( .A1(_00534__PTR0), .A2(_00534__PTR1), .ZN(_00535__PTR0) );
  OR2_X1 U935 ( .A1(_00534__PTR2), .A2(_02085__PTR216), .ZN(_00535__PTR1) );
  OR2_X1 U936 ( .A1(_00535__PTR0), .A2(_00535__PTR1), .ZN(_02087__PTR24) );
  OR2_X1 U937 ( .A1(_02085__PTR23), .A2(_02085__PTR55), .ZN(_00536__PTR0) );
  OR2_X1 U938 ( .A1(_02085__PTR87), .A2(_02085__PTR119), .ZN(_00536__PTR1) );
  OR2_X1 U939 ( .A1(_02085__PTR151), .A2(_02085__PTR183), .ZN(_00536__PTR2) );
  OR2_X1 U940 ( .A1(_00536__PTR0), .A2(_00536__PTR1), .ZN(_00537__PTR0) );
  OR2_X1 U941 ( .A1(_00536__PTR2), .A2(_02085__PTR215), .ZN(_00537__PTR1) );
  OR2_X1 U942 ( .A1(_00537__PTR0), .A2(_00537__PTR1), .ZN(_02087__PTR23) );
  OR2_X1 U943 ( .A1(_02085__PTR22), .A2(_02085__PTR54), .ZN(_00538__PTR0) );
  OR2_X1 U944 ( .A1(_02085__PTR86), .A2(_02085__PTR118), .ZN(_00538__PTR1) );
  OR2_X1 U945 ( .A1(_02085__PTR150), .A2(_02085__PTR182), .ZN(_00538__PTR2) );
  OR2_X1 U946 ( .A1(_00538__PTR0), .A2(_00538__PTR1), .ZN(_00539__PTR0) );
  OR2_X1 U947 ( .A1(_00538__PTR2), .A2(_02085__PTR214), .ZN(_00539__PTR1) );
  OR2_X1 U948 ( .A1(_00539__PTR0), .A2(_00539__PTR1), .ZN(_02087__PTR22) );
  OR2_X1 U949 ( .A1(_02085__PTR21), .A2(_02085__PTR53), .ZN(_00540__PTR0) );
  OR2_X1 U950 ( .A1(_02085__PTR85), .A2(_02085__PTR117), .ZN(_00540__PTR1) );
  OR2_X1 U951 ( .A1(_02085__PTR149), .A2(_02085__PTR181), .ZN(_00540__PTR2) );
  OR2_X1 U952 ( .A1(_00540__PTR0), .A2(_00540__PTR1), .ZN(_00541__PTR0) );
  OR2_X1 U953 ( .A1(_00540__PTR2), .A2(_02085__PTR213), .ZN(_00541__PTR1) );
  OR2_X1 U954 ( .A1(_00541__PTR0), .A2(_00541__PTR1), .ZN(_02087__PTR21) );
  OR2_X1 U955 ( .A1(_02085__PTR20), .A2(_02085__PTR52), .ZN(_00542__PTR0) );
  OR2_X1 U956 ( .A1(_02085__PTR84), .A2(_02085__PTR116), .ZN(_00542__PTR1) );
  OR2_X1 U957 ( .A1(_02085__PTR148), .A2(_02085__PTR180), .ZN(_00542__PTR2) );
  OR2_X1 U958 ( .A1(_00542__PTR0), .A2(_00542__PTR1), .ZN(_00543__PTR0) );
  OR2_X1 U959 ( .A1(_00542__PTR2), .A2(_02085__PTR212), .ZN(_00543__PTR1) );
  OR2_X1 U960 ( .A1(_00543__PTR0), .A2(_00543__PTR1), .ZN(_02087__PTR20) );
  OR2_X1 U961 ( .A1(_02085__PTR19), .A2(_02085__PTR51), .ZN(_00544__PTR0) );
  OR2_X1 U962 ( .A1(_02085__PTR83), .A2(_02085__PTR115), .ZN(_00544__PTR1) );
  OR2_X1 U963 ( .A1(_02085__PTR147), .A2(_02085__PTR179), .ZN(_00544__PTR2) );
  OR2_X1 U964 ( .A1(_00544__PTR0), .A2(_00544__PTR1), .ZN(_00545__PTR0) );
  OR2_X1 U965 ( .A1(_00544__PTR2), .A2(_02085__PTR211), .ZN(_00545__PTR1) );
  OR2_X1 U966 ( .A1(_00545__PTR0), .A2(_00545__PTR1), .ZN(_02087__PTR19) );
  OR2_X1 U967 ( .A1(_02085__PTR18), .A2(_02085__PTR50), .ZN(_00546__PTR0) );
  OR2_X1 U968 ( .A1(_02085__PTR82), .A2(_02085__PTR114), .ZN(_00546__PTR1) );
  OR2_X1 U969 ( .A1(_02085__PTR146), .A2(_02085__PTR178), .ZN(_00546__PTR2) );
  OR2_X1 U970 ( .A1(_00546__PTR0), .A2(_00546__PTR1), .ZN(_00547__PTR0) );
  OR2_X1 U971 ( .A1(_00546__PTR2), .A2(_02085__PTR210), .ZN(_00547__PTR1) );
  OR2_X1 U972 ( .A1(_00547__PTR0), .A2(_00547__PTR1), .ZN(_02087__PTR18) );
  OR2_X1 U973 ( .A1(_02085__PTR17), .A2(_02085__PTR49), .ZN(_00548__PTR0) );
  OR2_X1 U974 ( .A1(_02085__PTR81), .A2(_02085__PTR113), .ZN(_00548__PTR1) );
  OR2_X1 U975 ( .A1(_02085__PTR145), .A2(_02085__PTR177), .ZN(_00548__PTR2) );
  OR2_X1 U976 ( .A1(_00548__PTR0), .A2(_00548__PTR1), .ZN(_00549__PTR0) );
  OR2_X1 U977 ( .A1(_00548__PTR2), .A2(_02085__PTR209), .ZN(_00549__PTR1) );
  OR2_X1 U978 ( .A1(_00549__PTR0), .A2(_00549__PTR1), .ZN(_02087__PTR17) );
  OR2_X1 U979 ( .A1(_02085__PTR16), .A2(_02085__PTR48), .ZN(_00550__PTR0) );
  OR2_X1 U980 ( .A1(_02085__PTR80), .A2(_02085__PTR112), .ZN(_00550__PTR1) );
  OR2_X1 U981 ( .A1(_02085__PTR144), .A2(_02085__PTR176), .ZN(_00550__PTR2) );
  OR2_X1 U982 ( .A1(_00550__PTR0), .A2(_00550__PTR1), .ZN(_00551__PTR0) );
  OR2_X1 U983 ( .A1(_00550__PTR2), .A2(_02085__PTR208), .ZN(_00551__PTR1) );
  OR2_X1 U984 ( .A1(_00551__PTR0), .A2(_00551__PTR1), .ZN(_02087__PTR16) );
  OR2_X1 U985 ( .A1(_02085__PTR15), .A2(_02085__PTR47), .ZN(_00552__PTR0) );
  OR2_X1 U986 ( .A1(_02085__PTR79), .A2(_02085__PTR111), .ZN(_00552__PTR1) );
  OR2_X1 U987 ( .A1(_02085__PTR143), .A2(_02085__PTR175), .ZN(_00552__PTR2) );
  OR2_X1 U988 ( .A1(_00552__PTR0), .A2(_00552__PTR1), .ZN(_00553__PTR0) );
  OR2_X1 U989 ( .A1(_00552__PTR2), .A2(_02085__PTR207), .ZN(_00553__PTR1) );
  OR2_X1 U990 ( .A1(_00553__PTR0), .A2(_00553__PTR1), .ZN(_02087__PTR15) );
  OR2_X1 U991 ( .A1(_02085__PTR14), .A2(_02085__PTR46), .ZN(_00554__PTR0) );
  OR2_X1 U992 ( .A1(_02085__PTR78), .A2(_02085__PTR110), .ZN(_00554__PTR1) );
  OR2_X1 U993 ( .A1(_02085__PTR142), .A2(_02085__PTR174), .ZN(_00554__PTR2) );
  OR2_X1 U994 ( .A1(_00554__PTR0), .A2(_00554__PTR1), .ZN(_00555__PTR0) );
  OR2_X1 U995 ( .A1(_00554__PTR2), .A2(_02085__PTR206), .ZN(_00555__PTR1) );
  OR2_X1 U996 ( .A1(_00555__PTR0), .A2(_00555__PTR1), .ZN(_02087__PTR14) );
  OR2_X1 U997 ( .A1(_02085__PTR13), .A2(_02085__PTR45), .ZN(_00556__PTR0) );
  OR2_X1 U998 ( .A1(_02085__PTR77), .A2(_02085__PTR109), .ZN(_00556__PTR1) );
  OR2_X1 U999 ( .A1(_02085__PTR141), .A2(_02085__PTR173), .ZN(_00556__PTR2) );
  OR2_X1 U1000 ( .A1(_00556__PTR0), .A2(_00556__PTR1), .ZN(_00557__PTR0) );
  OR2_X1 U1001 ( .A1(_00556__PTR2), .A2(_02085__PTR205), .ZN(_00557__PTR1) );
  OR2_X1 U1002 ( .A1(_00557__PTR0), .A2(_00557__PTR1), .ZN(_02087__PTR13) );
  OR2_X1 U1003 ( .A1(_02085__PTR12), .A2(_02085__PTR44), .ZN(_00558__PTR0) );
  OR2_X1 U1004 ( .A1(_02085__PTR76), .A2(_02085__PTR108), .ZN(_00558__PTR1) );
  OR2_X1 U1005 ( .A1(_02085__PTR140), .A2(_02085__PTR172), .ZN(_00558__PTR2) );
  OR2_X1 U1006 ( .A1(_00558__PTR0), .A2(_00558__PTR1), .ZN(_00559__PTR0) );
  OR2_X1 U1007 ( .A1(_00558__PTR2), .A2(_02085__PTR204), .ZN(_00559__PTR1) );
  OR2_X1 U1008 ( .A1(_00559__PTR0), .A2(_00559__PTR1), .ZN(_02087__PTR12) );
  OR2_X1 U1009 ( .A1(_02085__PTR11), .A2(_02085__PTR43), .ZN(_00560__PTR0) );
  OR2_X1 U1010 ( .A1(_02085__PTR75), .A2(_02085__PTR107), .ZN(_00560__PTR1) );
  OR2_X1 U1011 ( .A1(_02085__PTR139), .A2(_02085__PTR171), .ZN(_00560__PTR2) );
  OR2_X1 U1012 ( .A1(_00560__PTR0), .A2(_00560__PTR1), .ZN(_00561__PTR0) );
  OR2_X1 U1013 ( .A1(_00560__PTR2), .A2(_02085__PTR203), .ZN(_00561__PTR1) );
  OR2_X1 U1014 ( .A1(_00561__PTR0), .A2(_00561__PTR1), .ZN(_02087__PTR11) );
  OR2_X1 U1015 ( .A1(_02085__PTR10), .A2(_02085__PTR42), .ZN(_00562__PTR0) );
  OR2_X1 U1016 ( .A1(_02085__PTR74), .A2(_02085__PTR106), .ZN(_00562__PTR1) );
  OR2_X1 U1017 ( .A1(_02085__PTR138), .A2(_02085__PTR170), .ZN(_00562__PTR2) );
  OR2_X1 U1018 ( .A1(_00562__PTR0), .A2(_00562__PTR1), .ZN(_00563__PTR0) );
  OR2_X1 U1019 ( .A1(_00562__PTR2), .A2(_02085__PTR202), .ZN(_00563__PTR1) );
  OR2_X1 U1020 ( .A1(_00563__PTR0), .A2(_00563__PTR1), .ZN(_02087__PTR10) );
  OR2_X1 U1021 ( .A1(_02085__PTR9), .A2(_02085__PTR41), .ZN(_00564__PTR0) );
  OR2_X1 U1022 ( .A1(_02085__PTR73), .A2(_02085__PTR105), .ZN(_00564__PTR1) );
  OR2_X1 U1023 ( .A1(_02085__PTR137), .A2(_02085__PTR169), .ZN(_00564__PTR2) );
  OR2_X1 U1024 ( .A1(_00564__PTR0), .A2(_00564__PTR1), .ZN(_00565__PTR0) );
  OR2_X1 U1025 ( .A1(_00564__PTR2), .A2(_02085__PTR201), .ZN(_00565__PTR1) );
  OR2_X1 U1026 ( .A1(_00565__PTR0), .A2(_00565__PTR1), .ZN(_02087__PTR9) );
  OR2_X1 U1027 ( .A1(_02085__PTR8), .A2(_02085__PTR40), .ZN(_00566__PTR0) );
  OR2_X1 U1028 ( .A1(_02085__PTR72), .A2(_02085__PTR104), .ZN(_00566__PTR1) );
  OR2_X1 U1029 ( .A1(_02085__PTR136), .A2(_02085__PTR168), .ZN(_00566__PTR2) );
  OR2_X1 U1030 ( .A1(_00566__PTR0), .A2(_00566__PTR1), .ZN(_00567__PTR0) );
  OR2_X1 U1031 ( .A1(_00566__PTR2), .A2(_02085__PTR200), .ZN(_00567__PTR1) );
  OR2_X1 U1032 ( .A1(_00567__PTR0), .A2(_00567__PTR1), .ZN(_02087__PTR8) );
  OR2_X1 U1033 ( .A1(_02085__PTR7), .A2(_02085__PTR39), .ZN(_00568__PTR0) );
  OR2_X1 U1034 ( .A1(_02085__PTR71), .A2(_02085__PTR103), .ZN(_00568__PTR1) );
  OR2_X1 U1035 ( .A1(_02085__PTR135), .A2(_02085__PTR167), .ZN(_00568__PTR2) );
  OR2_X1 U1036 ( .A1(_00568__PTR0), .A2(_00568__PTR1), .ZN(_00569__PTR0) );
  OR2_X1 U1037 ( .A1(_00568__PTR2), .A2(_02085__PTR199), .ZN(_00569__PTR1) );
  OR2_X1 U1038 ( .A1(_00569__PTR0), .A2(_00569__PTR1), .ZN(_02087__PTR7) );
  OR2_X1 U1039 ( .A1(_02085__PTR6), .A2(_02085__PTR38), .ZN(_00570__PTR0) );
  OR2_X1 U1040 ( .A1(_02085__PTR70), .A2(_02085__PTR102), .ZN(_00570__PTR1) );
  OR2_X1 U1041 ( .A1(_02085__PTR134), .A2(_02085__PTR166), .ZN(_00570__PTR2) );
  OR2_X1 U1042 ( .A1(_00570__PTR0), .A2(_00570__PTR1), .ZN(_00571__PTR0) );
  OR2_X1 U1043 ( .A1(_00570__PTR2), .A2(_02085__PTR198), .ZN(_00571__PTR1) );
  OR2_X1 U1044 ( .A1(_00571__PTR0), .A2(_00571__PTR1), .ZN(_02087__PTR6) );
  OR2_X1 U1045 ( .A1(_02085__PTR5), .A2(_02085__PTR37), .ZN(_00572__PTR0) );
  OR2_X1 U1046 ( .A1(_02085__PTR69), .A2(_02085__PTR101), .ZN(_00572__PTR1) );
  OR2_X1 U1047 ( .A1(_02085__PTR133), .A2(_02085__PTR165), .ZN(_00572__PTR2) );
  OR2_X1 U1048 ( .A1(_00572__PTR0), .A2(_00572__PTR1), .ZN(_00573__PTR0) );
  OR2_X1 U1049 ( .A1(_00572__PTR2), .A2(_02085__PTR197), .ZN(_00573__PTR1) );
  OR2_X1 U1050 ( .A1(_00573__PTR0), .A2(_00573__PTR1), .ZN(_02087__PTR5) );
  OR2_X1 U1051 ( .A1(_02085__PTR4), .A2(_02085__PTR36), .ZN(_00574__PTR0) );
  OR2_X1 U1052 ( .A1(_02085__PTR68), .A2(_02085__PTR100), .ZN(_00574__PTR1) );
  OR2_X1 U1053 ( .A1(_02085__PTR132), .A2(_02085__PTR164), .ZN(_00574__PTR2) );
  OR2_X1 U1054 ( .A1(_00574__PTR0), .A2(_00574__PTR1), .ZN(_00575__PTR0) );
  OR2_X1 U1055 ( .A1(_00574__PTR2), .A2(_02085__PTR196), .ZN(_00575__PTR1) );
  OR2_X1 U1056 ( .A1(_00575__PTR0), .A2(_00575__PTR1), .ZN(_02087__PTR4) );
  OR2_X1 U1057 ( .A1(_02085__PTR3), .A2(_02085__PTR35), .ZN(_00576__PTR0) );
  OR2_X1 U1058 ( .A1(_02085__PTR67), .A2(_02085__PTR99), .ZN(_00576__PTR1) );
  OR2_X1 U1059 ( .A1(_02085__PTR131), .A2(_02085__PTR163), .ZN(_00576__PTR2) );
  OR2_X1 U1060 ( .A1(_00576__PTR0), .A2(_00576__PTR1), .ZN(_00577__PTR0) );
  OR2_X1 U1061 ( .A1(_00576__PTR2), .A2(_02085__PTR195), .ZN(_00577__PTR1) );
  OR2_X1 U1062 ( .A1(_00577__PTR0), .A2(_00577__PTR1), .ZN(_02087__PTR3) );
  OR2_X1 U1063 ( .A1(_02085__PTR2), .A2(_02085__PTR34), .ZN(_00578__PTR0) );
  OR2_X1 U1064 ( .A1(_02085__PTR66), .A2(_02085__PTR98), .ZN(_00578__PTR1) );
  OR2_X1 U1065 ( .A1(_02085__PTR130), .A2(_02085__PTR162), .ZN(_00578__PTR2) );
  OR2_X1 U1066 ( .A1(_00578__PTR0), .A2(_00578__PTR1), .ZN(_00579__PTR0) );
  OR2_X1 U1067 ( .A1(_00578__PTR2), .A2(_02085__PTR194), .ZN(_00579__PTR1) );
  OR2_X1 U1068 ( .A1(_00579__PTR0), .A2(_00579__PTR1), .ZN(_02087__PTR2) );
  OR2_X1 U1069 ( .A1(_02085__PTR1), .A2(_02085__PTR33), .ZN(_00580__PTR0) );
  OR2_X1 U1070 ( .A1(_02085__PTR65), .A2(_02085__PTR97), .ZN(_00580__PTR1) );
  OR2_X1 U1071 ( .A1(_02085__PTR129), .A2(_02085__PTR161), .ZN(_00580__PTR2) );
  OR2_X1 U1072 ( .A1(_00580__PTR0), .A2(_00580__PTR1), .ZN(_00581__PTR0) );
  OR2_X1 U1073 ( .A1(_00580__PTR2), .A2(_02085__PTR193), .ZN(_00581__PTR1) );
  OR2_X1 U1074 ( .A1(_00581__PTR0), .A2(_00581__PTR1), .ZN(_02087__PTR1) );
  OR2_X1 U1075 ( .A1(_02085__PTR0), .A2(_02085__PTR32), .ZN(_00582__PTR0) );
  OR2_X1 U1076 ( .A1(_02085__PTR64), .A2(_02085__PTR96), .ZN(_00582__PTR1) );
  OR2_X1 U1077 ( .A1(_02085__PTR128), .A2(_02085__PTR160), .ZN(_00582__PTR2) );
  OR2_X1 U1078 ( .A1(_00582__PTR0), .A2(_00582__PTR1), .ZN(_00583__PTR0) );
  OR2_X1 U1079 ( .A1(_00582__PTR2), .A2(_02085__PTR192), .ZN(_00583__PTR1) );
  OR2_X1 U1080 ( .A1(_00583__PTR0), .A2(_00583__PTR1), .ZN(_02087__PTR0) );
  OR2_X1 U1081 ( .A1(_02086__PTR0), .A2(_02086__PTR1), .ZN(_00481__PTR0) );
  OR2_X1 U1082 ( .A1(_01855__PTR0), .A2(_01855__PTR1), .ZN(_00469__PTR0) );
  OR2_X1 U1083 ( .A1(_02086__PTR4), .A2(_01855__PTR2), .ZN(_01859__PTR2) );
  OR2_X1 U1084 ( .A1(_00481__PTR0), .A2(_00469__PTR0), .ZN(_00584__PTR0) );
  OR2_X1 U1085 ( .A1(_01859__PTR2), .A2(_01855__PTR3), .ZN(_00469__PTR1) );
  OR2_X1 U1086 ( .A1(_00584__PTR0), .A2(_00469__PTR1), .ZN(_02920_) );
  OR2_X1 U1087 ( .A1(_02093__PTR0), .A2(_02093__PTR32), .ZN(_00585_) );
  OR2_X1 U1088 ( .A1(_00585_), .A2(_02093__PTR64), .ZN(_02095__PTR0) );
  OR2_X1 U1089 ( .A1(_02093__PTR1), .A2(_02093__PTR33), .ZN(_00586_) );
  OR2_X1 U1090 ( .A1(_00586_), .A2(_02093__PTR65), .ZN(_02095__PTR1) );
  OR2_X1 U1091 ( .A1(_02093__PTR2), .A2(_02093__PTR34), .ZN(_00587_) );
  OR2_X1 U1092 ( .A1(_00587_), .A2(_02093__PTR66), .ZN(_02095__PTR2) );
  OR2_X1 U1093 ( .A1(_02093__PTR3), .A2(_02093__PTR35), .ZN(_00588_) );
  OR2_X1 U1094 ( .A1(_00588_), .A2(_02093__PTR67), .ZN(_02095__PTR3) );
  OR2_X1 U1095 ( .A1(_02093__PTR4), .A2(_02093__PTR36), .ZN(_00589_) );
  OR2_X1 U1096 ( .A1(_00589_), .A2(_02093__PTR68), .ZN(_02095__PTR4) );
  OR2_X1 U1097 ( .A1(_02093__PTR5), .A2(_02093__PTR37), .ZN(_00590_) );
  OR2_X1 U1098 ( .A1(_00590_), .A2(_02093__PTR69), .ZN(_02095__PTR5) );
  OR2_X1 U1099 ( .A1(_02093__PTR6), .A2(_02093__PTR38), .ZN(_00591_) );
  OR2_X1 U1100 ( .A1(_00591_), .A2(_02093__PTR70), .ZN(_02095__PTR6) );
  OR2_X1 U1101 ( .A1(_02093__PTR7), .A2(_02093__PTR39), .ZN(_00592_) );
  OR2_X1 U1102 ( .A1(_00592_), .A2(_02093__PTR71), .ZN(_02095__PTR7) );
  OR2_X1 U1103 ( .A1(_02093__PTR8), .A2(_02093__PTR40), .ZN(_00593_) );
  OR2_X1 U1104 ( .A1(_00593_), .A2(_02093__PTR72), .ZN(_02095__PTR8) );
  OR2_X1 U1105 ( .A1(_02093__PTR9), .A2(_02093__PTR41), .ZN(_00594_) );
  OR2_X1 U1106 ( .A1(_00594_), .A2(_02093__PTR73), .ZN(_02095__PTR9) );
  OR2_X1 U1107 ( .A1(_02093__PTR10), .A2(_02093__PTR42), .ZN(_00595_) );
  OR2_X1 U1108 ( .A1(_00595_), .A2(_02093__PTR74), .ZN(_02095__PTR10) );
  OR2_X1 U1109 ( .A1(_02093__PTR11), .A2(_02093__PTR43), .ZN(_00596_) );
  OR2_X1 U1110 ( .A1(_00596_), .A2(_02093__PTR75), .ZN(_02095__PTR11) );
  OR2_X1 U1111 ( .A1(_02093__PTR12), .A2(_02093__PTR44), .ZN(_00597_) );
  OR2_X1 U1112 ( .A1(_00597_), .A2(_02093__PTR76), .ZN(_02095__PTR12) );
  OR2_X1 U1113 ( .A1(_02093__PTR13), .A2(_02093__PTR45), .ZN(_00598_) );
  OR2_X1 U1114 ( .A1(_00598_), .A2(_02093__PTR77), .ZN(_02095__PTR13) );
  OR2_X1 U1115 ( .A1(_02093__PTR14), .A2(_02093__PTR46), .ZN(_00599_) );
  OR2_X1 U1116 ( .A1(_00599_), .A2(_02093__PTR78), .ZN(_02095__PTR14) );
  OR2_X1 U1117 ( .A1(_02093__PTR15), .A2(_02093__PTR47), .ZN(_00600_) );
  OR2_X1 U1118 ( .A1(_00600_), .A2(_02093__PTR79), .ZN(_02095__PTR15) );
  OR2_X1 U1119 ( .A1(_02093__PTR16), .A2(_02093__PTR48), .ZN(_00601_) );
  OR2_X1 U1120 ( .A1(_00601_), .A2(_02093__PTR80), .ZN(_02095__PTR16) );
  OR2_X1 U1121 ( .A1(_02093__PTR17), .A2(_02093__PTR49), .ZN(_00602_) );
  OR2_X1 U1122 ( .A1(_00602_), .A2(_02093__PTR81), .ZN(_02095__PTR17) );
  OR2_X1 U1123 ( .A1(_02093__PTR18), .A2(_02093__PTR50), .ZN(_00603_) );
  OR2_X1 U1124 ( .A1(_00603_), .A2(_02093__PTR82), .ZN(_02095__PTR18) );
  OR2_X1 U1125 ( .A1(_02093__PTR19), .A2(_02093__PTR51), .ZN(_00604_) );
  OR2_X1 U1126 ( .A1(_00604_), .A2(_02093__PTR83), .ZN(_02095__PTR19) );
  OR2_X1 U1127 ( .A1(_02093__PTR20), .A2(_02093__PTR52), .ZN(_00605_) );
  OR2_X1 U1128 ( .A1(_00605_), .A2(_02093__PTR84), .ZN(_02095__PTR20) );
  OR2_X1 U1129 ( .A1(_02093__PTR21), .A2(_02093__PTR53), .ZN(_00606_) );
  OR2_X1 U1130 ( .A1(_00606_), .A2(_02093__PTR85), .ZN(_02095__PTR21) );
  OR2_X1 U1131 ( .A1(_02093__PTR22), .A2(_02093__PTR54), .ZN(_00607_) );
  OR2_X1 U1132 ( .A1(_00607_), .A2(_02093__PTR86), .ZN(_02095__PTR22) );
  OR2_X1 U1133 ( .A1(_02093__PTR23), .A2(_02093__PTR55), .ZN(_00608_) );
  OR2_X1 U1134 ( .A1(_00608_), .A2(_02093__PTR87), .ZN(_02095__PTR23) );
  OR2_X1 U1135 ( .A1(_02093__PTR24), .A2(_02093__PTR56), .ZN(_00609_) );
  OR2_X1 U1136 ( .A1(_00609_), .A2(_02093__PTR88), .ZN(_02095__PTR24) );
  OR2_X1 U1137 ( .A1(_02093__PTR25), .A2(_02093__PTR57), .ZN(_00610_) );
  OR2_X1 U1138 ( .A1(_00610_), .A2(_02093__PTR89), .ZN(_02095__PTR25) );
  OR2_X1 U1139 ( .A1(_02093__PTR26), .A2(_02093__PTR58), .ZN(_00611_) );
  OR2_X1 U1140 ( .A1(_00611_), .A2(_02093__PTR90), .ZN(_02095__PTR26) );
  OR2_X1 U1141 ( .A1(_02093__PTR27), .A2(_02093__PTR59), .ZN(_00612_) );
  OR2_X1 U1142 ( .A1(_00612_), .A2(_02093__PTR91), .ZN(_02095__PTR27) );
  OR2_X1 U1143 ( .A1(_02093__PTR28), .A2(_02093__PTR60), .ZN(_00613_) );
  OR2_X1 U1144 ( .A1(_00613_), .A2(_02093__PTR92), .ZN(_02095__PTR28) );
  OR2_X1 U1145 ( .A1(_02093__PTR29), .A2(_02093__PTR61), .ZN(_00614_) );
  OR2_X1 U1146 ( .A1(_00614_), .A2(_02093__PTR93), .ZN(_02095__PTR29) );
  OR2_X1 U1147 ( .A1(_02093__PTR30), .A2(_02093__PTR62), .ZN(_00615_) );
  OR2_X1 U1148 ( .A1(_00615_), .A2(_02093__PTR94), .ZN(_02095__PTR30) );
  OR2_X1 U1149 ( .A1(_02093__PTR31), .A2(_02093__PTR63), .ZN(_00616_) );
  OR2_X1 U1150 ( .A1(_00616_), .A2(_02093__PTR95), .ZN(_02095__PTR31) );
  OR2_X1 U1151 ( .A1(_02094__PTR0), .A2(_01855__PTR2), .ZN(_00617_) );
  OR2_X1 U1152 ( .A1(_00617_), .A2(_01855__PTR3), .ZN(_02922_) );
  OR2_X1 U1153 ( .A1(_02752_), .A2(_02753_), .ZN(_01770__PTR2) );
  OR2_X1 U1154 ( .A1(_02119__PTR3), .A2(_02119__PTR7), .ZN(_02122__PTR3) );
  OR2_X1 U1155 ( .A1(_02119__PTR2), .A2(_02119__PTR6), .ZN(_02122__PTR2) );
  OR2_X1 U1156 ( .A1(_02119__PTR1), .A2(_02119__PTR5), .ZN(_02122__PTR1) );
  OR2_X1 U1157 ( .A1(_02119__PTR0), .A2(_02119__PTR4), .ZN(_02122__PTR0) );
  OR2_X1 U1158 ( .A1(_02120__PTR0), .A2(_01863__PTR2), .ZN(_02928_) );
  AND2_X1 U1159 ( .A1(_02718__PTR4), .A2(_02720__PTR5), .ZN(_00618__PTR2) );
  AND2_X1 U1160 ( .A1(_00618__PTR0), .A2(_02719__PTR3), .ZN(_00619_) );
  AND2_X1 U1161 ( .A1(_00619_), .A2(_00618__PTR2), .ZN(_02731_) );
  OR2_X1 U1162 ( .A1(_02730_), .A2(_02731_), .ZN(_02006_) );
  OR2_X1 U1163 ( .A1(_02727_), .A2(_02728_), .ZN(_01853__PTR2) );
  AND2_X1 U1164 ( .A1(_02717__PTR0), .A2(_02718__PTR1), .ZN(_00620__PTR0) );
  AND2_X1 U1165 ( .A1(_00620__PTR0), .A2(_00620__PTR1), .ZN(_00621_) );
  AND2_X1 U1166 ( .A1(_00621_), .A2(_00618__PTR2), .ZN(_02728_) );
  OR2_X1 U1167 ( .A1(_02721_), .A2(_02722_), .ZN(_01853__PTR3) );
  AND2_X1 U1168 ( .A1(_02717__PTR0), .A2(_02717__PTR1), .ZN(_00622__PTR0) );
  AND2_X1 U1169 ( .A1(_00622__PTR0), .A2(_02719__PTR3), .ZN(_00623_) );
  AND2_X1 U1170 ( .A1(_00623_), .A2(_00618__PTR2), .ZN(_02722_) );
  OR2_X1 U1171 ( .A1(_02412__PTR8), .A2(_02412__PTR12), .ZN(_00624__PTR1) );
  OR2_X1 U1172 ( .A1(_02412__PTR4), .A2(_00624__PTR1), .ZN(_02415__PTR0) );
  OR2_X1 U1173 ( .A1(_02412__PTR9), .A2(_02412__PTR13), .ZN(_00625__PTR1) );
  OR2_X1 U1174 ( .A1(_02412__PTR5), .A2(_00625__PTR1), .ZN(_02415__PTR1) );
  OR2_X1 U1175 ( .A1(_02412__PTR10), .A2(_02412__PTR14), .ZN(_00626__PTR1) );
  OR2_X1 U1176 ( .A1(_02412__PTR6), .A2(_00626__PTR1), .ZN(_02415__PTR2) );
  OR2_X1 U1177 ( .A1(_02412__PTR11), .A2(_02412__PTR15), .ZN(_02415__PTR3) );
  OR2_X1 U1178 ( .A1(_02413__PTR0), .A2(_02413__PTR1), .ZN(_00627__PTR0) );
  OR2_X1 U1179 ( .A1(_02413__PTR2), .A2(_02413__PTR3), .ZN(_00627__PTR1) );
  OR2_X1 U1180 ( .A1(_00627__PTR0), .A2(_00627__PTR1), .ZN(_03174_) );
  OR2_X1 U1181 ( .A1(_02404__PTR0), .A2(_02404__PTR32), .ZN(_00628_) );
  OR2_X1 U1182 ( .A1(_00628_), .A2(_02404__PTR64), .ZN(_02406__PTR0) );
  OR2_X1 U1183 ( .A1(_02404__PTR1), .A2(_02404__PTR33), .ZN(_00629_) );
  OR2_X1 U1184 ( .A1(_00629_), .A2(_02404__PTR65), .ZN(_02406__PTR1) );
  OR2_X1 U1185 ( .A1(_02404__PTR2), .A2(_02404__PTR34), .ZN(_00630_) );
  OR2_X1 U1186 ( .A1(_00630_), .A2(_02404__PTR66), .ZN(_02406__PTR2) );
  OR2_X1 U1187 ( .A1(_02404__PTR3), .A2(_02404__PTR35), .ZN(_00631_) );
  OR2_X1 U1188 ( .A1(_00631_), .A2(_02404__PTR67), .ZN(_02406__PTR3) );
  OR2_X1 U1189 ( .A1(_02404__PTR4), .A2(_02404__PTR36), .ZN(_00632_) );
  OR2_X1 U1190 ( .A1(_00632_), .A2(_02404__PTR68), .ZN(_02406__PTR4) );
  OR2_X1 U1191 ( .A1(_02404__PTR5), .A2(_02404__PTR37), .ZN(_00633_) );
  OR2_X1 U1192 ( .A1(_00633_), .A2(_02404__PTR69), .ZN(_02406__PTR5) );
  OR2_X1 U1193 ( .A1(_02404__PTR6), .A2(_02404__PTR38), .ZN(_00634_) );
  OR2_X1 U1194 ( .A1(_00634_), .A2(_02404__PTR70), .ZN(_02406__PTR6) );
  OR2_X1 U1195 ( .A1(_02404__PTR7), .A2(_02404__PTR39), .ZN(_00635_) );
  OR2_X1 U1196 ( .A1(_00635_), .A2(_02404__PTR71), .ZN(_02406__PTR7) );
  OR2_X1 U1197 ( .A1(_02404__PTR8), .A2(_02404__PTR40), .ZN(_00636_) );
  OR2_X1 U1198 ( .A1(_00636_), .A2(_02404__PTR72), .ZN(_02406__PTR8) );
  OR2_X1 U1199 ( .A1(_02404__PTR9), .A2(_02404__PTR41), .ZN(_00637_) );
  OR2_X1 U1200 ( .A1(_00637_), .A2(_02404__PTR73), .ZN(_02406__PTR9) );
  OR2_X1 U1201 ( .A1(_02404__PTR10), .A2(_02404__PTR42), .ZN(_00638_) );
  OR2_X1 U1202 ( .A1(_00638_), .A2(_02404__PTR74), .ZN(_02406__PTR10) );
  OR2_X1 U1203 ( .A1(_02404__PTR11), .A2(_02404__PTR43), .ZN(_00639_) );
  OR2_X1 U1204 ( .A1(_00639_), .A2(_02404__PTR75), .ZN(_02406__PTR11) );
  OR2_X1 U1205 ( .A1(_02404__PTR12), .A2(_02404__PTR44), .ZN(_00640_) );
  OR2_X1 U1206 ( .A1(_00640_), .A2(_02404__PTR76), .ZN(_02406__PTR12) );
  OR2_X1 U1207 ( .A1(_02404__PTR13), .A2(_02404__PTR45), .ZN(_00641_) );
  OR2_X1 U1208 ( .A1(_00641_), .A2(_02404__PTR77), .ZN(_02406__PTR13) );
  OR2_X1 U1209 ( .A1(_02404__PTR14), .A2(_02404__PTR46), .ZN(_00642_) );
  OR2_X1 U1210 ( .A1(_00642_), .A2(_02404__PTR78), .ZN(_02406__PTR14) );
  OR2_X1 U1211 ( .A1(_02404__PTR15), .A2(_02404__PTR47), .ZN(_00643_) );
  OR2_X1 U1212 ( .A1(_00643_), .A2(_02404__PTR79), .ZN(_02406__PTR15) );
  OR2_X1 U1213 ( .A1(_02404__PTR16), .A2(_02404__PTR48), .ZN(_00644_) );
  OR2_X1 U1214 ( .A1(_00644_), .A2(_02404__PTR80), .ZN(_02406__PTR16) );
  OR2_X1 U1215 ( .A1(_02404__PTR17), .A2(_02404__PTR49), .ZN(_00645_) );
  OR2_X1 U1216 ( .A1(_00645_), .A2(_02404__PTR81), .ZN(_02406__PTR17) );
  OR2_X1 U1217 ( .A1(_02404__PTR18), .A2(_02404__PTR50), .ZN(_00646_) );
  OR2_X1 U1218 ( .A1(_00646_), .A2(_02404__PTR82), .ZN(_02406__PTR18) );
  OR2_X1 U1219 ( .A1(_02404__PTR19), .A2(_02404__PTR51), .ZN(_00647_) );
  OR2_X1 U1220 ( .A1(_00647_), .A2(_02404__PTR83), .ZN(_02406__PTR19) );
  OR2_X1 U1221 ( .A1(_02404__PTR20), .A2(_02404__PTR52), .ZN(_00648_) );
  OR2_X1 U1222 ( .A1(_00648_), .A2(_02404__PTR84), .ZN(_02406__PTR20) );
  OR2_X1 U1223 ( .A1(_02404__PTR21), .A2(_02404__PTR53), .ZN(_00649_) );
  OR2_X1 U1224 ( .A1(_00649_), .A2(_02404__PTR85), .ZN(_02406__PTR21) );
  OR2_X1 U1225 ( .A1(_02404__PTR22), .A2(_02404__PTR54), .ZN(_00650_) );
  OR2_X1 U1226 ( .A1(_00650_), .A2(_02404__PTR86), .ZN(_02406__PTR22) );
  OR2_X1 U1227 ( .A1(_02404__PTR23), .A2(_02404__PTR55), .ZN(_00651_) );
  OR2_X1 U1228 ( .A1(_00651_), .A2(_02404__PTR87), .ZN(_02406__PTR23) );
  OR2_X1 U1229 ( .A1(_02404__PTR24), .A2(_02404__PTR56), .ZN(_00652_) );
  OR2_X1 U1230 ( .A1(_00652_), .A2(_02404__PTR88), .ZN(_02406__PTR24) );
  OR2_X1 U1231 ( .A1(_02404__PTR25), .A2(_02404__PTR57), .ZN(_00653_) );
  OR2_X1 U1232 ( .A1(_00653_), .A2(_02404__PTR89), .ZN(_02406__PTR25) );
  OR2_X1 U1233 ( .A1(_02404__PTR26), .A2(_02404__PTR58), .ZN(_00654_) );
  OR2_X1 U1234 ( .A1(_00654_), .A2(_02404__PTR90), .ZN(_02406__PTR26) );
  OR2_X1 U1235 ( .A1(_02404__PTR27), .A2(_02404__PTR59), .ZN(_00655_) );
  OR2_X1 U1236 ( .A1(_00655_), .A2(_02404__PTR91), .ZN(_02406__PTR27) );
  OR2_X1 U1237 ( .A1(_02404__PTR28), .A2(_02404__PTR60), .ZN(_00656_) );
  OR2_X1 U1238 ( .A1(_00656_), .A2(_02404__PTR92), .ZN(_02406__PTR28) );
  OR2_X1 U1239 ( .A1(_02404__PTR29), .A2(_02404__PTR61), .ZN(_00657_) );
  OR2_X1 U1240 ( .A1(_00657_), .A2(_02404__PTR93), .ZN(_02406__PTR29) );
  OR2_X1 U1241 ( .A1(_02404__PTR30), .A2(_02404__PTR62), .ZN(_00658_) );
  OR2_X1 U1242 ( .A1(_00658_), .A2(_02404__PTR94), .ZN(_02406__PTR30) );
  OR2_X1 U1243 ( .A1(_02404__PTR31), .A2(_02404__PTR63), .ZN(_00659_) );
  OR2_X1 U1244 ( .A1(_00659_), .A2(_02404__PTR95), .ZN(_02406__PTR31) );
  OR2_X1 U1245 ( .A1(_02405__PTR0), .A2(_02156__PTR0), .ZN(_00660_) );
  OR2_X1 U1246 ( .A1(_00660_), .A2(_02156__PTR2), .ZN(_03172_) );
  OR2_X1 U1247 ( .A1(_02401__PTR0), .A2(_02401__PTR16), .ZN(_00661_) );
  OR2_X1 U1248 ( .A1(_00661_), .A2(_02401__PTR32), .ZN(_02402__PTR0) );
  OR2_X1 U1249 ( .A1(_02401__PTR1), .A2(_02401__PTR17), .ZN(_00662_) );
  OR2_X1 U1250 ( .A1(_00662_), .A2(_02401__PTR33), .ZN(_02402__PTR1) );
  OR2_X1 U1251 ( .A1(_02401__PTR2), .A2(_02401__PTR18), .ZN(_00663_) );
  OR2_X1 U1252 ( .A1(_00663_), .A2(_02401__PTR34), .ZN(_02402__PTR2) );
  OR2_X1 U1253 ( .A1(_02401__PTR3), .A2(_02401__PTR19), .ZN(_00664_) );
  OR2_X1 U1254 ( .A1(_00664_), .A2(_02401__PTR35), .ZN(_02402__PTR3) );
  OR2_X1 U1255 ( .A1(_02401__PTR4), .A2(_02401__PTR20), .ZN(_00665_) );
  OR2_X1 U1256 ( .A1(_00665_), .A2(_02401__PTR36), .ZN(_02402__PTR4) );
  OR2_X1 U1257 ( .A1(_02401__PTR5), .A2(_02401__PTR21), .ZN(_00666_) );
  OR2_X1 U1258 ( .A1(_00666_), .A2(_02401__PTR37), .ZN(_02402__PTR5) );
  OR2_X1 U1259 ( .A1(_02401__PTR6), .A2(_02401__PTR22), .ZN(_00667_) );
  OR2_X1 U1260 ( .A1(_00667_), .A2(_02401__PTR38), .ZN(_02402__PTR6) );
  OR2_X1 U1261 ( .A1(_02401__PTR7), .A2(_02401__PTR23), .ZN(_00668_) );
  OR2_X1 U1262 ( .A1(_00668_), .A2(_02401__PTR39), .ZN(_02402__PTR7) );
  OR2_X1 U1263 ( .A1(_02401__PTR8), .A2(_02401__PTR24), .ZN(_00669_) );
  OR2_X1 U1264 ( .A1(_00669_), .A2(_02401__PTR40), .ZN(_02402__PTR8) );
  OR2_X1 U1265 ( .A1(_02401__PTR9), .A2(_02401__PTR25), .ZN(_00670_) );
  OR2_X1 U1266 ( .A1(_00670_), .A2(_02401__PTR41), .ZN(_02402__PTR9) );
  OR2_X1 U1267 ( .A1(_02401__PTR10), .A2(_02401__PTR26), .ZN(_00671_) );
  OR2_X1 U1268 ( .A1(_00671_), .A2(_02401__PTR42), .ZN(_02402__PTR10) );
  OR2_X1 U1269 ( .A1(_02401__PTR11), .A2(_02401__PTR27), .ZN(_00672_) );
  OR2_X1 U1270 ( .A1(_00672_), .A2(_02401__PTR43), .ZN(_02402__PTR11) );
  OR2_X1 U1271 ( .A1(_02401__PTR12), .A2(_02401__PTR28), .ZN(_00673_) );
  OR2_X1 U1272 ( .A1(_00673_), .A2(_02401__PTR44), .ZN(_02402__PTR12) );
  OR2_X1 U1273 ( .A1(_02401__PTR13), .A2(_02401__PTR29), .ZN(_00674_) );
  OR2_X1 U1274 ( .A1(_00674_), .A2(_02401__PTR45), .ZN(_02402__PTR13) );
  OR2_X1 U1275 ( .A1(_02401__PTR14), .A2(_02401__PTR30), .ZN(_00675_) );
  OR2_X1 U1276 ( .A1(_00675_), .A2(_02401__PTR46), .ZN(_02402__PTR14) );
  OR2_X1 U1277 ( .A1(_02401__PTR15), .A2(_02401__PTR31), .ZN(_00676_) );
  OR2_X1 U1278 ( .A1(_00676_), .A2(_02401__PTR47), .ZN(_02402__PTR15) );
  OR2_X1 U1279 ( .A1(_02397__PTR0), .A2(_02397__PTR15), .ZN(_00678_) );
  OR2_X1 U1280 ( .A1(_00678_), .A2(_02397__PTR30), .ZN(_02399__PTR0) );
  OR2_X1 U1281 ( .A1(_02397__PTR1), .A2(_02397__PTR16), .ZN(_00679_) );
  OR2_X1 U1282 ( .A1(_00679_), .A2(_02397__PTR31), .ZN(_02399__PTR1) );
  OR2_X1 U1283 ( .A1(_02397__PTR2), .A2(_02397__PTR17), .ZN(_00680_) );
  OR2_X1 U1284 ( .A1(_00680_), .A2(_02397__PTR32), .ZN(_02399__PTR2) );
  OR2_X1 U1285 ( .A1(_02397__PTR3), .A2(_02397__PTR18), .ZN(_00681_) );
  OR2_X1 U1286 ( .A1(_00681_), .A2(_02397__PTR33), .ZN(_02399__PTR3) );
  OR2_X1 U1287 ( .A1(_02397__PTR4), .A2(_02397__PTR19), .ZN(_00682_) );
  OR2_X1 U1288 ( .A1(_00682_), .A2(_02397__PTR34), .ZN(_02399__PTR4) );
  OR2_X1 U1289 ( .A1(_02397__PTR5), .A2(_02397__PTR20), .ZN(_00683_) );
  OR2_X1 U1290 ( .A1(_00683_), .A2(_02397__PTR35), .ZN(_02399__PTR5) );
  OR2_X1 U1291 ( .A1(_02397__PTR6), .A2(_02397__PTR21), .ZN(_00684_) );
  OR2_X1 U1292 ( .A1(_00684_), .A2(_02397__PTR36), .ZN(_02399__PTR6) );
  OR2_X1 U1293 ( .A1(_02397__PTR7), .A2(_02397__PTR22), .ZN(_00685_) );
  OR2_X1 U1294 ( .A1(_00685_), .A2(_02397__PTR37), .ZN(_02399__PTR7) );
  OR2_X1 U1295 ( .A1(_02397__PTR8), .A2(_02397__PTR23), .ZN(_00686_) );
  OR2_X1 U1296 ( .A1(_00686_), .A2(_02397__PTR38), .ZN(_02399__PTR8) );
  OR2_X1 U1297 ( .A1(_02397__PTR9), .A2(_02397__PTR24), .ZN(_00687_) );
  OR2_X1 U1298 ( .A1(_00687_), .A2(_02397__PTR39), .ZN(_02399__PTR9) );
  OR2_X1 U1299 ( .A1(_02397__PTR10), .A2(_02397__PTR25), .ZN(_00688_) );
  OR2_X1 U1300 ( .A1(_00688_), .A2(_02397__PTR40), .ZN(_02399__PTR10) );
  OR2_X1 U1301 ( .A1(_02397__PTR11), .A2(_02397__PTR26), .ZN(_00689_) );
  OR2_X1 U1302 ( .A1(_00689_), .A2(_02397__PTR41), .ZN(_02399__PTR11) );
  OR2_X1 U1303 ( .A1(_02397__PTR12), .A2(_02397__PTR27), .ZN(_00690_) );
  OR2_X1 U1304 ( .A1(_00690_), .A2(_02397__PTR42), .ZN(_02399__PTR12) );
  OR2_X1 U1305 ( .A1(_02397__PTR13), .A2(_02397__PTR28), .ZN(_00691_) );
  OR2_X1 U1306 ( .A1(_00691_), .A2(_02397__PTR43), .ZN(_02399__PTR13) );
  OR2_X1 U1307 ( .A1(_02397__PTR14), .A2(_02397__PTR29), .ZN(_00692_) );
  OR2_X1 U1308 ( .A1(_00692_), .A2(_02397__PTR44), .ZN(_02399__PTR14) );
  OR2_X1 U1309 ( .A1(_02398__PTR0), .A2(_02156__PTR2), .ZN(_00677_) );
  OR2_X1 U1310 ( .A1(_00677_), .A2(_02379__PTR4), .ZN(_03171_) );
  OR2_X1 U1311 ( .A1(_02390__PTR0), .A2(_02390__PTR32), .ZN(_00693_) );
  OR2_X1 U1312 ( .A1(_00693_), .A2(_02390__PTR64), .ZN(_02392__PTR0) );
  OR2_X1 U1313 ( .A1(_02390__PTR1), .A2(_02390__PTR33), .ZN(_00694_) );
  OR2_X1 U1314 ( .A1(_00694_), .A2(_02390__PTR65), .ZN(_02392__PTR1) );
  OR2_X1 U1315 ( .A1(_02390__PTR2), .A2(_02390__PTR34), .ZN(_00695_) );
  OR2_X1 U1316 ( .A1(_00695_), .A2(_02390__PTR66), .ZN(_02392__PTR2) );
  OR2_X1 U1317 ( .A1(_02390__PTR3), .A2(_02390__PTR35), .ZN(_00696_) );
  OR2_X1 U1318 ( .A1(_00696_), .A2(_02390__PTR67), .ZN(_02392__PTR3) );
  OR2_X1 U1319 ( .A1(_02390__PTR4), .A2(_02390__PTR36), .ZN(_00697_) );
  OR2_X1 U1320 ( .A1(_00697_), .A2(_02390__PTR68), .ZN(_02392__PTR4) );
  OR2_X1 U1321 ( .A1(_02390__PTR5), .A2(_02390__PTR37), .ZN(_00698_) );
  OR2_X1 U1322 ( .A1(_00698_), .A2(_02390__PTR69), .ZN(_02392__PTR5) );
  OR2_X1 U1323 ( .A1(_02390__PTR6), .A2(_02390__PTR38), .ZN(_00699_) );
  OR2_X1 U1324 ( .A1(_00699_), .A2(_02390__PTR70), .ZN(_02392__PTR6) );
  OR2_X1 U1325 ( .A1(_02390__PTR7), .A2(_02390__PTR39), .ZN(_00700_) );
  OR2_X1 U1326 ( .A1(_00700_), .A2(_02390__PTR71), .ZN(_02392__PTR7) );
  OR2_X1 U1327 ( .A1(_02390__PTR8), .A2(_02390__PTR40), .ZN(_00701_) );
  OR2_X1 U1328 ( .A1(_00701_), .A2(_02390__PTR72), .ZN(_02392__PTR8) );
  OR2_X1 U1329 ( .A1(_02390__PTR9), .A2(_02390__PTR41), .ZN(_00702_) );
  OR2_X1 U1330 ( .A1(_00702_), .A2(_02390__PTR73), .ZN(_02392__PTR9) );
  OR2_X1 U1331 ( .A1(_02390__PTR10), .A2(_02390__PTR42), .ZN(_00703_) );
  OR2_X1 U1332 ( .A1(_00703_), .A2(_02390__PTR74), .ZN(_02392__PTR10) );
  OR2_X1 U1333 ( .A1(_02390__PTR11), .A2(_02390__PTR43), .ZN(_00704_) );
  OR2_X1 U1334 ( .A1(_00704_), .A2(_02390__PTR75), .ZN(_02392__PTR11) );
  OR2_X1 U1335 ( .A1(_02390__PTR12), .A2(_02390__PTR44), .ZN(_00705_) );
  OR2_X1 U1336 ( .A1(_00705_), .A2(_02390__PTR76), .ZN(_02392__PTR12) );
  OR2_X1 U1337 ( .A1(_02390__PTR13), .A2(_02390__PTR45), .ZN(_00706_) );
  OR2_X1 U1338 ( .A1(_00706_), .A2(_02390__PTR77), .ZN(_02392__PTR13) );
  OR2_X1 U1339 ( .A1(_02390__PTR14), .A2(_02390__PTR46), .ZN(_00707_) );
  OR2_X1 U1340 ( .A1(_00707_), .A2(_02390__PTR78), .ZN(_02392__PTR14) );
  OR2_X1 U1341 ( .A1(_02390__PTR15), .A2(_02390__PTR47), .ZN(_00708_) );
  OR2_X1 U1342 ( .A1(_00708_), .A2(_02390__PTR79), .ZN(_02392__PTR15) );
  OR2_X1 U1343 ( .A1(_02390__PTR16), .A2(_02390__PTR48), .ZN(_00709_) );
  OR2_X1 U1344 ( .A1(_00709_), .A2(_02390__PTR80), .ZN(_02392__PTR16) );
  OR2_X1 U1345 ( .A1(_02390__PTR17), .A2(_02390__PTR49), .ZN(_00710_) );
  OR2_X1 U1346 ( .A1(_00710_), .A2(_02390__PTR81), .ZN(_02392__PTR17) );
  OR2_X1 U1347 ( .A1(_02390__PTR18), .A2(_02390__PTR50), .ZN(_00711_) );
  OR2_X1 U1348 ( .A1(_00711_), .A2(_02390__PTR82), .ZN(_02392__PTR18) );
  OR2_X1 U1349 ( .A1(_02390__PTR19), .A2(_02390__PTR51), .ZN(_00712_) );
  OR2_X1 U1350 ( .A1(_00712_), .A2(_02390__PTR83), .ZN(_02392__PTR19) );
  OR2_X1 U1351 ( .A1(_02390__PTR20), .A2(_02390__PTR52), .ZN(_00713_) );
  OR2_X1 U1352 ( .A1(_00713_), .A2(_02390__PTR84), .ZN(_02392__PTR20) );
  OR2_X1 U1353 ( .A1(_02390__PTR21), .A2(_02390__PTR53), .ZN(_00714_) );
  OR2_X1 U1354 ( .A1(_00714_), .A2(_02390__PTR85), .ZN(_02392__PTR21) );
  OR2_X1 U1355 ( .A1(_02390__PTR22), .A2(_02390__PTR54), .ZN(_00715_) );
  OR2_X1 U1356 ( .A1(_00715_), .A2(_02390__PTR86), .ZN(_02392__PTR22) );
  OR2_X1 U1357 ( .A1(_02390__PTR23), .A2(_02390__PTR55), .ZN(_00716_) );
  OR2_X1 U1358 ( .A1(_00716_), .A2(_02390__PTR87), .ZN(_02392__PTR23) );
  OR2_X1 U1359 ( .A1(_02390__PTR24), .A2(_02390__PTR56), .ZN(_00717_) );
  OR2_X1 U1360 ( .A1(_00717_), .A2(_02390__PTR88), .ZN(_02392__PTR24) );
  OR2_X1 U1361 ( .A1(_02390__PTR25), .A2(_02390__PTR57), .ZN(_00718_) );
  OR2_X1 U1362 ( .A1(_00718_), .A2(_02390__PTR89), .ZN(_02392__PTR25) );
  OR2_X1 U1363 ( .A1(_02390__PTR26), .A2(_02390__PTR58), .ZN(_00719_) );
  OR2_X1 U1364 ( .A1(_00719_), .A2(_02390__PTR90), .ZN(_02392__PTR26) );
  OR2_X1 U1365 ( .A1(_02390__PTR27), .A2(_02390__PTR59), .ZN(_00720_) );
  OR2_X1 U1366 ( .A1(_00720_), .A2(_02390__PTR91), .ZN(_02392__PTR27) );
  OR2_X1 U1367 ( .A1(_02390__PTR28), .A2(_02390__PTR60), .ZN(_00721_) );
  OR2_X1 U1368 ( .A1(_00721_), .A2(_02390__PTR92), .ZN(_02392__PTR28) );
  OR2_X1 U1369 ( .A1(_02390__PTR29), .A2(_02390__PTR61), .ZN(_00722_) );
  OR2_X1 U1370 ( .A1(_00722_), .A2(_02390__PTR93), .ZN(_02392__PTR29) );
  OR2_X1 U1371 ( .A1(_02390__PTR30), .A2(_02390__PTR62), .ZN(_00723_) );
  OR2_X1 U1372 ( .A1(_00723_), .A2(_02390__PTR94), .ZN(_02392__PTR30) );
  OR2_X1 U1373 ( .A1(_02390__PTR31), .A2(_02390__PTR63), .ZN(_00724_) );
  OR2_X1 U1374 ( .A1(_00724_), .A2(_02390__PTR95), .ZN(_02392__PTR31) );
  OR2_X1 U1375 ( .A1(_02391__PTR0), .A2(_02391__PTR1), .ZN(_00725_) );
  OR2_X1 U1376 ( .A1(_00725_), .A2(_02391__PTR2), .ZN(_03169_) );
  OR2_X1 U1377 ( .A1(_02386__PTR0), .A2(_02386__PTR32), .ZN(_00726__PTR0) );
  OR2_X1 U1378 ( .A1(_02386__PTR64), .A2(_02386__PTR96), .ZN(_00726__PTR1) );
  OR2_X1 U1379 ( .A1(_00726__PTR0), .A2(_00726__PTR1), .ZN(_00727_) );
  OR2_X1 U1380 ( .A1(_00727_), .A2(_02386__PTR128), .ZN(_02388__PTR0) );
  OR2_X1 U1381 ( .A1(_02386__PTR1), .A2(_02386__PTR33), .ZN(_00728__PTR0) );
  OR2_X1 U1382 ( .A1(_02386__PTR65), .A2(_02386__PTR97), .ZN(_00728__PTR1) );
  OR2_X1 U1383 ( .A1(_00728__PTR0), .A2(_00728__PTR1), .ZN(_00729_) );
  OR2_X1 U1384 ( .A1(_00729_), .A2(_02386__PTR129), .ZN(_02388__PTR1) );
  OR2_X1 U1385 ( .A1(_02386__PTR2), .A2(_02386__PTR34), .ZN(_00730__PTR0) );
  OR2_X1 U1386 ( .A1(_02386__PTR66), .A2(_02386__PTR98), .ZN(_00730__PTR1) );
  OR2_X1 U1387 ( .A1(_00730__PTR0), .A2(_00730__PTR1), .ZN(_00731_) );
  OR2_X1 U1388 ( .A1(_00731_), .A2(_02386__PTR130), .ZN(_02388__PTR2) );
  OR2_X1 U1389 ( .A1(_02386__PTR3), .A2(_02386__PTR35), .ZN(_00732__PTR0) );
  OR2_X1 U1390 ( .A1(_02386__PTR67), .A2(_02386__PTR99), .ZN(_00732__PTR1) );
  OR2_X1 U1391 ( .A1(_00732__PTR0), .A2(_00732__PTR1), .ZN(_00733_) );
  OR2_X1 U1392 ( .A1(_00733_), .A2(_02386__PTR131), .ZN(_02388__PTR3) );
  OR2_X1 U1393 ( .A1(_02386__PTR4), .A2(_02386__PTR36), .ZN(_00734__PTR0) );
  OR2_X1 U1394 ( .A1(_02386__PTR68), .A2(_02386__PTR100), .ZN(_00734__PTR1) );
  OR2_X1 U1395 ( .A1(_00734__PTR0), .A2(_00734__PTR1), .ZN(_00735_) );
  OR2_X1 U1396 ( .A1(_00735_), .A2(_02386__PTR132), .ZN(_02388__PTR4) );
  OR2_X1 U1397 ( .A1(_02386__PTR5), .A2(_02386__PTR37), .ZN(_00736__PTR0) );
  OR2_X1 U1398 ( .A1(_02386__PTR69), .A2(_02386__PTR101), .ZN(_00736__PTR1) );
  OR2_X1 U1399 ( .A1(_00736__PTR0), .A2(_00736__PTR1), .ZN(_00737_) );
  OR2_X1 U1400 ( .A1(_00737_), .A2(_02386__PTR133), .ZN(_02388__PTR5) );
  OR2_X1 U1401 ( .A1(_02386__PTR6), .A2(_02386__PTR38), .ZN(_00738__PTR0) );
  OR2_X1 U1402 ( .A1(_02386__PTR70), .A2(_02386__PTR102), .ZN(_00738__PTR1) );
  OR2_X1 U1403 ( .A1(_00738__PTR0), .A2(_00738__PTR1), .ZN(_00739_) );
  OR2_X1 U1404 ( .A1(_00739_), .A2(_02386__PTR134), .ZN(_02388__PTR6) );
  OR2_X1 U1405 ( .A1(_02386__PTR7), .A2(_02386__PTR39), .ZN(_00740__PTR0) );
  OR2_X1 U1406 ( .A1(_02386__PTR71), .A2(_02386__PTR103), .ZN(_00740__PTR1) );
  OR2_X1 U1407 ( .A1(_00740__PTR0), .A2(_00740__PTR1), .ZN(_00741_) );
  OR2_X1 U1408 ( .A1(_00741_), .A2(_02386__PTR135), .ZN(_02388__PTR7) );
  OR2_X1 U1409 ( .A1(_02386__PTR8), .A2(_02386__PTR40), .ZN(_00742__PTR0) );
  OR2_X1 U1410 ( .A1(_02386__PTR72), .A2(_02386__PTR104), .ZN(_00742__PTR1) );
  OR2_X1 U1411 ( .A1(_00742__PTR0), .A2(_00742__PTR1), .ZN(_00743_) );
  OR2_X1 U1412 ( .A1(_00743_), .A2(_02386__PTR136), .ZN(_02388__PTR8) );
  OR2_X1 U1413 ( .A1(_02386__PTR9), .A2(_02386__PTR41), .ZN(_00744__PTR0) );
  OR2_X1 U1414 ( .A1(_02386__PTR73), .A2(_02386__PTR105), .ZN(_00744__PTR1) );
  OR2_X1 U1415 ( .A1(_00744__PTR0), .A2(_00744__PTR1), .ZN(_00745_) );
  OR2_X1 U1416 ( .A1(_00745_), .A2(_02386__PTR137), .ZN(_02388__PTR9) );
  OR2_X1 U1417 ( .A1(_02386__PTR10), .A2(_02386__PTR42), .ZN(_00746__PTR0) );
  OR2_X1 U1418 ( .A1(_02386__PTR74), .A2(_02386__PTR106), .ZN(_00746__PTR1) );
  OR2_X1 U1419 ( .A1(_00746__PTR0), .A2(_00746__PTR1), .ZN(_00747_) );
  OR2_X1 U1420 ( .A1(_00747_), .A2(_02386__PTR138), .ZN(_02388__PTR10) );
  OR2_X1 U1421 ( .A1(_02386__PTR11), .A2(_02386__PTR43), .ZN(_00748__PTR0) );
  OR2_X1 U1422 ( .A1(_02386__PTR75), .A2(_02386__PTR107), .ZN(_00748__PTR1) );
  OR2_X1 U1423 ( .A1(_00748__PTR0), .A2(_00748__PTR1), .ZN(_00749_) );
  OR2_X1 U1424 ( .A1(_00749_), .A2(_02386__PTR139), .ZN(_02388__PTR11) );
  OR2_X1 U1425 ( .A1(_02386__PTR12), .A2(_02386__PTR44), .ZN(_00750__PTR0) );
  OR2_X1 U1426 ( .A1(_02386__PTR76), .A2(_02386__PTR108), .ZN(_00750__PTR1) );
  OR2_X1 U1427 ( .A1(_00750__PTR0), .A2(_00750__PTR1), .ZN(_00751_) );
  OR2_X1 U1428 ( .A1(_00751_), .A2(_02386__PTR140), .ZN(_02388__PTR12) );
  OR2_X1 U1429 ( .A1(_02386__PTR13), .A2(_02386__PTR45), .ZN(_00752__PTR0) );
  OR2_X1 U1430 ( .A1(_02386__PTR77), .A2(_02386__PTR109), .ZN(_00752__PTR1) );
  OR2_X1 U1431 ( .A1(_00752__PTR0), .A2(_00752__PTR1), .ZN(_00753_) );
  OR2_X1 U1432 ( .A1(_00753_), .A2(_02386__PTR141), .ZN(_02388__PTR13) );
  OR2_X1 U1433 ( .A1(_02386__PTR14), .A2(_02386__PTR46), .ZN(_00754__PTR0) );
  OR2_X1 U1434 ( .A1(_02386__PTR78), .A2(_02386__PTR110), .ZN(_00754__PTR1) );
  OR2_X1 U1435 ( .A1(_00754__PTR0), .A2(_00754__PTR1), .ZN(_00755_) );
  OR2_X1 U1436 ( .A1(_00755_), .A2(_02386__PTR142), .ZN(_02388__PTR14) );
  OR2_X1 U1437 ( .A1(_02386__PTR15), .A2(_02386__PTR47), .ZN(_00756__PTR0) );
  OR2_X1 U1438 ( .A1(_02386__PTR79), .A2(_02386__PTR111), .ZN(_00756__PTR1) );
  OR2_X1 U1439 ( .A1(_00756__PTR0), .A2(_00756__PTR1), .ZN(_00757_) );
  OR2_X1 U1440 ( .A1(_00757_), .A2(_02386__PTR143), .ZN(_02388__PTR15) );
  OR2_X1 U1441 ( .A1(_02386__PTR16), .A2(_02386__PTR48), .ZN(_00758__PTR0) );
  OR2_X1 U1442 ( .A1(_02386__PTR80), .A2(_02386__PTR112), .ZN(_00758__PTR1) );
  OR2_X1 U1443 ( .A1(_00758__PTR0), .A2(_00758__PTR1), .ZN(_00759_) );
  OR2_X1 U1444 ( .A1(_00759_), .A2(_02386__PTR144), .ZN(_02388__PTR16) );
  OR2_X1 U1445 ( .A1(_02386__PTR17), .A2(_02386__PTR49), .ZN(_00760__PTR0) );
  OR2_X1 U1446 ( .A1(_02386__PTR81), .A2(_02386__PTR113), .ZN(_00760__PTR1) );
  OR2_X1 U1447 ( .A1(_00760__PTR0), .A2(_00760__PTR1), .ZN(_00761_) );
  OR2_X1 U1448 ( .A1(_00761_), .A2(_02386__PTR145), .ZN(_02388__PTR17) );
  OR2_X1 U1449 ( .A1(_02386__PTR18), .A2(_02386__PTR50), .ZN(_00762__PTR0) );
  OR2_X1 U1450 ( .A1(_02386__PTR82), .A2(_02386__PTR114), .ZN(_00762__PTR1) );
  OR2_X1 U1451 ( .A1(_00762__PTR0), .A2(_00762__PTR1), .ZN(_00763_) );
  OR2_X1 U1452 ( .A1(_00763_), .A2(_02386__PTR146), .ZN(_02388__PTR18) );
  OR2_X1 U1453 ( .A1(_02386__PTR19), .A2(_02386__PTR51), .ZN(_00764__PTR0) );
  OR2_X1 U1454 ( .A1(_02386__PTR83), .A2(_02386__PTR115), .ZN(_00764__PTR1) );
  OR2_X1 U1455 ( .A1(_00764__PTR0), .A2(_00764__PTR1), .ZN(_00765_) );
  OR2_X1 U1456 ( .A1(_00765_), .A2(_02386__PTR147), .ZN(_02388__PTR19) );
  OR2_X1 U1457 ( .A1(_02386__PTR20), .A2(_02386__PTR52), .ZN(_00766__PTR0) );
  OR2_X1 U1458 ( .A1(_02386__PTR84), .A2(_02386__PTR116), .ZN(_00766__PTR1) );
  OR2_X1 U1459 ( .A1(_00766__PTR0), .A2(_00766__PTR1), .ZN(_00767_) );
  OR2_X1 U1460 ( .A1(_00767_), .A2(_02386__PTR148), .ZN(_02388__PTR20) );
  OR2_X1 U1461 ( .A1(_02386__PTR21), .A2(_02386__PTR53), .ZN(_00768__PTR0) );
  OR2_X1 U1462 ( .A1(_02386__PTR85), .A2(_02386__PTR117), .ZN(_00768__PTR1) );
  OR2_X1 U1463 ( .A1(_00768__PTR0), .A2(_00768__PTR1), .ZN(_00769_) );
  OR2_X1 U1464 ( .A1(_00769_), .A2(_02386__PTR149), .ZN(_02388__PTR21) );
  OR2_X1 U1465 ( .A1(_02386__PTR22), .A2(_02386__PTR54), .ZN(_00770__PTR0) );
  OR2_X1 U1466 ( .A1(_02386__PTR86), .A2(_02386__PTR118), .ZN(_00770__PTR1) );
  OR2_X1 U1467 ( .A1(_00770__PTR0), .A2(_00770__PTR1), .ZN(_00771_) );
  OR2_X1 U1468 ( .A1(_00771_), .A2(_02386__PTR150), .ZN(_02388__PTR22) );
  OR2_X1 U1469 ( .A1(_02386__PTR23), .A2(_02386__PTR55), .ZN(_00772__PTR0) );
  OR2_X1 U1470 ( .A1(_02386__PTR87), .A2(_02386__PTR119), .ZN(_00772__PTR1) );
  OR2_X1 U1471 ( .A1(_00772__PTR0), .A2(_00772__PTR1), .ZN(_00773_) );
  OR2_X1 U1472 ( .A1(_00773_), .A2(_02386__PTR151), .ZN(_02388__PTR23) );
  OR2_X1 U1473 ( .A1(_02386__PTR24), .A2(_02386__PTR56), .ZN(_00774__PTR0) );
  OR2_X1 U1474 ( .A1(_02386__PTR88), .A2(_02386__PTR120), .ZN(_00774__PTR1) );
  OR2_X1 U1475 ( .A1(_00774__PTR0), .A2(_00774__PTR1), .ZN(_00775_) );
  OR2_X1 U1476 ( .A1(_00775_), .A2(_02386__PTR152), .ZN(_02388__PTR24) );
  OR2_X1 U1477 ( .A1(_02386__PTR25), .A2(_02386__PTR57), .ZN(_00776__PTR0) );
  OR2_X1 U1478 ( .A1(_02386__PTR89), .A2(_02386__PTR121), .ZN(_00776__PTR1) );
  OR2_X1 U1479 ( .A1(_00776__PTR0), .A2(_00776__PTR1), .ZN(_00777_) );
  OR2_X1 U1480 ( .A1(_00777_), .A2(_02386__PTR153), .ZN(_02388__PTR25) );
  OR2_X1 U1481 ( .A1(_02386__PTR26), .A2(_02386__PTR58), .ZN(_00778__PTR0) );
  OR2_X1 U1482 ( .A1(_02386__PTR90), .A2(_02386__PTR122), .ZN(_00778__PTR1) );
  OR2_X1 U1483 ( .A1(_00778__PTR0), .A2(_00778__PTR1), .ZN(_00779_) );
  OR2_X1 U1484 ( .A1(_00779_), .A2(_02386__PTR154), .ZN(_02388__PTR26) );
  OR2_X1 U1485 ( .A1(_02386__PTR27), .A2(_02386__PTR59), .ZN(_00780__PTR0) );
  OR2_X1 U1486 ( .A1(_02386__PTR91), .A2(_02386__PTR123), .ZN(_00780__PTR1) );
  OR2_X1 U1487 ( .A1(_00780__PTR0), .A2(_00780__PTR1), .ZN(_00781_) );
  OR2_X1 U1488 ( .A1(_00781_), .A2(_02386__PTR155), .ZN(_02388__PTR27) );
  OR2_X1 U1489 ( .A1(_02386__PTR28), .A2(_02386__PTR60), .ZN(_00782__PTR0) );
  OR2_X1 U1490 ( .A1(_02386__PTR92), .A2(_02386__PTR124), .ZN(_00782__PTR1) );
  OR2_X1 U1491 ( .A1(_00782__PTR0), .A2(_00782__PTR1), .ZN(_00783_) );
  OR2_X1 U1492 ( .A1(_00783_), .A2(_02386__PTR156), .ZN(_02388__PTR28) );
  OR2_X1 U1493 ( .A1(_02386__PTR29), .A2(_02386__PTR61), .ZN(_00784__PTR0) );
  OR2_X1 U1494 ( .A1(_02386__PTR93), .A2(_02386__PTR125), .ZN(_00784__PTR1) );
  OR2_X1 U1495 ( .A1(_00784__PTR0), .A2(_00784__PTR1), .ZN(_00785_) );
  OR2_X1 U1496 ( .A1(_00785_), .A2(_02386__PTR157), .ZN(_02388__PTR29) );
  OR2_X1 U1497 ( .A1(_02386__PTR30), .A2(_02386__PTR62), .ZN(_00786__PTR0) );
  OR2_X1 U1498 ( .A1(_02386__PTR94), .A2(_02386__PTR126), .ZN(_00786__PTR1) );
  OR2_X1 U1499 ( .A1(_00786__PTR0), .A2(_00786__PTR1), .ZN(_00787_) );
  OR2_X1 U1500 ( .A1(_00787_), .A2(_02386__PTR158), .ZN(_02388__PTR30) );
  OR2_X1 U1501 ( .A1(_02386__PTR31), .A2(_02386__PTR63), .ZN(_00788__PTR0) );
  OR2_X1 U1502 ( .A1(_02386__PTR95), .A2(_02386__PTR127), .ZN(_00788__PTR1) );
  OR2_X1 U1503 ( .A1(_00788__PTR0), .A2(_00788__PTR1), .ZN(_00789_) );
  OR2_X1 U1504 ( .A1(_00789_), .A2(_02386__PTR159), .ZN(_02388__PTR31) );
  OR2_X1 U1505 ( .A1(_02387__PTR0), .A2(_02387__PTR1), .ZN(_00790__PTR0) );
  OR2_X1 U1506 ( .A1(_02379__PTR3), .A2(_02379__PTR4), .ZN(_02148__PTR1) );
  OR2_X1 U1507 ( .A1(_00790__PTR0), .A2(_02148__PTR1), .ZN(_00791_) );
  OR2_X1 U1508 ( .A1(_00791_), .A2(_02387__PTR4), .ZN(_03168_) );
  OR2_X1 U1509 ( .A1(_02151__PTR0), .A2(_02151__PTR1), .ZN(_00792__PTR0) );
  OR2_X1 U1510 ( .A1(_02151__PTR2), .A2(_02151__PTR3), .ZN(_00792__PTR1) );
  OR2_X1 U1511 ( .A1(_00792__PTR0), .A2(_00792__PTR1), .ZN(_02153_) );
  OR2_X1 U1512 ( .A1(_00793__PTR0), .A2(_00793__PTR1), .ZN(_03018_) );
  OR2_X1 U1513 ( .A1(_02147__PTR0), .A2(_02147__PTR1), .ZN(_00794__PTR0) );
  OR2_X1 U1514 ( .A1(_02147__PTR2), .A2(_02147__PTR3), .ZN(_00794__PTR1) );
  OR2_X1 U1515 ( .A1(_00794__PTR0), .A2(_00794__PTR1), .ZN(_02149_) );
  OR2_X1 U1516 ( .A1(_02148__PTR2), .A2(_02148__PTR3), .ZN(_02379__PTR6) );
  OR2_X1 U1517 ( .A1(_00793__PTR0), .A2(_02379__PTR6), .ZN(_03017_) );
  OR2_X1 U1518 ( .A1(_02378__PTR0), .A2(_02378__PTR5), .ZN(_00795__PTR0) );
  OR2_X1 U1519 ( .A1(_02378__PTR10), .A2(_02378__PTR15), .ZN(_00795__PTR1) );
  OR2_X1 U1520 ( .A1(_02378__PTR20), .A2(_02378__PTR25), .ZN(_00795__PTR2) );
  OR2_X1 U1521 ( .A1(_00795__PTR0), .A2(_00795__PTR1), .ZN(_00796__PTR0) );
  OR2_X1 U1522 ( .A1(_00795__PTR2), .A2(_02378__PTR30), .ZN(_00796__PTR1) );
  OR2_X1 U1523 ( .A1(_00796__PTR0), .A2(_00796__PTR1), .ZN(_02380__PTR0) );
  OR2_X1 U1524 ( .A1(_02378__PTR1), .A2(_02378__PTR6), .ZN(_00797__PTR0) );
  OR2_X1 U1525 ( .A1(_02378__PTR11), .A2(_02378__PTR16), .ZN(_00797__PTR1) );
  OR2_X1 U1526 ( .A1(_02378__PTR21), .A2(_02378__PTR26), .ZN(_00797__PTR2) );
  OR2_X1 U1527 ( .A1(_00797__PTR0), .A2(_00797__PTR1), .ZN(_00798__PTR0) );
  OR2_X1 U1528 ( .A1(_00797__PTR2), .A2(_02378__PTR31), .ZN(_00798__PTR1) );
  OR2_X1 U1529 ( .A1(_00798__PTR0), .A2(_00798__PTR1), .ZN(_02380__PTR1) );
  OR2_X1 U1530 ( .A1(_02378__PTR2), .A2(_02378__PTR7), .ZN(_00799__PTR0) );
  OR2_X1 U1531 ( .A1(_02378__PTR12), .A2(_02378__PTR17), .ZN(_00799__PTR1) );
  OR2_X1 U1532 ( .A1(_02378__PTR22), .A2(_02378__PTR27), .ZN(_00799__PTR2) );
  OR2_X1 U1533 ( .A1(_00799__PTR0), .A2(_00799__PTR1), .ZN(_00800__PTR0) );
  OR2_X1 U1534 ( .A1(_00799__PTR2), .A2(_02378__PTR32), .ZN(_00800__PTR1) );
  OR2_X1 U1535 ( .A1(_00800__PTR0), .A2(_00800__PTR1), .ZN(_02380__PTR2) );
  OR2_X1 U1536 ( .A1(_02378__PTR3), .A2(_02378__PTR8), .ZN(_00801__PTR0) );
  OR2_X1 U1537 ( .A1(_02378__PTR13), .A2(_02378__PTR18), .ZN(_00801__PTR1) );
  OR2_X1 U1538 ( .A1(_02378__PTR23), .A2(_02378__PTR28), .ZN(_00801__PTR2) );
  OR2_X1 U1539 ( .A1(_00801__PTR0), .A2(_00801__PTR1), .ZN(_00802__PTR0) );
  OR2_X1 U1540 ( .A1(_00801__PTR2), .A2(_02378__PTR33), .ZN(_00802__PTR1) );
  OR2_X1 U1541 ( .A1(_00802__PTR0), .A2(_00802__PTR1), .ZN(_02380__PTR3) );
  OR2_X1 U1542 ( .A1(_02378__PTR14), .A2(_02378__PTR19), .ZN(_00803__PTR1) );
  OR2_X1 U1543 ( .A1(_02378__PTR24), .A2(_02378__PTR29), .ZN(_00803__PTR2) );
  OR2_X1 U1544 ( .A1(_00803__PTR2), .A2(_02378__PTR34), .ZN(_00804__PTR1) );
  OR2_X1 U1545 ( .A1(_00803__PTR1), .A2(_00804__PTR1), .ZN(_02380__PTR4) );
  OR2_X1 U1546 ( .A1(_02148__PTR0), .A2(_02379__PTR3), .ZN(_00805__PTR1) );
  OR2_X1 U1547 ( .A1(_02379__PTR4), .A2(_02375__PTR4), .ZN(_00805__PTR2) );
  OR2_X1 U1548 ( .A1(_00805__PTR0), .A2(_00805__PTR1), .ZN(_00806__PTR0) );
  OR2_X1 U1549 ( .A1(_00805__PTR2), .A2(_02379__PTR6), .ZN(_00806__PTR1) );
  OR2_X1 U1550 ( .A1(_00806__PTR0), .A2(_00806__PTR1), .ZN(_03166_) );
  OR2_X1 U1551 ( .A1(_02166__PTR0), .A2(_02166__PTR1), .ZN(_02168_) );
  OR2_X1 U1552 ( .A1(_02155__PTR0), .A2(_02155__PTR1), .ZN(_00807__PTR0) );
  OR2_X1 U1553 ( .A1(_02155__PTR2), .A2(_02155__PTR3), .ZN(_00807__PTR1) );
  OR2_X1 U1554 ( .A1(_00807__PTR0), .A2(_00807__PTR1), .ZN(_02157_) );
  OR2_X1 U1555 ( .A1(_02156__PTR0), .A2(_02148__PTR1), .ZN(_00808__PTR0) );
  OR2_X1 U1556 ( .A1(_02156__PTR2), .A2(_02156__PTR3), .ZN(_00808__PTR1) );
  OR2_X1 U1557 ( .A1(_00808__PTR0), .A2(_00808__PTR1), .ZN(_03019_) );
  OR2_X1 U1558 ( .A1(_02162__PTR0), .A2(_02162__PTR1), .ZN(_00809_) );
  OR2_X1 U1559 ( .A1(_00809_), .A2(_02162__PTR2), .ZN(_02164_) );
  OR2_X1 U1560 ( .A1(_02163__PTR0), .A2(_02163__PTR1), .ZN(_02167__PTR0) );
  OR2_X1 U1561 ( .A1(_02167__PTR0), .A2(_02156__PTR3), .ZN(_03021_) );
  OR2_X1 U1562 ( .A1(_02159__PTR0), .A2(_02159__PTR1), .ZN(_00810_) );
  OR2_X1 U1563 ( .A1(_00810_), .A2(_02159__PTR2), .ZN(_02160_) );
  OR2_X1 U1564 ( .A1(_00793__PTR0), .A2(_02156__PTR3), .ZN(_03020_) );
  OR2_X1 U1565 ( .A1(_02394__PTR0), .A2(_02394__PTR32), .ZN(_00811__PTR0) );
  OR2_X1 U1566 ( .A1(_02394__PTR64), .A2(_02394__PTR96), .ZN(_00811__PTR1) );
  OR2_X1 U1567 ( .A1(_00811__PTR0), .A2(_00811__PTR1), .ZN(_02395__PTR0) );
  OR2_X1 U1568 ( .A1(_02394__PTR1), .A2(_02394__PTR33), .ZN(_00812__PTR0) );
  OR2_X1 U1569 ( .A1(_02394__PTR65), .A2(_02394__PTR97), .ZN(_00812__PTR1) );
  OR2_X1 U1570 ( .A1(_00812__PTR0), .A2(_00812__PTR1), .ZN(_02395__PTR1) );
  OR2_X1 U1571 ( .A1(_02394__PTR2), .A2(_02394__PTR34), .ZN(_00813__PTR0) );
  OR2_X1 U1572 ( .A1(_02394__PTR66), .A2(_02394__PTR98), .ZN(_00813__PTR1) );
  OR2_X1 U1573 ( .A1(_00813__PTR0), .A2(_00813__PTR1), .ZN(_02395__PTR2) );
  OR2_X1 U1574 ( .A1(_02394__PTR3), .A2(_02394__PTR35), .ZN(_00814__PTR0) );
  OR2_X1 U1575 ( .A1(_02394__PTR67), .A2(_02394__PTR99), .ZN(_00814__PTR1) );
  OR2_X1 U1576 ( .A1(_00814__PTR0), .A2(_00814__PTR1), .ZN(_02395__PTR3) );
  OR2_X1 U1577 ( .A1(_02394__PTR4), .A2(_02394__PTR36), .ZN(_00815__PTR0) );
  OR2_X1 U1578 ( .A1(_02394__PTR68), .A2(_02394__PTR100), .ZN(_00815__PTR1) );
  OR2_X1 U1579 ( .A1(_00815__PTR0), .A2(_00815__PTR1), .ZN(_02395__PTR4) );
  OR2_X1 U1580 ( .A1(_02394__PTR5), .A2(_02394__PTR37), .ZN(_00816__PTR0) );
  OR2_X1 U1581 ( .A1(_02394__PTR69), .A2(_02394__PTR101), .ZN(_00816__PTR1) );
  OR2_X1 U1582 ( .A1(_00816__PTR0), .A2(_00816__PTR1), .ZN(_02395__PTR5) );
  OR2_X1 U1583 ( .A1(_02394__PTR6), .A2(_02394__PTR38), .ZN(_00817__PTR0) );
  OR2_X1 U1584 ( .A1(_02394__PTR70), .A2(_02394__PTR102), .ZN(_00817__PTR1) );
  OR2_X1 U1585 ( .A1(_00817__PTR0), .A2(_00817__PTR1), .ZN(_02395__PTR6) );
  OR2_X1 U1586 ( .A1(_02394__PTR7), .A2(_02394__PTR39), .ZN(_00818__PTR0) );
  OR2_X1 U1587 ( .A1(_02394__PTR71), .A2(_02394__PTR103), .ZN(_00818__PTR1) );
  OR2_X1 U1588 ( .A1(_00818__PTR0), .A2(_00818__PTR1), .ZN(_02395__PTR7) );
  OR2_X1 U1589 ( .A1(_02394__PTR8), .A2(_02394__PTR40), .ZN(_00819__PTR0) );
  OR2_X1 U1590 ( .A1(_02394__PTR72), .A2(_02394__PTR104), .ZN(_00819__PTR1) );
  OR2_X1 U1591 ( .A1(_00819__PTR0), .A2(_00819__PTR1), .ZN(_02395__PTR8) );
  OR2_X1 U1592 ( .A1(_02394__PTR9), .A2(_02394__PTR41), .ZN(_00820__PTR0) );
  OR2_X1 U1593 ( .A1(_02394__PTR73), .A2(_02394__PTR105), .ZN(_00820__PTR1) );
  OR2_X1 U1594 ( .A1(_00820__PTR0), .A2(_00820__PTR1), .ZN(_02395__PTR9) );
  OR2_X1 U1595 ( .A1(_02394__PTR10), .A2(_02394__PTR42), .ZN(_00821__PTR0) );
  OR2_X1 U1596 ( .A1(_02394__PTR74), .A2(_02394__PTR106), .ZN(_00821__PTR1) );
  OR2_X1 U1597 ( .A1(_00821__PTR0), .A2(_00821__PTR1), .ZN(_02395__PTR10) );
  OR2_X1 U1598 ( .A1(_02394__PTR11), .A2(_02394__PTR43), .ZN(_00822__PTR0) );
  OR2_X1 U1599 ( .A1(_02394__PTR75), .A2(_02394__PTR107), .ZN(_00822__PTR1) );
  OR2_X1 U1600 ( .A1(_00822__PTR0), .A2(_00822__PTR1), .ZN(_02395__PTR11) );
  OR2_X1 U1601 ( .A1(_02394__PTR12), .A2(_02394__PTR44), .ZN(_00823__PTR0) );
  OR2_X1 U1602 ( .A1(_02394__PTR76), .A2(_02394__PTR108), .ZN(_00823__PTR1) );
  OR2_X1 U1603 ( .A1(_00823__PTR0), .A2(_00823__PTR1), .ZN(_02395__PTR12) );
  OR2_X1 U1604 ( .A1(_02394__PTR13), .A2(_02394__PTR45), .ZN(_00824__PTR0) );
  OR2_X1 U1605 ( .A1(_02394__PTR77), .A2(_02394__PTR109), .ZN(_00824__PTR1) );
  OR2_X1 U1606 ( .A1(_00824__PTR0), .A2(_00824__PTR1), .ZN(_02395__PTR13) );
  OR2_X1 U1607 ( .A1(_02394__PTR14), .A2(_02394__PTR46), .ZN(_00825__PTR0) );
  OR2_X1 U1608 ( .A1(_02394__PTR78), .A2(_02394__PTR110), .ZN(_00825__PTR1) );
  OR2_X1 U1609 ( .A1(_00825__PTR0), .A2(_00825__PTR1), .ZN(_02395__PTR14) );
  OR2_X1 U1610 ( .A1(_02394__PTR15), .A2(_02394__PTR47), .ZN(_00826__PTR0) );
  OR2_X1 U1611 ( .A1(_02394__PTR79), .A2(_02394__PTR111), .ZN(_00826__PTR1) );
  OR2_X1 U1612 ( .A1(_00826__PTR0), .A2(_00826__PTR1), .ZN(_02395__PTR15) );
  OR2_X1 U1613 ( .A1(_02394__PTR16), .A2(_02394__PTR48), .ZN(_00827__PTR0) );
  OR2_X1 U1614 ( .A1(_02394__PTR80), .A2(_02394__PTR112), .ZN(_00827__PTR1) );
  OR2_X1 U1615 ( .A1(_00827__PTR0), .A2(_00827__PTR1), .ZN(_02395__PTR16) );
  OR2_X1 U1616 ( .A1(_02394__PTR17), .A2(_02394__PTR49), .ZN(_00828__PTR0) );
  OR2_X1 U1617 ( .A1(_02394__PTR81), .A2(_02394__PTR113), .ZN(_00828__PTR1) );
  OR2_X1 U1618 ( .A1(_00828__PTR0), .A2(_00828__PTR1), .ZN(_02395__PTR17) );
  OR2_X1 U1619 ( .A1(_02394__PTR18), .A2(_02394__PTR50), .ZN(_00829__PTR0) );
  OR2_X1 U1620 ( .A1(_02394__PTR82), .A2(_02394__PTR114), .ZN(_00829__PTR1) );
  OR2_X1 U1621 ( .A1(_00829__PTR0), .A2(_00829__PTR1), .ZN(_02395__PTR18) );
  OR2_X1 U1622 ( .A1(_02394__PTR19), .A2(_02394__PTR51), .ZN(_00830__PTR0) );
  OR2_X1 U1623 ( .A1(_02394__PTR83), .A2(_02394__PTR115), .ZN(_00830__PTR1) );
  OR2_X1 U1624 ( .A1(_00830__PTR0), .A2(_00830__PTR1), .ZN(_02395__PTR19) );
  OR2_X1 U1625 ( .A1(_02394__PTR20), .A2(_02394__PTR52), .ZN(_00831__PTR0) );
  OR2_X1 U1626 ( .A1(_02394__PTR84), .A2(_02394__PTR116), .ZN(_00831__PTR1) );
  OR2_X1 U1627 ( .A1(_00831__PTR0), .A2(_00831__PTR1), .ZN(_02395__PTR20) );
  OR2_X1 U1628 ( .A1(_02394__PTR21), .A2(_02394__PTR53), .ZN(_00832__PTR0) );
  OR2_X1 U1629 ( .A1(_02394__PTR85), .A2(_02394__PTR117), .ZN(_00832__PTR1) );
  OR2_X1 U1630 ( .A1(_00832__PTR0), .A2(_00832__PTR1), .ZN(_02395__PTR21) );
  OR2_X1 U1631 ( .A1(_02394__PTR22), .A2(_02394__PTR54), .ZN(_00833__PTR0) );
  OR2_X1 U1632 ( .A1(_02394__PTR86), .A2(_02394__PTR118), .ZN(_00833__PTR1) );
  OR2_X1 U1633 ( .A1(_00833__PTR0), .A2(_00833__PTR1), .ZN(_02395__PTR22) );
  OR2_X1 U1634 ( .A1(_02394__PTR23), .A2(_02394__PTR55), .ZN(_00834__PTR0) );
  OR2_X1 U1635 ( .A1(_02394__PTR87), .A2(_02394__PTR119), .ZN(_00834__PTR1) );
  OR2_X1 U1636 ( .A1(_00834__PTR0), .A2(_00834__PTR1), .ZN(_02395__PTR23) );
  OR2_X1 U1637 ( .A1(_02394__PTR24), .A2(_02394__PTR56), .ZN(_00835__PTR0) );
  OR2_X1 U1638 ( .A1(_02394__PTR88), .A2(_02394__PTR120), .ZN(_00835__PTR1) );
  OR2_X1 U1639 ( .A1(_00835__PTR0), .A2(_00835__PTR1), .ZN(_02395__PTR24) );
  OR2_X1 U1640 ( .A1(_02394__PTR25), .A2(_02394__PTR57), .ZN(_00836__PTR0) );
  OR2_X1 U1641 ( .A1(_02394__PTR89), .A2(_02394__PTR121), .ZN(_00836__PTR1) );
  OR2_X1 U1642 ( .A1(_00836__PTR0), .A2(_00836__PTR1), .ZN(_02395__PTR25) );
  OR2_X1 U1643 ( .A1(_02394__PTR26), .A2(_02394__PTR58), .ZN(_00837__PTR0) );
  OR2_X1 U1644 ( .A1(_02394__PTR90), .A2(_02394__PTR122), .ZN(_00837__PTR1) );
  OR2_X1 U1645 ( .A1(_00837__PTR0), .A2(_00837__PTR1), .ZN(_02395__PTR26) );
  OR2_X1 U1646 ( .A1(_02394__PTR27), .A2(_02394__PTR59), .ZN(_00838__PTR0) );
  OR2_X1 U1647 ( .A1(_02394__PTR91), .A2(_02394__PTR123), .ZN(_00838__PTR1) );
  OR2_X1 U1648 ( .A1(_00838__PTR0), .A2(_00838__PTR1), .ZN(_02395__PTR27) );
  OR2_X1 U1649 ( .A1(_02394__PTR28), .A2(_02394__PTR60), .ZN(_00839__PTR0) );
  OR2_X1 U1650 ( .A1(_02394__PTR92), .A2(_02394__PTR124), .ZN(_00839__PTR1) );
  OR2_X1 U1651 ( .A1(_00839__PTR0), .A2(_00839__PTR1), .ZN(_02395__PTR28) );
  OR2_X1 U1652 ( .A1(_02394__PTR29), .A2(_02394__PTR61), .ZN(_00840__PTR0) );
  OR2_X1 U1653 ( .A1(_02394__PTR93), .A2(_02394__PTR125), .ZN(_00840__PTR1) );
  OR2_X1 U1654 ( .A1(_00840__PTR0), .A2(_00840__PTR1), .ZN(_02395__PTR29) );
  OR2_X1 U1655 ( .A1(_02394__PTR30), .A2(_02394__PTR62), .ZN(_00841__PTR0) );
  OR2_X1 U1656 ( .A1(_02394__PTR94), .A2(_02394__PTR126), .ZN(_00841__PTR1) );
  OR2_X1 U1657 ( .A1(_00841__PTR0), .A2(_00841__PTR1), .ZN(_02395__PTR30) );
  OR2_X1 U1658 ( .A1(_02394__PTR31), .A2(_02394__PTR63), .ZN(_00842__PTR0) );
  OR2_X1 U1659 ( .A1(_02394__PTR95), .A2(_02394__PTR127), .ZN(_00842__PTR1) );
  OR2_X1 U1660 ( .A1(_00842__PTR0), .A2(_00842__PTR1), .ZN(_02395__PTR31) );
  OR2_X1 U1661 ( .A1(_02156__PTR3), .A2(_02163__PTR0), .ZN(_00843__PTR0) );
  OR2_X1 U1662 ( .A1(_02156__PTR2), .A2(_02379__PTR4), .ZN(_02163__PTR1) );
  OR2_X1 U1663 ( .A1(_00843__PTR0), .A2(_02163__PTR1), .ZN(_03170_) );
  OR2_X1 U1664 ( .A1(_02374__PTR0), .A2(_02374__PTR32), .ZN(_00844__PTR0) );
  OR2_X1 U1665 ( .A1(_02374__PTR64), .A2(_02374__PTR96), .ZN(_00844__PTR1) );
  OR2_X1 U1666 ( .A1(_02374__PTR128), .A2(_02374__PTR160), .ZN(_00844__PTR2) );
  OR2_X1 U1667 ( .A1(_00844__PTR0), .A2(_00844__PTR1), .ZN(_00845__PTR0) );
  OR2_X1 U1668 ( .A1(_00844__PTR2), .A2(_02374__PTR192), .ZN(_00845__PTR1) );
  OR2_X1 U1669 ( .A1(_00845__PTR0), .A2(_00845__PTR1), .ZN(_02376__PTR0) );
  OR2_X1 U1670 ( .A1(_02374__PTR1), .A2(_02374__PTR33), .ZN(_00846__PTR0) );
  OR2_X1 U1671 ( .A1(_02374__PTR65), .A2(_02374__PTR97), .ZN(_00846__PTR1) );
  OR2_X1 U1672 ( .A1(_02374__PTR129), .A2(_02374__PTR161), .ZN(_00846__PTR2) );
  OR2_X1 U1673 ( .A1(_00846__PTR0), .A2(_00846__PTR1), .ZN(_00847__PTR0) );
  OR2_X1 U1674 ( .A1(_00846__PTR2), .A2(_02374__PTR193), .ZN(_00847__PTR1) );
  OR2_X1 U1675 ( .A1(_00847__PTR0), .A2(_00847__PTR1), .ZN(_02376__PTR1) );
  OR2_X1 U1676 ( .A1(_02374__PTR2), .A2(_02374__PTR34), .ZN(_00848__PTR0) );
  OR2_X1 U1677 ( .A1(_02374__PTR66), .A2(_02374__PTR98), .ZN(_00848__PTR1) );
  OR2_X1 U1678 ( .A1(_02374__PTR130), .A2(_02374__PTR162), .ZN(_00848__PTR2) );
  OR2_X1 U1679 ( .A1(_00848__PTR0), .A2(_00848__PTR1), .ZN(_00849__PTR0) );
  OR2_X1 U1680 ( .A1(_00848__PTR2), .A2(_02374__PTR194), .ZN(_00849__PTR1) );
  OR2_X1 U1681 ( .A1(_00849__PTR0), .A2(_00849__PTR1), .ZN(_02376__PTR2) );
  OR2_X1 U1682 ( .A1(_02374__PTR3), .A2(_02374__PTR35), .ZN(_00850__PTR0) );
  OR2_X1 U1683 ( .A1(_02374__PTR67), .A2(_02374__PTR99), .ZN(_00850__PTR1) );
  OR2_X1 U1684 ( .A1(_02374__PTR131), .A2(_02374__PTR163), .ZN(_00850__PTR2) );
  OR2_X1 U1685 ( .A1(_00850__PTR0), .A2(_00850__PTR1), .ZN(_00851__PTR0) );
  OR2_X1 U1686 ( .A1(_00850__PTR2), .A2(_02374__PTR195), .ZN(_00851__PTR1) );
  OR2_X1 U1687 ( .A1(_00851__PTR0), .A2(_00851__PTR1), .ZN(_02376__PTR3) );
  OR2_X1 U1688 ( .A1(_02374__PTR4), .A2(_02374__PTR36), .ZN(_00852__PTR0) );
  OR2_X1 U1689 ( .A1(_02374__PTR68), .A2(_02374__PTR100), .ZN(_00852__PTR1) );
  OR2_X1 U1690 ( .A1(_02374__PTR132), .A2(_02374__PTR164), .ZN(_00852__PTR2) );
  OR2_X1 U1691 ( .A1(_00852__PTR0), .A2(_00852__PTR1), .ZN(_00853__PTR0) );
  OR2_X1 U1692 ( .A1(_00852__PTR2), .A2(_02374__PTR196), .ZN(_00853__PTR1) );
  OR2_X1 U1693 ( .A1(_00853__PTR0), .A2(_00853__PTR1), .ZN(_02376__PTR4) );
  OR2_X1 U1694 ( .A1(_02374__PTR5), .A2(_02374__PTR37), .ZN(_00854__PTR0) );
  OR2_X1 U1695 ( .A1(_02374__PTR69), .A2(_02374__PTR101), .ZN(_00854__PTR1) );
  OR2_X1 U1696 ( .A1(_02374__PTR133), .A2(_02374__PTR165), .ZN(_00854__PTR2) );
  OR2_X1 U1697 ( .A1(_00854__PTR0), .A2(_00854__PTR1), .ZN(_00855__PTR0) );
  OR2_X1 U1698 ( .A1(_00854__PTR2), .A2(_02374__PTR197), .ZN(_00855__PTR1) );
  OR2_X1 U1699 ( .A1(_00855__PTR0), .A2(_00855__PTR1), .ZN(_02376__PTR5) );
  OR2_X1 U1700 ( .A1(_02374__PTR6), .A2(_02374__PTR38), .ZN(_00856__PTR0) );
  OR2_X1 U1701 ( .A1(_02374__PTR70), .A2(_02374__PTR102), .ZN(_00856__PTR1) );
  OR2_X1 U1702 ( .A1(_02374__PTR134), .A2(_02374__PTR166), .ZN(_00856__PTR2) );
  OR2_X1 U1703 ( .A1(_00856__PTR0), .A2(_00856__PTR1), .ZN(_00857__PTR0) );
  OR2_X1 U1704 ( .A1(_00856__PTR2), .A2(_02374__PTR198), .ZN(_00857__PTR1) );
  OR2_X1 U1705 ( .A1(_00857__PTR0), .A2(_00857__PTR1), .ZN(_02376__PTR6) );
  OR2_X1 U1706 ( .A1(_02374__PTR7), .A2(_02374__PTR39), .ZN(_00858__PTR0) );
  OR2_X1 U1707 ( .A1(_02374__PTR71), .A2(_02374__PTR103), .ZN(_00858__PTR1) );
  OR2_X1 U1708 ( .A1(_02374__PTR135), .A2(_02374__PTR167), .ZN(_00858__PTR2) );
  OR2_X1 U1709 ( .A1(_00858__PTR0), .A2(_00858__PTR1), .ZN(_00859__PTR0) );
  OR2_X1 U1710 ( .A1(_00858__PTR2), .A2(_02374__PTR199), .ZN(_00859__PTR1) );
  OR2_X1 U1711 ( .A1(_00859__PTR0), .A2(_00859__PTR1), .ZN(_02376__PTR7) );
  OR2_X1 U1712 ( .A1(_02374__PTR8), .A2(_02374__PTR40), .ZN(_00860__PTR0) );
  OR2_X1 U1713 ( .A1(_02374__PTR72), .A2(_02374__PTR104), .ZN(_00860__PTR1) );
  OR2_X1 U1714 ( .A1(_02374__PTR136), .A2(_02374__PTR168), .ZN(_00860__PTR2) );
  OR2_X1 U1715 ( .A1(_00860__PTR0), .A2(_00860__PTR1), .ZN(_00861__PTR0) );
  OR2_X1 U1716 ( .A1(_00860__PTR2), .A2(_02374__PTR200), .ZN(_00861__PTR1) );
  OR2_X1 U1717 ( .A1(_00861__PTR0), .A2(_00861__PTR1), .ZN(_02376__PTR8) );
  OR2_X1 U1718 ( .A1(_02374__PTR9), .A2(_02374__PTR41), .ZN(_00862__PTR0) );
  OR2_X1 U1719 ( .A1(_02374__PTR73), .A2(_02374__PTR105), .ZN(_00862__PTR1) );
  OR2_X1 U1720 ( .A1(_02374__PTR137), .A2(_02374__PTR169), .ZN(_00862__PTR2) );
  OR2_X1 U1721 ( .A1(_00862__PTR0), .A2(_00862__PTR1), .ZN(_00863__PTR0) );
  OR2_X1 U1722 ( .A1(_00862__PTR2), .A2(_02374__PTR201), .ZN(_00863__PTR1) );
  OR2_X1 U1723 ( .A1(_00863__PTR0), .A2(_00863__PTR1), .ZN(_02376__PTR9) );
  OR2_X1 U1724 ( .A1(_02374__PTR10), .A2(_02374__PTR42), .ZN(_00864__PTR0) );
  OR2_X1 U1725 ( .A1(_02374__PTR74), .A2(_02374__PTR106), .ZN(_00864__PTR1) );
  OR2_X1 U1726 ( .A1(_02374__PTR138), .A2(_02374__PTR170), .ZN(_00864__PTR2) );
  OR2_X1 U1727 ( .A1(_00864__PTR0), .A2(_00864__PTR1), .ZN(_00865__PTR0) );
  OR2_X1 U1728 ( .A1(_00864__PTR2), .A2(_02374__PTR202), .ZN(_00865__PTR1) );
  OR2_X1 U1729 ( .A1(_00865__PTR0), .A2(_00865__PTR1), .ZN(_02376__PTR10) );
  OR2_X1 U1730 ( .A1(_02374__PTR11), .A2(_02374__PTR43), .ZN(_00866__PTR0) );
  OR2_X1 U1731 ( .A1(_02374__PTR75), .A2(_02374__PTR107), .ZN(_00866__PTR1) );
  OR2_X1 U1732 ( .A1(_02374__PTR139), .A2(_02374__PTR171), .ZN(_00866__PTR2) );
  OR2_X1 U1733 ( .A1(_00866__PTR0), .A2(_00866__PTR1), .ZN(_00867__PTR0) );
  OR2_X1 U1734 ( .A1(_00866__PTR2), .A2(_02374__PTR203), .ZN(_00867__PTR1) );
  OR2_X1 U1735 ( .A1(_00867__PTR0), .A2(_00867__PTR1), .ZN(_02376__PTR11) );
  OR2_X1 U1736 ( .A1(_02374__PTR12), .A2(_02374__PTR44), .ZN(_00868__PTR0) );
  OR2_X1 U1737 ( .A1(_02374__PTR76), .A2(_02374__PTR108), .ZN(_00868__PTR1) );
  OR2_X1 U1738 ( .A1(_02374__PTR140), .A2(_02374__PTR172), .ZN(_00868__PTR2) );
  OR2_X1 U1739 ( .A1(_00868__PTR0), .A2(_00868__PTR1), .ZN(_00869__PTR0) );
  OR2_X1 U1740 ( .A1(_00868__PTR2), .A2(_02374__PTR204), .ZN(_00869__PTR1) );
  OR2_X1 U1741 ( .A1(_00869__PTR0), .A2(_00869__PTR1), .ZN(_02376__PTR12) );
  OR2_X1 U1742 ( .A1(_02374__PTR13), .A2(_02374__PTR45), .ZN(_00870__PTR0) );
  OR2_X1 U1743 ( .A1(_02374__PTR77), .A2(_02374__PTR109), .ZN(_00870__PTR1) );
  OR2_X1 U1744 ( .A1(_02374__PTR141), .A2(_02374__PTR173), .ZN(_00870__PTR2) );
  OR2_X1 U1745 ( .A1(_00870__PTR0), .A2(_00870__PTR1), .ZN(_00871__PTR0) );
  OR2_X1 U1746 ( .A1(_00870__PTR2), .A2(_02374__PTR205), .ZN(_00871__PTR1) );
  OR2_X1 U1747 ( .A1(_00871__PTR0), .A2(_00871__PTR1), .ZN(_02376__PTR13) );
  OR2_X1 U1748 ( .A1(_02374__PTR14), .A2(_02374__PTR46), .ZN(_00872__PTR0) );
  OR2_X1 U1749 ( .A1(_02374__PTR78), .A2(_02374__PTR110), .ZN(_00872__PTR1) );
  OR2_X1 U1750 ( .A1(_02374__PTR142), .A2(_02374__PTR174), .ZN(_00872__PTR2) );
  OR2_X1 U1751 ( .A1(_00872__PTR0), .A2(_00872__PTR1), .ZN(_00873__PTR0) );
  OR2_X1 U1752 ( .A1(_00872__PTR2), .A2(_02374__PTR206), .ZN(_00873__PTR1) );
  OR2_X1 U1753 ( .A1(_00873__PTR0), .A2(_00873__PTR1), .ZN(_02376__PTR14) );
  OR2_X1 U1754 ( .A1(_02374__PTR15), .A2(_02374__PTR47), .ZN(_00874__PTR0) );
  OR2_X1 U1755 ( .A1(_02374__PTR79), .A2(_02374__PTR111), .ZN(_00874__PTR1) );
  OR2_X1 U1756 ( .A1(_02374__PTR143), .A2(_02374__PTR175), .ZN(_00874__PTR2) );
  OR2_X1 U1757 ( .A1(_00874__PTR0), .A2(_00874__PTR1), .ZN(_00875__PTR0) );
  OR2_X1 U1758 ( .A1(_00874__PTR2), .A2(_02374__PTR207), .ZN(_00875__PTR1) );
  OR2_X1 U1759 ( .A1(_00875__PTR0), .A2(_00875__PTR1), .ZN(_02376__PTR15) );
  OR2_X1 U1760 ( .A1(_02374__PTR16), .A2(_02374__PTR48), .ZN(_00876__PTR0) );
  OR2_X1 U1761 ( .A1(_02374__PTR80), .A2(_02374__PTR112), .ZN(_00876__PTR1) );
  OR2_X1 U1762 ( .A1(_02374__PTR144), .A2(_02374__PTR176), .ZN(_00876__PTR2) );
  OR2_X1 U1763 ( .A1(_00876__PTR0), .A2(_00876__PTR1), .ZN(_00877__PTR0) );
  OR2_X1 U1764 ( .A1(_00876__PTR2), .A2(_02374__PTR208), .ZN(_00877__PTR1) );
  OR2_X1 U1765 ( .A1(_00877__PTR0), .A2(_00877__PTR1), .ZN(_02376__PTR16) );
  OR2_X1 U1766 ( .A1(_02374__PTR17), .A2(_02374__PTR49), .ZN(_00878__PTR0) );
  OR2_X1 U1767 ( .A1(_02374__PTR81), .A2(_02374__PTR113), .ZN(_00878__PTR1) );
  OR2_X1 U1768 ( .A1(_02374__PTR145), .A2(_02374__PTR177), .ZN(_00878__PTR2) );
  OR2_X1 U1769 ( .A1(_00878__PTR0), .A2(_00878__PTR1), .ZN(_00879__PTR0) );
  OR2_X1 U1770 ( .A1(_00878__PTR2), .A2(_02374__PTR209), .ZN(_00879__PTR1) );
  OR2_X1 U1771 ( .A1(_00879__PTR0), .A2(_00879__PTR1), .ZN(_02376__PTR17) );
  OR2_X1 U1772 ( .A1(_02374__PTR18), .A2(_02374__PTR50), .ZN(_00880__PTR0) );
  OR2_X1 U1773 ( .A1(_02374__PTR82), .A2(_02374__PTR114), .ZN(_00880__PTR1) );
  OR2_X1 U1774 ( .A1(_02374__PTR146), .A2(_02374__PTR178), .ZN(_00880__PTR2) );
  OR2_X1 U1775 ( .A1(_00880__PTR0), .A2(_00880__PTR1), .ZN(_00881__PTR0) );
  OR2_X1 U1776 ( .A1(_00880__PTR2), .A2(_02374__PTR210), .ZN(_00881__PTR1) );
  OR2_X1 U1777 ( .A1(_00881__PTR0), .A2(_00881__PTR1), .ZN(_02376__PTR18) );
  OR2_X1 U1778 ( .A1(_02374__PTR19), .A2(_02374__PTR51), .ZN(_00882__PTR0) );
  OR2_X1 U1779 ( .A1(_02374__PTR83), .A2(_02374__PTR115), .ZN(_00882__PTR1) );
  OR2_X1 U1780 ( .A1(_02374__PTR147), .A2(_02374__PTR179), .ZN(_00882__PTR2) );
  OR2_X1 U1781 ( .A1(_00882__PTR0), .A2(_00882__PTR1), .ZN(_00883__PTR0) );
  OR2_X1 U1782 ( .A1(_00882__PTR2), .A2(_02374__PTR211), .ZN(_00883__PTR1) );
  OR2_X1 U1783 ( .A1(_00883__PTR0), .A2(_00883__PTR1), .ZN(_02376__PTR19) );
  OR2_X1 U1784 ( .A1(_02374__PTR20), .A2(_02374__PTR52), .ZN(_00884__PTR0) );
  OR2_X1 U1785 ( .A1(_02374__PTR84), .A2(_02374__PTR116), .ZN(_00884__PTR1) );
  OR2_X1 U1786 ( .A1(_02374__PTR148), .A2(_02374__PTR180), .ZN(_00884__PTR2) );
  OR2_X1 U1787 ( .A1(_00884__PTR0), .A2(_00884__PTR1), .ZN(_00885__PTR0) );
  OR2_X1 U1788 ( .A1(_00884__PTR2), .A2(_02374__PTR212), .ZN(_00885__PTR1) );
  OR2_X1 U1789 ( .A1(_00885__PTR0), .A2(_00885__PTR1), .ZN(_02376__PTR20) );
  OR2_X1 U1790 ( .A1(_02374__PTR21), .A2(_02374__PTR53), .ZN(_00886__PTR0) );
  OR2_X1 U1791 ( .A1(_02374__PTR85), .A2(_02374__PTR117), .ZN(_00886__PTR1) );
  OR2_X1 U1792 ( .A1(_02374__PTR149), .A2(_02374__PTR181), .ZN(_00886__PTR2) );
  OR2_X1 U1793 ( .A1(_00886__PTR0), .A2(_00886__PTR1), .ZN(_00887__PTR0) );
  OR2_X1 U1794 ( .A1(_00886__PTR2), .A2(_02374__PTR213), .ZN(_00887__PTR1) );
  OR2_X1 U1795 ( .A1(_00887__PTR0), .A2(_00887__PTR1), .ZN(_02376__PTR21) );
  OR2_X1 U1796 ( .A1(_02374__PTR22), .A2(_02374__PTR54), .ZN(_00888__PTR0) );
  OR2_X1 U1797 ( .A1(_02374__PTR86), .A2(_02374__PTR118), .ZN(_00888__PTR1) );
  OR2_X1 U1798 ( .A1(_02374__PTR150), .A2(_02374__PTR182), .ZN(_00888__PTR2) );
  OR2_X1 U1799 ( .A1(_00888__PTR0), .A2(_00888__PTR1), .ZN(_00889__PTR0) );
  OR2_X1 U1800 ( .A1(_00888__PTR2), .A2(_02374__PTR214), .ZN(_00889__PTR1) );
  OR2_X1 U1801 ( .A1(_00889__PTR0), .A2(_00889__PTR1), .ZN(_02376__PTR22) );
  OR2_X1 U1802 ( .A1(_02374__PTR23), .A2(_02374__PTR55), .ZN(_00890__PTR0) );
  OR2_X1 U1803 ( .A1(_02374__PTR87), .A2(_02374__PTR119), .ZN(_00890__PTR1) );
  OR2_X1 U1804 ( .A1(_02374__PTR151), .A2(_02374__PTR183), .ZN(_00890__PTR2) );
  OR2_X1 U1805 ( .A1(_00890__PTR0), .A2(_00890__PTR1), .ZN(_00891__PTR0) );
  OR2_X1 U1806 ( .A1(_00890__PTR2), .A2(_02374__PTR215), .ZN(_00891__PTR1) );
  OR2_X1 U1807 ( .A1(_00891__PTR0), .A2(_00891__PTR1), .ZN(_02376__PTR23) );
  OR2_X1 U1808 ( .A1(_02374__PTR24), .A2(_02374__PTR56), .ZN(_00892__PTR0) );
  OR2_X1 U1809 ( .A1(_02374__PTR88), .A2(_02374__PTR120), .ZN(_00892__PTR1) );
  OR2_X1 U1810 ( .A1(_02374__PTR152), .A2(_02374__PTR184), .ZN(_00892__PTR2) );
  OR2_X1 U1811 ( .A1(_00892__PTR0), .A2(_00892__PTR1), .ZN(_00893__PTR0) );
  OR2_X1 U1812 ( .A1(_00892__PTR2), .A2(_02374__PTR216), .ZN(_00893__PTR1) );
  OR2_X1 U1813 ( .A1(_00893__PTR0), .A2(_00893__PTR1), .ZN(_02376__PTR24) );
  OR2_X1 U1814 ( .A1(_02374__PTR25), .A2(_02374__PTR57), .ZN(_00894__PTR0) );
  OR2_X1 U1815 ( .A1(_02374__PTR89), .A2(_02374__PTR121), .ZN(_00894__PTR1) );
  OR2_X1 U1816 ( .A1(_02374__PTR153), .A2(_02374__PTR185), .ZN(_00894__PTR2) );
  OR2_X1 U1817 ( .A1(_00894__PTR0), .A2(_00894__PTR1), .ZN(_00895__PTR0) );
  OR2_X1 U1818 ( .A1(_00894__PTR2), .A2(_02374__PTR217), .ZN(_00895__PTR1) );
  OR2_X1 U1819 ( .A1(_00895__PTR0), .A2(_00895__PTR1), .ZN(_02376__PTR25) );
  OR2_X1 U1820 ( .A1(_02374__PTR26), .A2(_02374__PTR58), .ZN(_00896__PTR0) );
  OR2_X1 U1821 ( .A1(_02374__PTR90), .A2(_02374__PTR122), .ZN(_00896__PTR1) );
  OR2_X1 U1822 ( .A1(_02374__PTR154), .A2(_02374__PTR186), .ZN(_00896__PTR2) );
  OR2_X1 U1823 ( .A1(_00896__PTR0), .A2(_00896__PTR1), .ZN(_00897__PTR0) );
  OR2_X1 U1824 ( .A1(_00896__PTR2), .A2(_02374__PTR218), .ZN(_00897__PTR1) );
  OR2_X1 U1825 ( .A1(_00897__PTR0), .A2(_00897__PTR1), .ZN(_02376__PTR26) );
  OR2_X1 U1826 ( .A1(_02374__PTR27), .A2(_02374__PTR59), .ZN(_00898__PTR0) );
  OR2_X1 U1827 ( .A1(_02374__PTR91), .A2(_02374__PTR123), .ZN(_00898__PTR1) );
  OR2_X1 U1828 ( .A1(_02374__PTR155), .A2(_02374__PTR187), .ZN(_00898__PTR2) );
  OR2_X1 U1829 ( .A1(_00898__PTR0), .A2(_00898__PTR1), .ZN(_00899__PTR0) );
  OR2_X1 U1830 ( .A1(_00898__PTR2), .A2(_02374__PTR219), .ZN(_00899__PTR1) );
  OR2_X1 U1831 ( .A1(_00899__PTR0), .A2(_00899__PTR1), .ZN(_02376__PTR27) );
  OR2_X1 U1832 ( .A1(_02374__PTR28), .A2(_02374__PTR60), .ZN(_00900__PTR0) );
  OR2_X1 U1833 ( .A1(_02374__PTR92), .A2(_02374__PTR124), .ZN(_00900__PTR1) );
  OR2_X1 U1834 ( .A1(_02374__PTR156), .A2(_02374__PTR188), .ZN(_00900__PTR2) );
  OR2_X1 U1835 ( .A1(_00900__PTR0), .A2(_00900__PTR1), .ZN(_00901__PTR0) );
  OR2_X1 U1836 ( .A1(_00900__PTR2), .A2(_02374__PTR220), .ZN(_00901__PTR1) );
  OR2_X1 U1837 ( .A1(_00901__PTR0), .A2(_00901__PTR1), .ZN(_02376__PTR28) );
  OR2_X1 U1838 ( .A1(_02374__PTR29), .A2(_02374__PTR61), .ZN(_00902__PTR0) );
  OR2_X1 U1839 ( .A1(_02374__PTR93), .A2(_02374__PTR125), .ZN(_00902__PTR1) );
  OR2_X1 U1840 ( .A1(_02374__PTR157), .A2(_02374__PTR189), .ZN(_00902__PTR2) );
  OR2_X1 U1841 ( .A1(_00902__PTR0), .A2(_00902__PTR1), .ZN(_00903__PTR0) );
  OR2_X1 U1842 ( .A1(_00902__PTR2), .A2(_02374__PTR221), .ZN(_00903__PTR1) );
  OR2_X1 U1843 ( .A1(_00903__PTR0), .A2(_00903__PTR1), .ZN(_02376__PTR29) );
  OR2_X1 U1844 ( .A1(_02374__PTR30), .A2(_02374__PTR62), .ZN(_00904__PTR0) );
  OR2_X1 U1845 ( .A1(_02374__PTR94), .A2(_02374__PTR126), .ZN(_00904__PTR1) );
  OR2_X1 U1846 ( .A1(_02374__PTR158), .A2(_02374__PTR190), .ZN(_00904__PTR2) );
  OR2_X1 U1847 ( .A1(_00904__PTR0), .A2(_00904__PTR1), .ZN(_00905__PTR0) );
  OR2_X1 U1848 ( .A1(_00904__PTR2), .A2(_02374__PTR222), .ZN(_00905__PTR1) );
  OR2_X1 U1849 ( .A1(_00905__PTR0), .A2(_00905__PTR1), .ZN(_02376__PTR30) );
  OR2_X1 U1850 ( .A1(_02374__PTR31), .A2(_02374__PTR63), .ZN(_00906__PTR0) );
  OR2_X1 U1851 ( .A1(_02374__PTR95), .A2(_02374__PTR127), .ZN(_00906__PTR1) );
  OR2_X1 U1852 ( .A1(_02374__PTR159), .A2(_02374__PTR191), .ZN(_00906__PTR2) );
  OR2_X1 U1853 ( .A1(_00906__PTR0), .A2(_00906__PTR1), .ZN(_00907__PTR0) );
  OR2_X1 U1854 ( .A1(_00906__PTR2), .A2(_02374__PTR223), .ZN(_00907__PTR1) );
  OR2_X1 U1855 ( .A1(_00907__PTR0), .A2(_00907__PTR1), .ZN(_02376__PTR31) );
  OR2_X1 U1856 ( .A1(_02375__PTR0), .A2(_02375__PTR1), .ZN(_00805__PTR0) );
  OR2_X1 U1857 ( .A1(_02148__PTR0), .A2(_02148__PTR1), .ZN(_00793__PTR0) );
  OR2_X1 U1858 ( .A1(_02375__PTR4), .A2(_02148__PTR2), .ZN(_02152__PTR2) );
  OR2_X1 U1859 ( .A1(_00805__PTR0), .A2(_00793__PTR0), .ZN(_00908__PTR0) );
  OR2_X1 U1860 ( .A1(_02152__PTR2), .A2(_02148__PTR3), .ZN(_00793__PTR1) );
  OR2_X1 U1861 ( .A1(_00908__PTR0), .A2(_00793__PTR1), .ZN(_03165_) );
  OR2_X1 U1862 ( .A1(_02382__PTR0), .A2(_02382__PTR32), .ZN(_00909_) );
  OR2_X1 U1863 ( .A1(_00909_), .A2(_02382__PTR64), .ZN(_02384__PTR0) );
  OR2_X1 U1864 ( .A1(_02382__PTR1), .A2(_02382__PTR33), .ZN(_00910_) );
  OR2_X1 U1865 ( .A1(_00910_), .A2(_02382__PTR65), .ZN(_02384__PTR1) );
  OR2_X1 U1866 ( .A1(_02382__PTR2), .A2(_02382__PTR34), .ZN(_00911_) );
  OR2_X1 U1867 ( .A1(_00911_), .A2(_02382__PTR66), .ZN(_02384__PTR2) );
  OR2_X1 U1868 ( .A1(_02382__PTR3), .A2(_02382__PTR35), .ZN(_00912_) );
  OR2_X1 U1869 ( .A1(_00912_), .A2(_02382__PTR67), .ZN(_02384__PTR3) );
  OR2_X1 U1870 ( .A1(_02382__PTR4), .A2(_02382__PTR36), .ZN(_00913_) );
  OR2_X1 U1871 ( .A1(_00913_), .A2(_02382__PTR68), .ZN(_02384__PTR4) );
  OR2_X1 U1872 ( .A1(_02382__PTR5), .A2(_02382__PTR37), .ZN(_00914_) );
  OR2_X1 U1873 ( .A1(_00914_), .A2(_02382__PTR69), .ZN(_02384__PTR5) );
  OR2_X1 U1874 ( .A1(_02382__PTR6), .A2(_02382__PTR38), .ZN(_00915_) );
  OR2_X1 U1875 ( .A1(_00915_), .A2(_02382__PTR70), .ZN(_02384__PTR6) );
  OR2_X1 U1876 ( .A1(_02382__PTR7), .A2(_02382__PTR39), .ZN(_00916_) );
  OR2_X1 U1877 ( .A1(_00916_), .A2(_02382__PTR71), .ZN(_02384__PTR7) );
  OR2_X1 U1878 ( .A1(_02382__PTR8), .A2(_02382__PTR40), .ZN(_00917_) );
  OR2_X1 U1879 ( .A1(_00917_), .A2(_02382__PTR72), .ZN(_02384__PTR8) );
  OR2_X1 U1880 ( .A1(_02382__PTR9), .A2(_02382__PTR41), .ZN(_00918_) );
  OR2_X1 U1881 ( .A1(_00918_), .A2(_02382__PTR73), .ZN(_02384__PTR9) );
  OR2_X1 U1882 ( .A1(_02382__PTR10), .A2(_02382__PTR42), .ZN(_00919_) );
  OR2_X1 U1883 ( .A1(_00919_), .A2(_02382__PTR74), .ZN(_02384__PTR10) );
  OR2_X1 U1884 ( .A1(_02382__PTR11), .A2(_02382__PTR43), .ZN(_00920_) );
  OR2_X1 U1885 ( .A1(_00920_), .A2(_02382__PTR75), .ZN(_02384__PTR11) );
  OR2_X1 U1886 ( .A1(_02382__PTR12), .A2(_02382__PTR44), .ZN(_00921_) );
  OR2_X1 U1887 ( .A1(_00921_), .A2(_02382__PTR76), .ZN(_02384__PTR12) );
  OR2_X1 U1888 ( .A1(_02382__PTR13), .A2(_02382__PTR45), .ZN(_00922_) );
  OR2_X1 U1889 ( .A1(_00922_), .A2(_02382__PTR77), .ZN(_02384__PTR13) );
  OR2_X1 U1890 ( .A1(_02382__PTR14), .A2(_02382__PTR46), .ZN(_00923_) );
  OR2_X1 U1891 ( .A1(_00923_), .A2(_02382__PTR78), .ZN(_02384__PTR14) );
  OR2_X1 U1892 ( .A1(_02382__PTR15), .A2(_02382__PTR47), .ZN(_00924_) );
  OR2_X1 U1893 ( .A1(_00924_), .A2(_02382__PTR79), .ZN(_02384__PTR15) );
  OR2_X1 U1894 ( .A1(_02382__PTR16), .A2(_02382__PTR48), .ZN(_00925_) );
  OR2_X1 U1895 ( .A1(_00925_), .A2(_02382__PTR80), .ZN(_02384__PTR16) );
  OR2_X1 U1896 ( .A1(_02382__PTR17), .A2(_02382__PTR49), .ZN(_00926_) );
  OR2_X1 U1897 ( .A1(_00926_), .A2(_02382__PTR81), .ZN(_02384__PTR17) );
  OR2_X1 U1898 ( .A1(_02382__PTR18), .A2(_02382__PTR50), .ZN(_00927_) );
  OR2_X1 U1899 ( .A1(_00927_), .A2(_02382__PTR82), .ZN(_02384__PTR18) );
  OR2_X1 U1900 ( .A1(_02382__PTR19), .A2(_02382__PTR51), .ZN(_00928_) );
  OR2_X1 U1901 ( .A1(_00928_), .A2(_02382__PTR83), .ZN(_02384__PTR19) );
  OR2_X1 U1902 ( .A1(_02382__PTR20), .A2(_02382__PTR52), .ZN(_00929_) );
  OR2_X1 U1903 ( .A1(_00929_), .A2(_02382__PTR84), .ZN(_02384__PTR20) );
  OR2_X1 U1904 ( .A1(_02382__PTR21), .A2(_02382__PTR53), .ZN(_00930_) );
  OR2_X1 U1905 ( .A1(_00930_), .A2(_02382__PTR85), .ZN(_02384__PTR21) );
  OR2_X1 U1906 ( .A1(_02382__PTR22), .A2(_02382__PTR54), .ZN(_00931_) );
  OR2_X1 U1907 ( .A1(_00931_), .A2(_02382__PTR86), .ZN(_02384__PTR22) );
  OR2_X1 U1908 ( .A1(_02382__PTR23), .A2(_02382__PTR55), .ZN(_00932_) );
  OR2_X1 U1909 ( .A1(_00932_), .A2(_02382__PTR87), .ZN(_02384__PTR23) );
  OR2_X1 U1910 ( .A1(_02382__PTR24), .A2(_02382__PTR56), .ZN(_00933_) );
  OR2_X1 U1911 ( .A1(_00933_), .A2(_02382__PTR88), .ZN(_02384__PTR24) );
  OR2_X1 U1912 ( .A1(_02382__PTR25), .A2(_02382__PTR57), .ZN(_00934_) );
  OR2_X1 U1913 ( .A1(_00934_), .A2(_02382__PTR89), .ZN(_02384__PTR25) );
  OR2_X1 U1914 ( .A1(_02382__PTR26), .A2(_02382__PTR58), .ZN(_00935_) );
  OR2_X1 U1915 ( .A1(_00935_), .A2(_02382__PTR90), .ZN(_02384__PTR26) );
  OR2_X1 U1916 ( .A1(_02382__PTR27), .A2(_02382__PTR59), .ZN(_00936_) );
  OR2_X1 U1917 ( .A1(_00936_), .A2(_02382__PTR91), .ZN(_02384__PTR27) );
  OR2_X1 U1918 ( .A1(_02382__PTR28), .A2(_02382__PTR60), .ZN(_00937_) );
  OR2_X1 U1919 ( .A1(_00937_), .A2(_02382__PTR92), .ZN(_02384__PTR28) );
  OR2_X1 U1920 ( .A1(_02382__PTR29), .A2(_02382__PTR61), .ZN(_00938_) );
  OR2_X1 U1921 ( .A1(_00938_), .A2(_02382__PTR93), .ZN(_02384__PTR29) );
  OR2_X1 U1922 ( .A1(_02382__PTR30), .A2(_02382__PTR62), .ZN(_00939_) );
  OR2_X1 U1923 ( .A1(_00939_), .A2(_02382__PTR94), .ZN(_02384__PTR30) );
  OR2_X1 U1924 ( .A1(_02382__PTR31), .A2(_02382__PTR63), .ZN(_00940_) );
  OR2_X1 U1925 ( .A1(_00940_), .A2(_02382__PTR95), .ZN(_02384__PTR31) );
  OR2_X1 U1926 ( .A1(_02383__PTR0), .A2(_02148__PTR2), .ZN(_00941_) );
  OR2_X1 U1927 ( .A1(_00941_), .A2(_02148__PTR3), .ZN(_03167_) );
  OR2_X1 U1928 ( .A1(_02997_), .A2(_02998_), .ZN(_01768__PTR2) );
  OR2_X1 U1929 ( .A1(_02408__PTR0), .A2(_02408__PTR4), .ZN(_02411__PTR0) );
  OR2_X1 U1930 ( .A1(_02408__PTR1), .A2(_02408__PTR5), .ZN(_02411__PTR1) );
  OR2_X1 U1931 ( .A1(_02408__PTR2), .A2(_02408__PTR6), .ZN(_02411__PTR2) );
  OR2_X1 U1932 ( .A1(_02408__PTR3), .A2(_02408__PTR7), .ZN(_02411__PTR3) );
  OR2_X1 U1933 ( .A1(_02409__PTR0), .A2(_02156__PTR2), .ZN(_03173_) );
  OR2_X1 U1934 ( .A1(_02975_), .A2(_02976_), .ZN(_02296_) );
  AND2_X1 U1935 ( .A1(_00942__PTR0), .A2(_02964__PTR3), .ZN(_00943_) );
  AND2_X1 U1936 ( .A1(_00943_), .A2(_00942__PTR2), .ZN(_02976_) );
  OR2_X1 U1937 ( .A1(_02972_), .A2(_02973_), .ZN(_02146__PTR2) );
  AND2_X1 U1938 ( .A1(_02962__PTR0), .A2(_02963__PTR1), .ZN(_00944__PTR0) );
  AND2_X1 U1939 ( .A1(_00944__PTR0), .A2(_00944__PTR1), .ZN(_00945_) );
  AND2_X1 U1940 ( .A1(_00945_), .A2(_00942__PTR2), .ZN(_02973_) );
  OR2_X1 U1941 ( .A1(_02966_), .A2(_02967_), .ZN(_02146__PTR3) );
  AND2_X1 U1942 ( .A1(_02962__PTR0), .A2(_02962__PTR1), .ZN(_00946__PTR0) );
  AND2_X1 U1943 ( .A1(_00946__PTR0), .A2(_02964__PTR3), .ZN(_00947_) );
  AND2_X1 U1944 ( .A1(_00947_), .A2(_00942__PTR2), .ZN(_02967_) );
  OR2_X1 U1945 ( .A1(_02701__PTR8), .A2(_02701__PTR12), .ZN(_00948__PTR1) );
  OR2_X1 U1946 ( .A1(_02701__PTR4), .A2(_00948__PTR1), .ZN(_02704__PTR0) );
  OR2_X1 U1947 ( .A1(_02701__PTR9), .A2(_02701__PTR13), .ZN(_00949__PTR1) );
  OR2_X1 U1948 ( .A1(_02701__PTR5), .A2(_00949__PTR1), .ZN(_02704__PTR1) );
  OR2_X1 U1949 ( .A1(_02701__PTR10), .A2(_02701__PTR14), .ZN(_00950__PTR1) );
  OR2_X1 U1950 ( .A1(_02701__PTR6), .A2(_00950__PTR1), .ZN(_02704__PTR2) );
  OR2_X1 U1951 ( .A1(_02701__PTR11), .A2(_02701__PTR15), .ZN(_02704__PTR3) );
  OR2_X1 U1952 ( .A1(_02702__PTR0), .A2(_02702__PTR1), .ZN(_00951__PTR0) );
  OR2_X1 U1953 ( .A1(_02702__PTR2), .A2(_02702__PTR3), .ZN(_00951__PTR1) );
  OR2_X1 U1954 ( .A1(_00951__PTR0), .A2(_00951__PTR1), .ZN(_03419_) );
  OR2_X1 U1955 ( .A1(_02693__PTR0), .A2(_02693__PTR32), .ZN(_00952_) );
  OR2_X1 U1956 ( .A1(_00952_), .A2(_02693__PTR64), .ZN(_02695__PTR0) );
  OR2_X1 U1957 ( .A1(_02693__PTR1), .A2(_02693__PTR33), .ZN(_00953_) );
  OR2_X1 U1958 ( .A1(_00953_), .A2(_02693__PTR65), .ZN(_02695__PTR1) );
  OR2_X1 U1959 ( .A1(_02693__PTR2), .A2(_02693__PTR34), .ZN(_00954_) );
  OR2_X1 U1960 ( .A1(_00954_), .A2(_02693__PTR66), .ZN(_02695__PTR2) );
  OR2_X1 U1961 ( .A1(_02693__PTR3), .A2(_02693__PTR35), .ZN(_00955_) );
  OR2_X1 U1962 ( .A1(_00955_), .A2(_02693__PTR67), .ZN(_02695__PTR3) );
  OR2_X1 U1963 ( .A1(_02693__PTR4), .A2(_02693__PTR36), .ZN(_00956_) );
  OR2_X1 U1964 ( .A1(_00956_), .A2(_02693__PTR68), .ZN(_02695__PTR4) );
  OR2_X1 U1965 ( .A1(_02693__PTR5), .A2(_02693__PTR37), .ZN(_00957_) );
  OR2_X1 U1966 ( .A1(_00957_), .A2(_02693__PTR69), .ZN(_02695__PTR5) );
  OR2_X1 U1967 ( .A1(_02693__PTR6), .A2(_02693__PTR38), .ZN(_00958_) );
  OR2_X1 U1968 ( .A1(_00958_), .A2(_02693__PTR70), .ZN(_02695__PTR6) );
  OR2_X1 U1969 ( .A1(_02693__PTR7), .A2(_02693__PTR39), .ZN(_00959_) );
  OR2_X1 U1970 ( .A1(_00959_), .A2(_02693__PTR71), .ZN(_02695__PTR7) );
  OR2_X1 U1971 ( .A1(_02693__PTR8), .A2(_02693__PTR40), .ZN(_00960_) );
  OR2_X1 U1972 ( .A1(_00960_), .A2(_02693__PTR72), .ZN(_02695__PTR8) );
  OR2_X1 U1973 ( .A1(_02693__PTR9), .A2(_02693__PTR41), .ZN(_00961_) );
  OR2_X1 U1974 ( .A1(_00961_), .A2(_02693__PTR73), .ZN(_02695__PTR9) );
  OR2_X1 U1975 ( .A1(_02693__PTR10), .A2(_02693__PTR42), .ZN(_00962_) );
  OR2_X1 U1976 ( .A1(_00962_), .A2(_02693__PTR74), .ZN(_02695__PTR10) );
  OR2_X1 U1977 ( .A1(_02693__PTR11), .A2(_02693__PTR43), .ZN(_00963_) );
  OR2_X1 U1978 ( .A1(_00963_), .A2(_02693__PTR75), .ZN(_02695__PTR11) );
  OR2_X1 U1979 ( .A1(_02693__PTR12), .A2(_02693__PTR44), .ZN(_00964_) );
  OR2_X1 U1980 ( .A1(_00964_), .A2(_02693__PTR76), .ZN(_02695__PTR12) );
  OR2_X1 U1981 ( .A1(_02693__PTR13), .A2(_02693__PTR45), .ZN(_00965_) );
  OR2_X1 U1982 ( .A1(_00965_), .A2(_02693__PTR77), .ZN(_02695__PTR13) );
  OR2_X1 U1983 ( .A1(_02693__PTR14), .A2(_02693__PTR46), .ZN(_00966_) );
  OR2_X1 U1984 ( .A1(_00966_), .A2(_02693__PTR78), .ZN(_02695__PTR14) );
  OR2_X1 U1985 ( .A1(_02693__PTR15), .A2(_02693__PTR47), .ZN(_00967_) );
  OR2_X1 U1986 ( .A1(_00967_), .A2(_02693__PTR79), .ZN(_02695__PTR15) );
  OR2_X1 U1987 ( .A1(_02693__PTR16), .A2(_02693__PTR48), .ZN(_00968_) );
  OR2_X1 U1988 ( .A1(_00968_), .A2(_02693__PTR80), .ZN(_02695__PTR16) );
  OR2_X1 U1989 ( .A1(_02693__PTR17), .A2(_02693__PTR49), .ZN(_00969_) );
  OR2_X1 U1990 ( .A1(_00969_), .A2(_02693__PTR81), .ZN(_02695__PTR17) );
  OR2_X1 U1991 ( .A1(_02693__PTR18), .A2(_02693__PTR50), .ZN(_00970_) );
  OR2_X1 U1992 ( .A1(_00970_), .A2(_02693__PTR82), .ZN(_02695__PTR18) );
  OR2_X1 U1993 ( .A1(_02693__PTR19), .A2(_02693__PTR51), .ZN(_00971_) );
  OR2_X1 U1994 ( .A1(_00971_), .A2(_02693__PTR83), .ZN(_02695__PTR19) );
  OR2_X1 U1995 ( .A1(_02693__PTR20), .A2(_02693__PTR52), .ZN(_00972_) );
  OR2_X1 U1996 ( .A1(_00972_), .A2(_02693__PTR84), .ZN(_02695__PTR20) );
  OR2_X1 U1997 ( .A1(_02693__PTR21), .A2(_02693__PTR53), .ZN(_00973_) );
  OR2_X1 U1998 ( .A1(_00973_), .A2(_02693__PTR85), .ZN(_02695__PTR21) );
  OR2_X1 U1999 ( .A1(_02693__PTR22), .A2(_02693__PTR54), .ZN(_00974_) );
  OR2_X1 U2000 ( .A1(_00974_), .A2(_02693__PTR86), .ZN(_02695__PTR22) );
  OR2_X1 U2001 ( .A1(_02693__PTR23), .A2(_02693__PTR55), .ZN(_00975_) );
  OR2_X1 U2002 ( .A1(_00975_), .A2(_02693__PTR87), .ZN(_02695__PTR23) );
  OR2_X1 U2003 ( .A1(_02693__PTR24), .A2(_02693__PTR56), .ZN(_00976_) );
  OR2_X1 U2004 ( .A1(_00976_), .A2(_02693__PTR88), .ZN(_02695__PTR24) );
  OR2_X1 U2005 ( .A1(_02693__PTR25), .A2(_02693__PTR57), .ZN(_00977_) );
  OR2_X1 U2006 ( .A1(_00977_), .A2(_02693__PTR89), .ZN(_02695__PTR25) );
  OR2_X1 U2007 ( .A1(_02693__PTR26), .A2(_02693__PTR58), .ZN(_00978_) );
  OR2_X1 U2008 ( .A1(_00978_), .A2(_02693__PTR90), .ZN(_02695__PTR26) );
  OR2_X1 U2009 ( .A1(_02693__PTR27), .A2(_02693__PTR59), .ZN(_00979_) );
  OR2_X1 U2010 ( .A1(_00979_), .A2(_02693__PTR91), .ZN(_02695__PTR27) );
  OR2_X1 U2011 ( .A1(_02693__PTR28), .A2(_02693__PTR60), .ZN(_00980_) );
  OR2_X1 U2012 ( .A1(_00980_), .A2(_02693__PTR92), .ZN(_02695__PTR28) );
  OR2_X1 U2013 ( .A1(_02693__PTR29), .A2(_02693__PTR61), .ZN(_00981_) );
  OR2_X1 U2014 ( .A1(_00981_), .A2(_02693__PTR93), .ZN(_02695__PTR29) );
  OR2_X1 U2015 ( .A1(_02693__PTR30), .A2(_02693__PTR62), .ZN(_00982_) );
  OR2_X1 U2016 ( .A1(_00982_), .A2(_02693__PTR94), .ZN(_02695__PTR30) );
  OR2_X1 U2017 ( .A1(_02693__PTR31), .A2(_02693__PTR63), .ZN(_00983_) );
  OR2_X1 U2018 ( .A1(_00983_), .A2(_02693__PTR95), .ZN(_02695__PTR31) );
  OR2_X1 U2019 ( .A1(_02694__PTR0), .A2(_02445__PTR0), .ZN(_00984_) );
  OR2_X1 U2020 ( .A1(_00984_), .A2(_02445__PTR2), .ZN(_03417_) );
  OR2_X1 U2021 ( .A1(_02690__PTR0), .A2(_02690__PTR16), .ZN(_00985_) );
  OR2_X1 U2022 ( .A1(_00985_), .A2(_02690__PTR32), .ZN(_02691__PTR0) );
  OR2_X1 U2023 ( .A1(_02690__PTR1), .A2(_02690__PTR17), .ZN(_00986_) );
  OR2_X1 U2024 ( .A1(_00986_), .A2(_02690__PTR33), .ZN(_02691__PTR1) );
  OR2_X1 U2025 ( .A1(_02690__PTR2), .A2(_02690__PTR18), .ZN(_00987_) );
  OR2_X1 U2026 ( .A1(_00987_), .A2(_02690__PTR34), .ZN(_02691__PTR2) );
  OR2_X1 U2027 ( .A1(_02690__PTR3), .A2(_02690__PTR19), .ZN(_00988_) );
  OR2_X1 U2028 ( .A1(_00988_), .A2(_02690__PTR35), .ZN(_02691__PTR3) );
  OR2_X1 U2029 ( .A1(_02690__PTR4), .A2(_02690__PTR20), .ZN(_00989_) );
  OR2_X1 U2030 ( .A1(_00989_), .A2(_02690__PTR36), .ZN(_02691__PTR4) );
  OR2_X1 U2031 ( .A1(_02690__PTR5), .A2(_02690__PTR21), .ZN(_00990_) );
  OR2_X1 U2032 ( .A1(_00990_), .A2(_02690__PTR37), .ZN(_02691__PTR5) );
  OR2_X1 U2033 ( .A1(_02690__PTR6), .A2(_02690__PTR22), .ZN(_00991_) );
  OR2_X1 U2034 ( .A1(_00991_), .A2(_02690__PTR38), .ZN(_02691__PTR6) );
  OR2_X1 U2035 ( .A1(_02690__PTR7), .A2(_02690__PTR23), .ZN(_00992_) );
  OR2_X1 U2036 ( .A1(_00992_), .A2(_02690__PTR39), .ZN(_02691__PTR7) );
  OR2_X1 U2037 ( .A1(_02690__PTR8), .A2(_02690__PTR24), .ZN(_00993_) );
  OR2_X1 U2038 ( .A1(_00993_), .A2(_02690__PTR40), .ZN(_02691__PTR8) );
  OR2_X1 U2039 ( .A1(_02690__PTR9), .A2(_02690__PTR25), .ZN(_00994_) );
  OR2_X1 U2040 ( .A1(_00994_), .A2(_02690__PTR41), .ZN(_02691__PTR9) );
  OR2_X1 U2041 ( .A1(_02690__PTR10), .A2(_02690__PTR26), .ZN(_00995_) );
  OR2_X1 U2042 ( .A1(_00995_), .A2(_02690__PTR42), .ZN(_02691__PTR10) );
  OR2_X1 U2043 ( .A1(_02690__PTR11), .A2(_02690__PTR27), .ZN(_00996_) );
  OR2_X1 U2044 ( .A1(_00996_), .A2(_02690__PTR43), .ZN(_02691__PTR11) );
  OR2_X1 U2045 ( .A1(_02690__PTR12), .A2(_02690__PTR28), .ZN(_00997_) );
  OR2_X1 U2046 ( .A1(_00997_), .A2(_02690__PTR44), .ZN(_02691__PTR12) );
  OR2_X1 U2047 ( .A1(_02690__PTR13), .A2(_02690__PTR29), .ZN(_00998_) );
  OR2_X1 U2048 ( .A1(_00998_), .A2(_02690__PTR45), .ZN(_02691__PTR13) );
  OR2_X1 U2049 ( .A1(_02690__PTR14), .A2(_02690__PTR30), .ZN(_00999_) );
  OR2_X1 U2050 ( .A1(_00999_), .A2(_02690__PTR46), .ZN(_02691__PTR14) );
  OR2_X1 U2051 ( .A1(_02690__PTR15), .A2(_02690__PTR31), .ZN(_01000_) );
  OR2_X1 U2052 ( .A1(_01000_), .A2(_02690__PTR47), .ZN(_02691__PTR15) );
  OR2_X1 U2053 ( .A1(_02686__PTR0), .A2(_02686__PTR15), .ZN(_01002_) );
  OR2_X1 U2054 ( .A1(_01002_), .A2(_02686__PTR30), .ZN(_02688__PTR0) );
  OR2_X1 U2055 ( .A1(_02686__PTR1), .A2(_02686__PTR16), .ZN(_01003_) );
  OR2_X1 U2056 ( .A1(_01003_), .A2(_02686__PTR31), .ZN(_02688__PTR1) );
  OR2_X1 U2057 ( .A1(_02686__PTR2), .A2(_02686__PTR17), .ZN(_01004_) );
  OR2_X1 U2058 ( .A1(_01004_), .A2(_02686__PTR32), .ZN(_02688__PTR2) );
  OR2_X1 U2059 ( .A1(_02686__PTR3), .A2(_02686__PTR18), .ZN(_01005_) );
  OR2_X1 U2060 ( .A1(_01005_), .A2(_02686__PTR33), .ZN(_02688__PTR3) );
  OR2_X1 U2061 ( .A1(_02686__PTR4), .A2(_02686__PTR19), .ZN(_01006_) );
  OR2_X1 U2062 ( .A1(_01006_), .A2(_02686__PTR34), .ZN(_02688__PTR4) );
  OR2_X1 U2063 ( .A1(_02686__PTR5), .A2(_02686__PTR20), .ZN(_01007_) );
  OR2_X1 U2064 ( .A1(_01007_), .A2(_02686__PTR35), .ZN(_02688__PTR5) );
  OR2_X1 U2065 ( .A1(_02686__PTR6), .A2(_02686__PTR21), .ZN(_01008_) );
  OR2_X1 U2066 ( .A1(_01008_), .A2(_02686__PTR36), .ZN(_02688__PTR6) );
  OR2_X1 U2067 ( .A1(_02686__PTR7), .A2(_02686__PTR22), .ZN(_01009_) );
  OR2_X1 U2068 ( .A1(_01009_), .A2(_02686__PTR37), .ZN(_02688__PTR7) );
  OR2_X1 U2069 ( .A1(_02686__PTR8), .A2(_02686__PTR23), .ZN(_01010_) );
  OR2_X1 U2070 ( .A1(_01010_), .A2(_02686__PTR38), .ZN(_02688__PTR8) );
  OR2_X1 U2071 ( .A1(_02686__PTR9), .A2(_02686__PTR24), .ZN(_01011_) );
  OR2_X1 U2072 ( .A1(_01011_), .A2(_02686__PTR39), .ZN(_02688__PTR9) );
  OR2_X1 U2073 ( .A1(_02686__PTR10), .A2(_02686__PTR25), .ZN(_01012_) );
  OR2_X1 U2074 ( .A1(_01012_), .A2(_02686__PTR40), .ZN(_02688__PTR10) );
  OR2_X1 U2075 ( .A1(_02686__PTR11), .A2(_02686__PTR26), .ZN(_01013_) );
  OR2_X1 U2076 ( .A1(_01013_), .A2(_02686__PTR41), .ZN(_02688__PTR11) );
  OR2_X1 U2077 ( .A1(_02686__PTR12), .A2(_02686__PTR27), .ZN(_01014_) );
  OR2_X1 U2078 ( .A1(_01014_), .A2(_02686__PTR42), .ZN(_02688__PTR12) );
  OR2_X1 U2079 ( .A1(_02686__PTR13), .A2(_02686__PTR28), .ZN(_01015_) );
  OR2_X1 U2080 ( .A1(_01015_), .A2(_02686__PTR43), .ZN(_02688__PTR13) );
  OR2_X1 U2081 ( .A1(_02686__PTR14), .A2(_02686__PTR29), .ZN(_01016_) );
  OR2_X1 U2082 ( .A1(_01016_), .A2(_02686__PTR44), .ZN(_02688__PTR14) );
  OR2_X1 U2083 ( .A1(_02687__PTR0), .A2(_02445__PTR2), .ZN(_01001_) );
  OR2_X1 U2084 ( .A1(_01001_), .A2(_02668__PTR4), .ZN(_03416_) );
  OR2_X1 U2085 ( .A1(_02679__PTR0), .A2(_02679__PTR32), .ZN(_01017_) );
  OR2_X1 U2086 ( .A1(_01017_), .A2(_02679__PTR64), .ZN(_02681__PTR0) );
  OR2_X1 U2087 ( .A1(_02679__PTR1), .A2(_02679__PTR33), .ZN(_01018_) );
  OR2_X1 U2088 ( .A1(_01018_), .A2(_02679__PTR65), .ZN(_02681__PTR1) );
  OR2_X1 U2089 ( .A1(_02679__PTR2), .A2(_02679__PTR34), .ZN(_01019_) );
  OR2_X1 U2090 ( .A1(_01019_), .A2(_02679__PTR66), .ZN(_02681__PTR2) );
  OR2_X1 U2091 ( .A1(_02679__PTR3), .A2(_02679__PTR35), .ZN(_01020_) );
  OR2_X1 U2092 ( .A1(_01020_), .A2(_02679__PTR67), .ZN(_02681__PTR3) );
  OR2_X1 U2093 ( .A1(_02679__PTR4), .A2(_02679__PTR36), .ZN(_01021_) );
  OR2_X1 U2094 ( .A1(_01021_), .A2(_02679__PTR68), .ZN(_02681__PTR4) );
  OR2_X1 U2095 ( .A1(_02679__PTR5), .A2(_02679__PTR37), .ZN(_01022_) );
  OR2_X1 U2096 ( .A1(_01022_), .A2(_02679__PTR69), .ZN(_02681__PTR5) );
  OR2_X1 U2097 ( .A1(_02679__PTR6), .A2(_02679__PTR38), .ZN(_01023_) );
  OR2_X1 U2098 ( .A1(_01023_), .A2(_02679__PTR70), .ZN(_02681__PTR6) );
  OR2_X1 U2099 ( .A1(_02679__PTR7), .A2(_02679__PTR39), .ZN(_01024_) );
  OR2_X1 U2100 ( .A1(_01024_), .A2(_02679__PTR71), .ZN(_02681__PTR7) );
  OR2_X1 U2101 ( .A1(_02679__PTR8), .A2(_02679__PTR40), .ZN(_01025_) );
  OR2_X1 U2102 ( .A1(_01025_), .A2(_02679__PTR72), .ZN(_02681__PTR8) );
  OR2_X1 U2103 ( .A1(_02679__PTR9), .A2(_02679__PTR41), .ZN(_01026_) );
  OR2_X1 U2104 ( .A1(_01026_), .A2(_02679__PTR73), .ZN(_02681__PTR9) );
  OR2_X1 U2105 ( .A1(_02679__PTR10), .A2(_02679__PTR42), .ZN(_01027_) );
  OR2_X1 U2106 ( .A1(_01027_), .A2(_02679__PTR74), .ZN(_02681__PTR10) );
  OR2_X1 U2107 ( .A1(_02679__PTR11), .A2(_02679__PTR43), .ZN(_01028_) );
  OR2_X1 U2108 ( .A1(_01028_), .A2(_02679__PTR75), .ZN(_02681__PTR11) );
  OR2_X1 U2109 ( .A1(_02679__PTR12), .A2(_02679__PTR44), .ZN(_01029_) );
  OR2_X1 U2110 ( .A1(_01029_), .A2(_02679__PTR76), .ZN(_02681__PTR12) );
  OR2_X1 U2111 ( .A1(_02679__PTR13), .A2(_02679__PTR45), .ZN(_01030_) );
  OR2_X1 U2112 ( .A1(_01030_), .A2(_02679__PTR77), .ZN(_02681__PTR13) );
  OR2_X1 U2113 ( .A1(_02679__PTR14), .A2(_02679__PTR46), .ZN(_01031_) );
  OR2_X1 U2114 ( .A1(_01031_), .A2(_02679__PTR78), .ZN(_02681__PTR14) );
  OR2_X1 U2115 ( .A1(_02679__PTR15), .A2(_02679__PTR47), .ZN(_01032_) );
  OR2_X1 U2116 ( .A1(_01032_), .A2(_02679__PTR79), .ZN(_02681__PTR15) );
  OR2_X1 U2117 ( .A1(_02679__PTR16), .A2(_02679__PTR48), .ZN(_01033_) );
  OR2_X1 U2118 ( .A1(_01033_), .A2(_02679__PTR80), .ZN(_02681__PTR16) );
  OR2_X1 U2119 ( .A1(_02679__PTR17), .A2(_02679__PTR49), .ZN(_01034_) );
  OR2_X1 U2120 ( .A1(_01034_), .A2(_02679__PTR81), .ZN(_02681__PTR17) );
  OR2_X1 U2121 ( .A1(_02679__PTR18), .A2(_02679__PTR50), .ZN(_01035_) );
  OR2_X1 U2122 ( .A1(_01035_), .A2(_02679__PTR82), .ZN(_02681__PTR18) );
  OR2_X1 U2123 ( .A1(_02679__PTR19), .A2(_02679__PTR51), .ZN(_01036_) );
  OR2_X1 U2124 ( .A1(_01036_), .A2(_02679__PTR83), .ZN(_02681__PTR19) );
  OR2_X1 U2125 ( .A1(_02679__PTR20), .A2(_02679__PTR52), .ZN(_01037_) );
  OR2_X1 U2126 ( .A1(_01037_), .A2(_02679__PTR84), .ZN(_02681__PTR20) );
  OR2_X1 U2127 ( .A1(_02679__PTR21), .A2(_02679__PTR53), .ZN(_01038_) );
  OR2_X1 U2128 ( .A1(_01038_), .A2(_02679__PTR85), .ZN(_02681__PTR21) );
  OR2_X1 U2129 ( .A1(_02679__PTR22), .A2(_02679__PTR54), .ZN(_01039_) );
  OR2_X1 U2130 ( .A1(_01039_), .A2(_02679__PTR86), .ZN(_02681__PTR22) );
  OR2_X1 U2131 ( .A1(_02679__PTR23), .A2(_02679__PTR55), .ZN(_01040_) );
  OR2_X1 U2132 ( .A1(_01040_), .A2(_02679__PTR87), .ZN(_02681__PTR23) );
  OR2_X1 U2133 ( .A1(_02679__PTR24), .A2(_02679__PTR56), .ZN(_01041_) );
  OR2_X1 U2134 ( .A1(_01041_), .A2(_02679__PTR88), .ZN(_02681__PTR24) );
  OR2_X1 U2135 ( .A1(_02679__PTR25), .A2(_02679__PTR57), .ZN(_01042_) );
  OR2_X1 U2136 ( .A1(_01042_), .A2(_02679__PTR89), .ZN(_02681__PTR25) );
  OR2_X1 U2137 ( .A1(_02679__PTR26), .A2(_02679__PTR58), .ZN(_01043_) );
  OR2_X1 U2138 ( .A1(_01043_), .A2(_02679__PTR90), .ZN(_02681__PTR26) );
  OR2_X1 U2139 ( .A1(_02679__PTR27), .A2(_02679__PTR59), .ZN(_01044_) );
  OR2_X1 U2140 ( .A1(_01044_), .A2(_02679__PTR91), .ZN(_02681__PTR27) );
  OR2_X1 U2141 ( .A1(_02679__PTR28), .A2(_02679__PTR60), .ZN(_01045_) );
  OR2_X1 U2142 ( .A1(_01045_), .A2(_02679__PTR92), .ZN(_02681__PTR28) );
  OR2_X1 U2143 ( .A1(_02679__PTR29), .A2(_02679__PTR61), .ZN(_01046_) );
  OR2_X1 U2144 ( .A1(_01046_), .A2(_02679__PTR93), .ZN(_02681__PTR29) );
  OR2_X1 U2145 ( .A1(_02679__PTR30), .A2(_02679__PTR62), .ZN(_01047_) );
  OR2_X1 U2146 ( .A1(_01047_), .A2(_02679__PTR94), .ZN(_02681__PTR30) );
  OR2_X1 U2147 ( .A1(_02679__PTR31), .A2(_02679__PTR63), .ZN(_01048_) );
  OR2_X1 U2148 ( .A1(_01048_), .A2(_02679__PTR95), .ZN(_02681__PTR31) );
  OR2_X1 U2149 ( .A1(_02680__PTR0), .A2(_02680__PTR1), .ZN(_01049_) );
  OR2_X1 U2150 ( .A1(_01049_), .A2(_02680__PTR2), .ZN(_03414_) );
  OR2_X1 U2151 ( .A1(_02675__PTR0), .A2(_02675__PTR32), .ZN(_01050__PTR0) );
  OR2_X1 U2152 ( .A1(_02675__PTR64), .A2(_02675__PTR96), .ZN(_01050__PTR1) );
  OR2_X1 U2153 ( .A1(_01050__PTR0), .A2(_01050__PTR1), .ZN(_01051_) );
  OR2_X1 U2154 ( .A1(_01051_), .A2(_02675__PTR128), .ZN(_02677__PTR0) );
  OR2_X1 U2155 ( .A1(_02675__PTR1), .A2(_02675__PTR33), .ZN(_01052__PTR0) );
  OR2_X1 U2156 ( .A1(_02675__PTR65), .A2(_02675__PTR97), .ZN(_01052__PTR1) );
  OR2_X1 U2157 ( .A1(_01052__PTR0), .A2(_01052__PTR1), .ZN(_01053_) );
  OR2_X1 U2158 ( .A1(_01053_), .A2(_02675__PTR129), .ZN(_02677__PTR1) );
  OR2_X1 U2159 ( .A1(_02675__PTR2), .A2(_02675__PTR34), .ZN(_01054__PTR0) );
  OR2_X1 U2160 ( .A1(_02675__PTR66), .A2(_02675__PTR98), .ZN(_01054__PTR1) );
  OR2_X1 U2161 ( .A1(_01054__PTR0), .A2(_01054__PTR1), .ZN(_01055_) );
  OR2_X1 U2162 ( .A1(_01055_), .A2(_02675__PTR130), .ZN(_02677__PTR2) );
  OR2_X1 U2163 ( .A1(_02675__PTR3), .A2(_02675__PTR35), .ZN(_01056__PTR0) );
  OR2_X1 U2164 ( .A1(_02675__PTR67), .A2(_02675__PTR99), .ZN(_01056__PTR1) );
  OR2_X1 U2165 ( .A1(_01056__PTR0), .A2(_01056__PTR1), .ZN(_01057_) );
  OR2_X1 U2166 ( .A1(_01057_), .A2(_02675__PTR131), .ZN(_02677__PTR3) );
  OR2_X1 U2167 ( .A1(_02675__PTR4), .A2(_02675__PTR36), .ZN(_01058__PTR0) );
  OR2_X1 U2168 ( .A1(_02675__PTR68), .A2(_02675__PTR100), .ZN(_01058__PTR1) );
  OR2_X1 U2169 ( .A1(_01058__PTR0), .A2(_01058__PTR1), .ZN(_01059_) );
  OR2_X1 U2170 ( .A1(_01059_), .A2(_02675__PTR132), .ZN(_02677__PTR4) );
  OR2_X1 U2171 ( .A1(_02675__PTR5), .A2(_02675__PTR37), .ZN(_01060__PTR0) );
  OR2_X1 U2172 ( .A1(_02675__PTR69), .A2(_02675__PTR101), .ZN(_01060__PTR1) );
  OR2_X1 U2173 ( .A1(_01060__PTR0), .A2(_01060__PTR1), .ZN(_01061_) );
  OR2_X1 U2174 ( .A1(_01061_), .A2(_02675__PTR133), .ZN(_02677__PTR5) );
  OR2_X1 U2175 ( .A1(_02675__PTR6), .A2(_02675__PTR38), .ZN(_01062__PTR0) );
  OR2_X1 U2176 ( .A1(_02675__PTR70), .A2(_02675__PTR102), .ZN(_01062__PTR1) );
  OR2_X1 U2177 ( .A1(_01062__PTR0), .A2(_01062__PTR1), .ZN(_01063_) );
  OR2_X1 U2178 ( .A1(_01063_), .A2(_02675__PTR134), .ZN(_02677__PTR6) );
  OR2_X1 U2179 ( .A1(_02675__PTR7), .A2(_02675__PTR39), .ZN(_01064__PTR0) );
  OR2_X1 U2180 ( .A1(_02675__PTR71), .A2(_02675__PTR103), .ZN(_01064__PTR1) );
  OR2_X1 U2181 ( .A1(_01064__PTR0), .A2(_01064__PTR1), .ZN(_01065_) );
  OR2_X1 U2182 ( .A1(_01065_), .A2(_02675__PTR135), .ZN(_02677__PTR7) );
  OR2_X1 U2183 ( .A1(_02675__PTR8), .A2(_02675__PTR40), .ZN(_01066__PTR0) );
  OR2_X1 U2184 ( .A1(_02675__PTR72), .A2(_02675__PTR104), .ZN(_01066__PTR1) );
  OR2_X1 U2185 ( .A1(_01066__PTR0), .A2(_01066__PTR1), .ZN(_01067_) );
  OR2_X1 U2186 ( .A1(_01067_), .A2(_02675__PTR136), .ZN(_02677__PTR8) );
  OR2_X1 U2187 ( .A1(_02675__PTR9), .A2(_02675__PTR41), .ZN(_01068__PTR0) );
  OR2_X1 U2188 ( .A1(_02675__PTR73), .A2(_02675__PTR105), .ZN(_01068__PTR1) );
  OR2_X1 U2189 ( .A1(_01068__PTR0), .A2(_01068__PTR1), .ZN(_01069_) );
  OR2_X1 U2190 ( .A1(_01069_), .A2(_02675__PTR137), .ZN(_02677__PTR9) );
  OR2_X1 U2191 ( .A1(_02675__PTR10), .A2(_02675__PTR42), .ZN(_01070__PTR0) );
  OR2_X1 U2192 ( .A1(_02675__PTR74), .A2(_02675__PTR106), .ZN(_01070__PTR1) );
  OR2_X1 U2193 ( .A1(_01070__PTR0), .A2(_01070__PTR1), .ZN(_01071_) );
  OR2_X1 U2194 ( .A1(_01071_), .A2(_02675__PTR138), .ZN(_02677__PTR10) );
  OR2_X1 U2195 ( .A1(_02675__PTR11), .A2(_02675__PTR43), .ZN(_01072__PTR0) );
  OR2_X1 U2196 ( .A1(_02675__PTR75), .A2(_02675__PTR107), .ZN(_01072__PTR1) );
  OR2_X1 U2197 ( .A1(_01072__PTR0), .A2(_01072__PTR1), .ZN(_01073_) );
  OR2_X1 U2198 ( .A1(_01073_), .A2(_02675__PTR139), .ZN(_02677__PTR11) );
  OR2_X1 U2199 ( .A1(_02675__PTR12), .A2(_02675__PTR44), .ZN(_01074__PTR0) );
  OR2_X1 U2200 ( .A1(_02675__PTR76), .A2(_02675__PTR108), .ZN(_01074__PTR1) );
  OR2_X1 U2201 ( .A1(_01074__PTR0), .A2(_01074__PTR1), .ZN(_01075_) );
  OR2_X1 U2202 ( .A1(_01075_), .A2(_02675__PTR140), .ZN(_02677__PTR12) );
  OR2_X1 U2203 ( .A1(_02675__PTR13), .A2(_02675__PTR45), .ZN(_01076__PTR0) );
  OR2_X1 U2204 ( .A1(_02675__PTR77), .A2(_02675__PTR109), .ZN(_01076__PTR1) );
  OR2_X1 U2205 ( .A1(_01076__PTR0), .A2(_01076__PTR1), .ZN(_01077_) );
  OR2_X1 U2206 ( .A1(_01077_), .A2(_02675__PTR141), .ZN(_02677__PTR13) );
  OR2_X1 U2207 ( .A1(_02675__PTR14), .A2(_02675__PTR46), .ZN(_01078__PTR0) );
  OR2_X1 U2208 ( .A1(_02675__PTR78), .A2(_02675__PTR110), .ZN(_01078__PTR1) );
  OR2_X1 U2209 ( .A1(_01078__PTR0), .A2(_01078__PTR1), .ZN(_01079_) );
  OR2_X1 U2210 ( .A1(_01079_), .A2(_02675__PTR142), .ZN(_02677__PTR14) );
  OR2_X1 U2211 ( .A1(_02675__PTR15), .A2(_02675__PTR47), .ZN(_01080__PTR0) );
  OR2_X1 U2212 ( .A1(_02675__PTR79), .A2(_02675__PTR111), .ZN(_01080__PTR1) );
  OR2_X1 U2213 ( .A1(_01080__PTR0), .A2(_01080__PTR1), .ZN(_01081_) );
  OR2_X1 U2214 ( .A1(_01081_), .A2(_02675__PTR143), .ZN(_02677__PTR15) );
  OR2_X1 U2215 ( .A1(_02675__PTR16), .A2(_02675__PTR48), .ZN(_01082__PTR0) );
  OR2_X1 U2216 ( .A1(_02675__PTR80), .A2(_02675__PTR112), .ZN(_01082__PTR1) );
  OR2_X1 U2217 ( .A1(_01082__PTR0), .A2(_01082__PTR1), .ZN(_01083_) );
  OR2_X1 U2218 ( .A1(_01083_), .A2(_02675__PTR144), .ZN(_02677__PTR16) );
  OR2_X1 U2219 ( .A1(_02675__PTR17), .A2(_02675__PTR49), .ZN(_01084__PTR0) );
  OR2_X1 U2220 ( .A1(_02675__PTR81), .A2(_02675__PTR113), .ZN(_01084__PTR1) );
  OR2_X1 U2221 ( .A1(_01084__PTR0), .A2(_01084__PTR1), .ZN(_01085_) );
  OR2_X1 U2222 ( .A1(_01085_), .A2(_02675__PTR145), .ZN(_02677__PTR17) );
  OR2_X1 U2223 ( .A1(_02675__PTR18), .A2(_02675__PTR50), .ZN(_01086__PTR0) );
  OR2_X1 U2224 ( .A1(_02675__PTR82), .A2(_02675__PTR114), .ZN(_01086__PTR1) );
  OR2_X1 U2225 ( .A1(_01086__PTR0), .A2(_01086__PTR1), .ZN(_01087_) );
  OR2_X1 U2226 ( .A1(_01087_), .A2(_02675__PTR146), .ZN(_02677__PTR18) );
  OR2_X1 U2227 ( .A1(_02675__PTR19), .A2(_02675__PTR51), .ZN(_01088__PTR0) );
  OR2_X1 U2228 ( .A1(_02675__PTR83), .A2(_02675__PTR115), .ZN(_01088__PTR1) );
  OR2_X1 U2229 ( .A1(_01088__PTR0), .A2(_01088__PTR1), .ZN(_01089_) );
  OR2_X1 U2230 ( .A1(_01089_), .A2(_02675__PTR147), .ZN(_02677__PTR19) );
  OR2_X1 U2231 ( .A1(_02675__PTR20), .A2(_02675__PTR52), .ZN(_01090__PTR0) );
  OR2_X1 U2232 ( .A1(_02675__PTR84), .A2(_02675__PTR116), .ZN(_01090__PTR1) );
  OR2_X1 U2233 ( .A1(_01090__PTR0), .A2(_01090__PTR1), .ZN(_01091_) );
  OR2_X1 U2234 ( .A1(_01091_), .A2(_02675__PTR148), .ZN(_02677__PTR20) );
  OR2_X1 U2235 ( .A1(_02675__PTR21), .A2(_02675__PTR53), .ZN(_01092__PTR0) );
  OR2_X1 U2236 ( .A1(_02675__PTR85), .A2(_02675__PTR117), .ZN(_01092__PTR1) );
  OR2_X1 U2237 ( .A1(_01092__PTR0), .A2(_01092__PTR1), .ZN(_01093_) );
  OR2_X1 U2238 ( .A1(_01093_), .A2(_02675__PTR149), .ZN(_02677__PTR21) );
  OR2_X1 U2239 ( .A1(_02675__PTR22), .A2(_02675__PTR54), .ZN(_01094__PTR0) );
  OR2_X1 U2240 ( .A1(_02675__PTR86), .A2(_02675__PTR118), .ZN(_01094__PTR1) );
  OR2_X1 U2241 ( .A1(_01094__PTR0), .A2(_01094__PTR1), .ZN(_01095_) );
  OR2_X1 U2242 ( .A1(_01095_), .A2(_02675__PTR150), .ZN(_02677__PTR22) );
  OR2_X1 U2243 ( .A1(_02675__PTR23), .A2(_02675__PTR55), .ZN(_01096__PTR0) );
  OR2_X1 U2244 ( .A1(_02675__PTR87), .A2(_02675__PTR119), .ZN(_01096__PTR1) );
  OR2_X1 U2245 ( .A1(_01096__PTR0), .A2(_01096__PTR1), .ZN(_01097_) );
  OR2_X1 U2246 ( .A1(_01097_), .A2(_02675__PTR151), .ZN(_02677__PTR23) );
  OR2_X1 U2247 ( .A1(_02675__PTR24), .A2(_02675__PTR56), .ZN(_01098__PTR0) );
  OR2_X1 U2248 ( .A1(_02675__PTR88), .A2(_02675__PTR120), .ZN(_01098__PTR1) );
  OR2_X1 U2249 ( .A1(_01098__PTR0), .A2(_01098__PTR1), .ZN(_01099_) );
  OR2_X1 U2250 ( .A1(_01099_), .A2(_02675__PTR152), .ZN(_02677__PTR24) );
  OR2_X1 U2251 ( .A1(_02675__PTR25), .A2(_02675__PTR57), .ZN(_01100__PTR0) );
  OR2_X1 U2252 ( .A1(_02675__PTR89), .A2(_02675__PTR121), .ZN(_01100__PTR1) );
  OR2_X1 U2253 ( .A1(_01100__PTR0), .A2(_01100__PTR1), .ZN(_01101_) );
  OR2_X1 U2254 ( .A1(_01101_), .A2(_02675__PTR153), .ZN(_02677__PTR25) );
  OR2_X1 U2255 ( .A1(_02675__PTR26), .A2(_02675__PTR58), .ZN(_01102__PTR0) );
  OR2_X1 U2256 ( .A1(_02675__PTR90), .A2(_02675__PTR122), .ZN(_01102__PTR1) );
  OR2_X1 U2257 ( .A1(_01102__PTR0), .A2(_01102__PTR1), .ZN(_01103_) );
  OR2_X1 U2258 ( .A1(_01103_), .A2(_02675__PTR154), .ZN(_02677__PTR26) );
  OR2_X1 U2259 ( .A1(_02675__PTR27), .A2(_02675__PTR59), .ZN(_01104__PTR0) );
  OR2_X1 U2260 ( .A1(_02675__PTR91), .A2(_02675__PTR123), .ZN(_01104__PTR1) );
  OR2_X1 U2261 ( .A1(_01104__PTR0), .A2(_01104__PTR1), .ZN(_01105_) );
  OR2_X1 U2262 ( .A1(_01105_), .A2(_02675__PTR155), .ZN(_02677__PTR27) );
  OR2_X1 U2263 ( .A1(_02675__PTR28), .A2(_02675__PTR60), .ZN(_01106__PTR0) );
  OR2_X1 U2264 ( .A1(_02675__PTR92), .A2(_02675__PTR124), .ZN(_01106__PTR1) );
  OR2_X1 U2265 ( .A1(_01106__PTR0), .A2(_01106__PTR1), .ZN(_01107_) );
  OR2_X1 U2266 ( .A1(_01107_), .A2(_02675__PTR156), .ZN(_02677__PTR28) );
  OR2_X1 U2267 ( .A1(_02675__PTR29), .A2(_02675__PTR61), .ZN(_01108__PTR0) );
  OR2_X1 U2268 ( .A1(_02675__PTR93), .A2(_02675__PTR125), .ZN(_01108__PTR1) );
  OR2_X1 U2269 ( .A1(_01108__PTR0), .A2(_01108__PTR1), .ZN(_01109_) );
  OR2_X1 U2270 ( .A1(_01109_), .A2(_02675__PTR157), .ZN(_02677__PTR29) );
  OR2_X1 U2271 ( .A1(_02675__PTR30), .A2(_02675__PTR62), .ZN(_01110__PTR0) );
  OR2_X1 U2272 ( .A1(_02675__PTR94), .A2(_02675__PTR126), .ZN(_01110__PTR1) );
  OR2_X1 U2273 ( .A1(_01110__PTR0), .A2(_01110__PTR1), .ZN(_01111_) );
  OR2_X1 U2274 ( .A1(_01111_), .A2(_02675__PTR158), .ZN(_02677__PTR30) );
  OR2_X1 U2275 ( .A1(_02675__PTR31), .A2(_02675__PTR63), .ZN(_01112__PTR0) );
  OR2_X1 U2276 ( .A1(_02675__PTR95), .A2(_02675__PTR127), .ZN(_01112__PTR1) );
  OR2_X1 U2277 ( .A1(_01112__PTR0), .A2(_01112__PTR1), .ZN(_01113_) );
  OR2_X1 U2278 ( .A1(_01113_), .A2(_02675__PTR159), .ZN(_02677__PTR31) );
  OR2_X1 U2279 ( .A1(_02676__PTR0), .A2(_02676__PTR1), .ZN(_01114__PTR0) );
  OR2_X1 U2280 ( .A1(_02668__PTR3), .A2(_02668__PTR4), .ZN(_02437__PTR1) );
  OR2_X1 U2281 ( .A1(_01114__PTR0), .A2(_02437__PTR1), .ZN(_01115_) );
  OR2_X1 U2282 ( .A1(_01115_), .A2(_02676__PTR4), .ZN(_03413_) );
  OR2_X1 U2283 ( .A1(_02440__PTR0), .A2(_02440__PTR1), .ZN(_01116__PTR0) );
  OR2_X1 U2284 ( .A1(_02440__PTR2), .A2(_02440__PTR3), .ZN(_01116__PTR1) );
  OR2_X1 U2285 ( .A1(_01116__PTR0), .A2(_01116__PTR1), .ZN(_02442_) );
  OR2_X1 U2286 ( .A1(_01117__PTR0), .A2(_01117__PTR1), .ZN(_03263_) );
  OR2_X1 U2287 ( .A1(_02436__PTR0), .A2(_02436__PTR1), .ZN(_01118__PTR0) );
  OR2_X1 U2288 ( .A1(_02436__PTR2), .A2(_02436__PTR3), .ZN(_01118__PTR1) );
  OR2_X1 U2289 ( .A1(_01118__PTR0), .A2(_01118__PTR1), .ZN(_02438_) );
  OR2_X1 U2290 ( .A1(_02437__PTR2), .A2(_02437__PTR3), .ZN(_02668__PTR6) );
  OR2_X1 U2291 ( .A1(_01117__PTR0), .A2(_02668__PTR6), .ZN(_03262_) );
  OR2_X1 U2292 ( .A1(_02667__PTR0), .A2(_02667__PTR5), .ZN(_01119__PTR0) );
  OR2_X1 U2293 ( .A1(_02667__PTR10), .A2(_02667__PTR15), .ZN(_01119__PTR1) );
  OR2_X1 U2294 ( .A1(_02667__PTR20), .A2(_02667__PTR25), .ZN(_01119__PTR2) );
  OR2_X1 U2295 ( .A1(_01119__PTR0), .A2(_01119__PTR1), .ZN(_01120__PTR0) );
  OR2_X1 U2296 ( .A1(_01119__PTR2), .A2(_02667__PTR30), .ZN(_01120__PTR1) );
  OR2_X1 U2297 ( .A1(_01120__PTR0), .A2(_01120__PTR1), .ZN(_02669__PTR0) );
  OR2_X1 U2298 ( .A1(_02667__PTR1), .A2(_02667__PTR6), .ZN(_01121__PTR0) );
  OR2_X1 U2299 ( .A1(_02667__PTR11), .A2(_02667__PTR16), .ZN(_01121__PTR1) );
  OR2_X1 U2300 ( .A1(_02667__PTR21), .A2(_02667__PTR26), .ZN(_01121__PTR2) );
  OR2_X1 U2301 ( .A1(_01121__PTR0), .A2(_01121__PTR1), .ZN(_01122__PTR0) );
  OR2_X1 U2302 ( .A1(_01121__PTR2), .A2(_02667__PTR31), .ZN(_01122__PTR1) );
  OR2_X1 U2303 ( .A1(_01122__PTR0), .A2(_01122__PTR1), .ZN(_02669__PTR1) );
  OR2_X1 U2304 ( .A1(_02667__PTR2), .A2(_02667__PTR7), .ZN(_01123__PTR0) );
  OR2_X1 U2305 ( .A1(_02667__PTR12), .A2(_02667__PTR17), .ZN(_01123__PTR1) );
  OR2_X1 U2306 ( .A1(_02667__PTR22), .A2(_02667__PTR27), .ZN(_01123__PTR2) );
  OR2_X1 U2307 ( .A1(_01123__PTR0), .A2(_01123__PTR1), .ZN(_01124__PTR0) );
  OR2_X1 U2308 ( .A1(_01123__PTR2), .A2(_02667__PTR32), .ZN(_01124__PTR1) );
  OR2_X1 U2309 ( .A1(_01124__PTR0), .A2(_01124__PTR1), .ZN(_02669__PTR2) );
  OR2_X1 U2310 ( .A1(_02667__PTR3), .A2(_02667__PTR8), .ZN(_01125__PTR0) );
  OR2_X1 U2311 ( .A1(_02667__PTR13), .A2(_02667__PTR18), .ZN(_01125__PTR1) );
  OR2_X1 U2312 ( .A1(_02667__PTR23), .A2(_02667__PTR28), .ZN(_01125__PTR2) );
  OR2_X1 U2313 ( .A1(_01125__PTR0), .A2(_01125__PTR1), .ZN(_01126__PTR0) );
  OR2_X1 U2314 ( .A1(_01125__PTR2), .A2(_02667__PTR33), .ZN(_01126__PTR1) );
  OR2_X1 U2315 ( .A1(_01126__PTR0), .A2(_01126__PTR1), .ZN(_02669__PTR3) );
  OR2_X1 U2316 ( .A1(_02667__PTR14), .A2(_02667__PTR19), .ZN(_01127__PTR1) );
  OR2_X1 U2317 ( .A1(_02667__PTR24), .A2(_02667__PTR29), .ZN(_01127__PTR2) );
  OR2_X1 U2318 ( .A1(_01127__PTR2), .A2(_02667__PTR34), .ZN(_01128__PTR1) );
  OR2_X1 U2319 ( .A1(_01127__PTR1), .A2(_01128__PTR1), .ZN(_02669__PTR4) );
  OR2_X1 U2320 ( .A1(_02437__PTR0), .A2(_02668__PTR3), .ZN(_01129__PTR1) );
  OR2_X1 U2321 ( .A1(_02668__PTR4), .A2(_02664__PTR4), .ZN(_01129__PTR2) );
  OR2_X1 U2322 ( .A1(_01129__PTR0), .A2(_01129__PTR1), .ZN(_01130__PTR0) );
  OR2_X1 U2323 ( .A1(_01129__PTR2), .A2(_02668__PTR6), .ZN(_01130__PTR1) );
  OR2_X1 U2324 ( .A1(_01130__PTR0), .A2(_01130__PTR1), .ZN(_03411_) );
  OR2_X1 U2325 ( .A1(_02455__PTR0), .A2(_02455__PTR1), .ZN(_02457_) );
  OR2_X1 U2326 ( .A1(_02444__PTR0), .A2(_02444__PTR1), .ZN(_01131__PTR0) );
  OR2_X1 U2327 ( .A1(_02444__PTR2), .A2(_02444__PTR3), .ZN(_01131__PTR1) );
  OR2_X1 U2328 ( .A1(_01131__PTR0), .A2(_01131__PTR1), .ZN(_02446_) );
  OR2_X1 U2329 ( .A1(_02445__PTR0), .A2(_02437__PTR1), .ZN(_01132__PTR0) );
  OR2_X1 U2330 ( .A1(_02445__PTR2), .A2(_02445__PTR3), .ZN(_01132__PTR1) );
  OR2_X1 U2331 ( .A1(_01132__PTR0), .A2(_01132__PTR1), .ZN(_03264_) );
  OR2_X1 U2332 ( .A1(_02451__PTR0), .A2(_02451__PTR1), .ZN(_01133_) );
  OR2_X1 U2333 ( .A1(_01133_), .A2(_02451__PTR2), .ZN(_02453_) );
  OR2_X1 U2334 ( .A1(_02452__PTR0), .A2(_02452__PTR1), .ZN(_02456__PTR0) );
  OR2_X1 U2335 ( .A1(_02456__PTR0), .A2(_02445__PTR3), .ZN(_03266_) );
  OR2_X1 U2336 ( .A1(_02448__PTR0), .A2(_02448__PTR1), .ZN(_01134_) );
  OR2_X1 U2337 ( .A1(_01134_), .A2(_02448__PTR2), .ZN(_02449_) );
  OR2_X1 U2338 ( .A1(_01117__PTR0), .A2(_02445__PTR3), .ZN(_03265_) );
  OR2_X1 U2339 ( .A1(_02683__PTR0), .A2(_02683__PTR32), .ZN(_01135__PTR0) );
  OR2_X1 U2340 ( .A1(_02683__PTR64), .A2(_02683__PTR96), .ZN(_01135__PTR1) );
  OR2_X1 U2341 ( .A1(_01135__PTR0), .A2(_01135__PTR1), .ZN(_02684__PTR0) );
  OR2_X1 U2342 ( .A1(_02683__PTR1), .A2(_02683__PTR33), .ZN(_01136__PTR0) );
  OR2_X1 U2343 ( .A1(_02683__PTR65), .A2(_02683__PTR97), .ZN(_01136__PTR1) );
  OR2_X1 U2344 ( .A1(_01136__PTR0), .A2(_01136__PTR1), .ZN(_02684__PTR1) );
  OR2_X1 U2345 ( .A1(_02683__PTR2), .A2(_02683__PTR34), .ZN(_01137__PTR0) );
  OR2_X1 U2346 ( .A1(_02683__PTR66), .A2(_02683__PTR98), .ZN(_01137__PTR1) );
  OR2_X1 U2347 ( .A1(_01137__PTR0), .A2(_01137__PTR1), .ZN(_02684__PTR2) );
  OR2_X1 U2348 ( .A1(_02683__PTR3), .A2(_02683__PTR35), .ZN(_01138__PTR0) );
  OR2_X1 U2349 ( .A1(_02683__PTR67), .A2(_02683__PTR99), .ZN(_01138__PTR1) );
  OR2_X1 U2350 ( .A1(_01138__PTR0), .A2(_01138__PTR1), .ZN(_02684__PTR3) );
  OR2_X1 U2351 ( .A1(_02683__PTR4), .A2(_02683__PTR36), .ZN(_01139__PTR0) );
  OR2_X1 U2352 ( .A1(_02683__PTR68), .A2(_02683__PTR100), .ZN(_01139__PTR1) );
  OR2_X1 U2353 ( .A1(_01139__PTR0), .A2(_01139__PTR1), .ZN(_02684__PTR4) );
  OR2_X1 U2354 ( .A1(_02683__PTR5), .A2(_02683__PTR37), .ZN(_01140__PTR0) );
  OR2_X1 U2355 ( .A1(_02683__PTR69), .A2(_02683__PTR101), .ZN(_01140__PTR1) );
  OR2_X1 U2356 ( .A1(_01140__PTR0), .A2(_01140__PTR1), .ZN(_02684__PTR5) );
  OR2_X1 U2357 ( .A1(_02683__PTR6), .A2(_02683__PTR38), .ZN(_01141__PTR0) );
  OR2_X1 U2358 ( .A1(_02683__PTR70), .A2(_02683__PTR102), .ZN(_01141__PTR1) );
  OR2_X1 U2359 ( .A1(_01141__PTR0), .A2(_01141__PTR1), .ZN(_02684__PTR6) );
  OR2_X1 U2360 ( .A1(_02683__PTR7), .A2(_02683__PTR39), .ZN(_01142__PTR0) );
  OR2_X1 U2361 ( .A1(_02683__PTR71), .A2(_02683__PTR103), .ZN(_01142__PTR1) );
  OR2_X1 U2362 ( .A1(_01142__PTR0), .A2(_01142__PTR1), .ZN(_02684__PTR7) );
  OR2_X1 U2363 ( .A1(_02683__PTR8), .A2(_02683__PTR40), .ZN(_01143__PTR0) );
  OR2_X1 U2364 ( .A1(_02683__PTR72), .A2(_02683__PTR104), .ZN(_01143__PTR1) );
  OR2_X1 U2365 ( .A1(_01143__PTR0), .A2(_01143__PTR1), .ZN(_02684__PTR8) );
  OR2_X1 U2366 ( .A1(_02683__PTR9), .A2(_02683__PTR41), .ZN(_01144__PTR0) );
  OR2_X1 U2367 ( .A1(_02683__PTR73), .A2(_02683__PTR105), .ZN(_01144__PTR1) );
  OR2_X1 U2368 ( .A1(_01144__PTR0), .A2(_01144__PTR1), .ZN(_02684__PTR9) );
  OR2_X1 U2369 ( .A1(_02683__PTR10), .A2(_02683__PTR42), .ZN(_01145__PTR0) );
  OR2_X1 U2370 ( .A1(_02683__PTR74), .A2(_02683__PTR106), .ZN(_01145__PTR1) );
  OR2_X1 U2371 ( .A1(_01145__PTR0), .A2(_01145__PTR1), .ZN(_02684__PTR10) );
  OR2_X1 U2372 ( .A1(_02683__PTR11), .A2(_02683__PTR43), .ZN(_01146__PTR0) );
  OR2_X1 U2373 ( .A1(_02683__PTR75), .A2(_02683__PTR107), .ZN(_01146__PTR1) );
  OR2_X1 U2374 ( .A1(_01146__PTR0), .A2(_01146__PTR1), .ZN(_02684__PTR11) );
  OR2_X1 U2375 ( .A1(_02683__PTR12), .A2(_02683__PTR44), .ZN(_01147__PTR0) );
  OR2_X1 U2376 ( .A1(_02683__PTR76), .A2(_02683__PTR108), .ZN(_01147__PTR1) );
  OR2_X1 U2377 ( .A1(_01147__PTR0), .A2(_01147__PTR1), .ZN(_02684__PTR12) );
  OR2_X1 U2378 ( .A1(_02683__PTR13), .A2(_02683__PTR45), .ZN(_01148__PTR0) );
  OR2_X1 U2379 ( .A1(_02683__PTR77), .A2(_02683__PTR109), .ZN(_01148__PTR1) );
  OR2_X1 U2380 ( .A1(_01148__PTR0), .A2(_01148__PTR1), .ZN(_02684__PTR13) );
  OR2_X1 U2381 ( .A1(_02683__PTR14), .A2(_02683__PTR46), .ZN(_01149__PTR0) );
  OR2_X1 U2382 ( .A1(_02683__PTR78), .A2(_02683__PTR110), .ZN(_01149__PTR1) );
  OR2_X1 U2383 ( .A1(_01149__PTR0), .A2(_01149__PTR1), .ZN(_02684__PTR14) );
  OR2_X1 U2384 ( .A1(_02683__PTR15), .A2(_02683__PTR47), .ZN(_01150__PTR0) );
  OR2_X1 U2385 ( .A1(_02683__PTR79), .A2(_02683__PTR111), .ZN(_01150__PTR1) );
  OR2_X1 U2386 ( .A1(_01150__PTR0), .A2(_01150__PTR1), .ZN(_02684__PTR15) );
  OR2_X1 U2387 ( .A1(_02683__PTR16), .A2(_02683__PTR48), .ZN(_01151__PTR0) );
  OR2_X1 U2388 ( .A1(_02683__PTR80), .A2(_02683__PTR112), .ZN(_01151__PTR1) );
  OR2_X1 U2389 ( .A1(_01151__PTR0), .A2(_01151__PTR1), .ZN(_02684__PTR16) );
  OR2_X1 U2390 ( .A1(_02683__PTR17), .A2(_02683__PTR49), .ZN(_01152__PTR0) );
  OR2_X1 U2391 ( .A1(_02683__PTR81), .A2(_02683__PTR113), .ZN(_01152__PTR1) );
  OR2_X1 U2392 ( .A1(_01152__PTR0), .A2(_01152__PTR1), .ZN(_02684__PTR17) );
  OR2_X1 U2393 ( .A1(_02683__PTR18), .A2(_02683__PTR50), .ZN(_01153__PTR0) );
  OR2_X1 U2394 ( .A1(_02683__PTR82), .A2(_02683__PTR114), .ZN(_01153__PTR1) );
  OR2_X1 U2395 ( .A1(_01153__PTR0), .A2(_01153__PTR1), .ZN(_02684__PTR18) );
  OR2_X1 U2396 ( .A1(_02683__PTR19), .A2(_02683__PTR51), .ZN(_01154__PTR0) );
  OR2_X1 U2397 ( .A1(_02683__PTR83), .A2(_02683__PTR115), .ZN(_01154__PTR1) );
  OR2_X1 U2398 ( .A1(_01154__PTR0), .A2(_01154__PTR1), .ZN(_02684__PTR19) );
  OR2_X1 U2399 ( .A1(_02683__PTR20), .A2(_02683__PTR52), .ZN(_01155__PTR0) );
  OR2_X1 U2400 ( .A1(_02683__PTR84), .A2(_02683__PTR116), .ZN(_01155__PTR1) );
  OR2_X1 U2401 ( .A1(_01155__PTR0), .A2(_01155__PTR1), .ZN(_02684__PTR20) );
  OR2_X1 U2402 ( .A1(_02683__PTR21), .A2(_02683__PTR53), .ZN(_01156__PTR0) );
  OR2_X1 U2403 ( .A1(_02683__PTR85), .A2(_02683__PTR117), .ZN(_01156__PTR1) );
  OR2_X1 U2404 ( .A1(_01156__PTR0), .A2(_01156__PTR1), .ZN(_02684__PTR21) );
  OR2_X1 U2405 ( .A1(_02683__PTR22), .A2(_02683__PTR54), .ZN(_01157__PTR0) );
  OR2_X1 U2406 ( .A1(_02683__PTR86), .A2(_02683__PTR118), .ZN(_01157__PTR1) );
  OR2_X1 U2407 ( .A1(_01157__PTR0), .A2(_01157__PTR1), .ZN(_02684__PTR22) );
  OR2_X1 U2408 ( .A1(_02683__PTR23), .A2(_02683__PTR55), .ZN(_01158__PTR0) );
  OR2_X1 U2409 ( .A1(_02683__PTR87), .A2(_02683__PTR119), .ZN(_01158__PTR1) );
  OR2_X1 U2410 ( .A1(_01158__PTR0), .A2(_01158__PTR1), .ZN(_02684__PTR23) );
  OR2_X1 U2411 ( .A1(_02683__PTR24), .A2(_02683__PTR56), .ZN(_01159__PTR0) );
  OR2_X1 U2412 ( .A1(_02683__PTR88), .A2(_02683__PTR120), .ZN(_01159__PTR1) );
  OR2_X1 U2413 ( .A1(_01159__PTR0), .A2(_01159__PTR1), .ZN(_02684__PTR24) );
  OR2_X1 U2414 ( .A1(_02683__PTR25), .A2(_02683__PTR57), .ZN(_01160__PTR0) );
  OR2_X1 U2415 ( .A1(_02683__PTR89), .A2(_02683__PTR121), .ZN(_01160__PTR1) );
  OR2_X1 U2416 ( .A1(_01160__PTR0), .A2(_01160__PTR1), .ZN(_02684__PTR25) );
  OR2_X1 U2417 ( .A1(_02683__PTR26), .A2(_02683__PTR58), .ZN(_01161__PTR0) );
  OR2_X1 U2418 ( .A1(_02683__PTR90), .A2(_02683__PTR122), .ZN(_01161__PTR1) );
  OR2_X1 U2419 ( .A1(_01161__PTR0), .A2(_01161__PTR1), .ZN(_02684__PTR26) );
  OR2_X1 U2420 ( .A1(_02683__PTR27), .A2(_02683__PTR59), .ZN(_01162__PTR0) );
  OR2_X1 U2421 ( .A1(_02683__PTR91), .A2(_02683__PTR123), .ZN(_01162__PTR1) );
  OR2_X1 U2422 ( .A1(_01162__PTR0), .A2(_01162__PTR1), .ZN(_02684__PTR27) );
  OR2_X1 U2423 ( .A1(_02683__PTR28), .A2(_02683__PTR60), .ZN(_01163__PTR0) );
  OR2_X1 U2424 ( .A1(_02683__PTR92), .A2(_02683__PTR124), .ZN(_01163__PTR1) );
  OR2_X1 U2425 ( .A1(_01163__PTR0), .A2(_01163__PTR1), .ZN(_02684__PTR28) );
  OR2_X1 U2426 ( .A1(_02683__PTR29), .A2(_02683__PTR61), .ZN(_01164__PTR0) );
  OR2_X1 U2427 ( .A1(_02683__PTR93), .A2(_02683__PTR125), .ZN(_01164__PTR1) );
  OR2_X1 U2428 ( .A1(_01164__PTR0), .A2(_01164__PTR1), .ZN(_02684__PTR29) );
  OR2_X1 U2429 ( .A1(_02683__PTR30), .A2(_02683__PTR62), .ZN(_01165__PTR0) );
  OR2_X1 U2430 ( .A1(_02683__PTR94), .A2(_02683__PTR126), .ZN(_01165__PTR1) );
  OR2_X1 U2431 ( .A1(_01165__PTR0), .A2(_01165__PTR1), .ZN(_02684__PTR30) );
  OR2_X1 U2432 ( .A1(_02683__PTR31), .A2(_02683__PTR63), .ZN(_01166__PTR0) );
  OR2_X1 U2433 ( .A1(_02683__PTR95), .A2(_02683__PTR127), .ZN(_01166__PTR1) );
  OR2_X1 U2434 ( .A1(_01166__PTR0), .A2(_01166__PTR1), .ZN(_02684__PTR31) );
  OR2_X1 U2435 ( .A1(_02445__PTR3), .A2(_02452__PTR0), .ZN(_01167__PTR0) );
  OR2_X1 U2436 ( .A1(_02445__PTR2), .A2(_02668__PTR4), .ZN(_02452__PTR1) );
  OR2_X1 U2437 ( .A1(_01167__PTR0), .A2(_02452__PTR1), .ZN(_03415_) );
  OR2_X1 U2438 ( .A1(_02663__PTR0), .A2(_02663__PTR32), .ZN(_01168__PTR0) );
  OR2_X1 U2439 ( .A1(_02663__PTR64), .A2(_02663__PTR96), .ZN(_01168__PTR1) );
  OR2_X1 U2440 ( .A1(_02663__PTR128), .A2(_02663__PTR160), .ZN(_01168__PTR2) );
  OR2_X1 U2441 ( .A1(_01168__PTR0), .A2(_01168__PTR1), .ZN(_01169__PTR0) );
  OR2_X1 U2442 ( .A1(_01168__PTR2), .A2(_02663__PTR192), .ZN(_01169__PTR1) );
  OR2_X1 U2443 ( .A1(_01169__PTR0), .A2(_01169__PTR1), .ZN(_02665__PTR0) );
  OR2_X1 U2444 ( .A1(_02663__PTR1), .A2(_02663__PTR33), .ZN(_01170__PTR0) );
  OR2_X1 U2445 ( .A1(_02663__PTR65), .A2(_02663__PTR97), .ZN(_01170__PTR1) );
  OR2_X1 U2446 ( .A1(_02663__PTR129), .A2(_02663__PTR161), .ZN(_01170__PTR2) );
  OR2_X1 U2447 ( .A1(_01170__PTR0), .A2(_01170__PTR1), .ZN(_01171__PTR0) );
  OR2_X1 U2448 ( .A1(_01170__PTR2), .A2(_02663__PTR193), .ZN(_01171__PTR1) );
  OR2_X1 U2449 ( .A1(_01171__PTR0), .A2(_01171__PTR1), .ZN(_02665__PTR1) );
  OR2_X1 U2450 ( .A1(_02663__PTR2), .A2(_02663__PTR34), .ZN(_01172__PTR0) );
  OR2_X1 U2451 ( .A1(_02663__PTR66), .A2(_02663__PTR98), .ZN(_01172__PTR1) );
  OR2_X1 U2452 ( .A1(_02663__PTR130), .A2(_02663__PTR162), .ZN(_01172__PTR2) );
  OR2_X1 U2453 ( .A1(_01172__PTR0), .A2(_01172__PTR1), .ZN(_01173__PTR0) );
  OR2_X1 U2454 ( .A1(_01172__PTR2), .A2(_02663__PTR194), .ZN(_01173__PTR1) );
  OR2_X1 U2455 ( .A1(_01173__PTR0), .A2(_01173__PTR1), .ZN(_02665__PTR2) );
  OR2_X1 U2456 ( .A1(_02663__PTR3), .A2(_02663__PTR35), .ZN(_01174__PTR0) );
  OR2_X1 U2457 ( .A1(_02663__PTR67), .A2(_02663__PTR99), .ZN(_01174__PTR1) );
  OR2_X1 U2458 ( .A1(_02663__PTR131), .A2(_02663__PTR163), .ZN(_01174__PTR2) );
  OR2_X1 U2459 ( .A1(_01174__PTR0), .A2(_01174__PTR1), .ZN(_01175__PTR0) );
  OR2_X1 U2460 ( .A1(_01174__PTR2), .A2(_02663__PTR195), .ZN(_01175__PTR1) );
  OR2_X1 U2461 ( .A1(_01175__PTR0), .A2(_01175__PTR1), .ZN(_02665__PTR3) );
  OR2_X1 U2462 ( .A1(_02663__PTR4), .A2(_02663__PTR36), .ZN(_01176__PTR0) );
  OR2_X1 U2463 ( .A1(_02663__PTR68), .A2(_02663__PTR100), .ZN(_01176__PTR1) );
  OR2_X1 U2464 ( .A1(_02663__PTR132), .A2(_02663__PTR164), .ZN(_01176__PTR2) );
  OR2_X1 U2465 ( .A1(_01176__PTR0), .A2(_01176__PTR1), .ZN(_01177__PTR0) );
  OR2_X1 U2466 ( .A1(_01176__PTR2), .A2(_02663__PTR196), .ZN(_01177__PTR1) );
  OR2_X1 U2467 ( .A1(_01177__PTR0), .A2(_01177__PTR1), .ZN(_02665__PTR4) );
  OR2_X1 U2468 ( .A1(_02663__PTR5), .A2(_02663__PTR37), .ZN(_01178__PTR0) );
  OR2_X1 U2469 ( .A1(_02663__PTR69), .A2(_02663__PTR101), .ZN(_01178__PTR1) );
  OR2_X1 U2470 ( .A1(_02663__PTR133), .A2(_02663__PTR165), .ZN(_01178__PTR2) );
  OR2_X1 U2471 ( .A1(_01178__PTR0), .A2(_01178__PTR1), .ZN(_01179__PTR0) );
  OR2_X1 U2472 ( .A1(_01178__PTR2), .A2(_02663__PTR197), .ZN(_01179__PTR1) );
  OR2_X1 U2473 ( .A1(_01179__PTR0), .A2(_01179__PTR1), .ZN(_02665__PTR5) );
  OR2_X1 U2474 ( .A1(_02663__PTR6), .A2(_02663__PTR38), .ZN(_01180__PTR0) );
  OR2_X1 U2475 ( .A1(_02663__PTR70), .A2(_02663__PTR102), .ZN(_01180__PTR1) );
  OR2_X1 U2476 ( .A1(_02663__PTR134), .A2(_02663__PTR166), .ZN(_01180__PTR2) );
  OR2_X1 U2477 ( .A1(_01180__PTR0), .A2(_01180__PTR1), .ZN(_01181__PTR0) );
  OR2_X1 U2478 ( .A1(_01180__PTR2), .A2(_02663__PTR198), .ZN(_01181__PTR1) );
  OR2_X1 U2479 ( .A1(_01181__PTR0), .A2(_01181__PTR1), .ZN(_02665__PTR6) );
  OR2_X1 U2480 ( .A1(_02663__PTR7), .A2(_02663__PTR39), .ZN(_01182__PTR0) );
  OR2_X1 U2481 ( .A1(_02663__PTR71), .A2(_02663__PTR103), .ZN(_01182__PTR1) );
  OR2_X1 U2482 ( .A1(_02663__PTR135), .A2(_02663__PTR167), .ZN(_01182__PTR2) );
  OR2_X1 U2483 ( .A1(_01182__PTR0), .A2(_01182__PTR1), .ZN(_01183__PTR0) );
  OR2_X1 U2484 ( .A1(_01182__PTR2), .A2(_02663__PTR199), .ZN(_01183__PTR1) );
  OR2_X1 U2485 ( .A1(_01183__PTR0), .A2(_01183__PTR1), .ZN(_02665__PTR7) );
  OR2_X1 U2486 ( .A1(_02663__PTR8), .A2(_02663__PTR40), .ZN(_01184__PTR0) );
  OR2_X1 U2487 ( .A1(_02663__PTR72), .A2(_02663__PTR104), .ZN(_01184__PTR1) );
  OR2_X1 U2488 ( .A1(_02663__PTR136), .A2(_02663__PTR168), .ZN(_01184__PTR2) );
  OR2_X1 U2489 ( .A1(_01184__PTR0), .A2(_01184__PTR1), .ZN(_01185__PTR0) );
  OR2_X1 U2490 ( .A1(_01184__PTR2), .A2(_02663__PTR200), .ZN(_01185__PTR1) );
  OR2_X1 U2491 ( .A1(_01185__PTR0), .A2(_01185__PTR1), .ZN(_02665__PTR8) );
  OR2_X1 U2492 ( .A1(_02663__PTR9), .A2(_02663__PTR41), .ZN(_01186__PTR0) );
  OR2_X1 U2493 ( .A1(_02663__PTR73), .A2(_02663__PTR105), .ZN(_01186__PTR1) );
  OR2_X1 U2494 ( .A1(_02663__PTR137), .A2(_02663__PTR169), .ZN(_01186__PTR2) );
  OR2_X1 U2495 ( .A1(_01186__PTR0), .A2(_01186__PTR1), .ZN(_01187__PTR0) );
  OR2_X1 U2496 ( .A1(_01186__PTR2), .A2(_02663__PTR201), .ZN(_01187__PTR1) );
  OR2_X1 U2497 ( .A1(_01187__PTR0), .A2(_01187__PTR1), .ZN(_02665__PTR9) );
  OR2_X1 U2498 ( .A1(_02663__PTR10), .A2(_02663__PTR42), .ZN(_01188__PTR0) );
  OR2_X1 U2499 ( .A1(_02663__PTR74), .A2(_02663__PTR106), .ZN(_01188__PTR1) );
  OR2_X1 U2500 ( .A1(_02663__PTR138), .A2(_02663__PTR170), .ZN(_01188__PTR2) );
  OR2_X1 U2501 ( .A1(_01188__PTR0), .A2(_01188__PTR1), .ZN(_01189__PTR0) );
  OR2_X1 U2502 ( .A1(_01188__PTR2), .A2(_02663__PTR202), .ZN(_01189__PTR1) );
  OR2_X1 U2503 ( .A1(_01189__PTR0), .A2(_01189__PTR1), .ZN(_02665__PTR10) );
  OR2_X1 U2504 ( .A1(_02663__PTR11), .A2(_02663__PTR43), .ZN(_01190__PTR0) );
  OR2_X1 U2505 ( .A1(_02663__PTR75), .A2(_02663__PTR107), .ZN(_01190__PTR1) );
  OR2_X1 U2506 ( .A1(_02663__PTR139), .A2(_02663__PTR171), .ZN(_01190__PTR2) );
  OR2_X1 U2507 ( .A1(_01190__PTR0), .A2(_01190__PTR1), .ZN(_01191__PTR0) );
  OR2_X1 U2508 ( .A1(_01190__PTR2), .A2(_02663__PTR203), .ZN(_01191__PTR1) );
  OR2_X1 U2509 ( .A1(_01191__PTR0), .A2(_01191__PTR1), .ZN(_02665__PTR11) );
  OR2_X1 U2510 ( .A1(_02663__PTR12), .A2(_02663__PTR44), .ZN(_01192__PTR0) );
  OR2_X1 U2511 ( .A1(_02663__PTR76), .A2(_02663__PTR108), .ZN(_01192__PTR1) );
  OR2_X1 U2512 ( .A1(_02663__PTR140), .A2(_02663__PTR172), .ZN(_01192__PTR2) );
  OR2_X1 U2513 ( .A1(_01192__PTR0), .A2(_01192__PTR1), .ZN(_01193__PTR0) );
  OR2_X1 U2514 ( .A1(_01192__PTR2), .A2(_02663__PTR204), .ZN(_01193__PTR1) );
  OR2_X1 U2515 ( .A1(_01193__PTR0), .A2(_01193__PTR1), .ZN(_02665__PTR12) );
  OR2_X1 U2516 ( .A1(_02663__PTR13), .A2(_02663__PTR45), .ZN(_01194__PTR0) );
  OR2_X1 U2517 ( .A1(_02663__PTR77), .A2(_02663__PTR109), .ZN(_01194__PTR1) );
  OR2_X1 U2518 ( .A1(_02663__PTR141), .A2(_02663__PTR173), .ZN(_01194__PTR2) );
  OR2_X1 U2519 ( .A1(_01194__PTR0), .A2(_01194__PTR1), .ZN(_01195__PTR0) );
  OR2_X1 U2520 ( .A1(_01194__PTR2), .A2(_02663__PTR205), .ZN(_01195__PTR1) );
  OR2_X1 U2521 ( .A1(_01195__PTR0), .A2(_01195__PTR1), .ZN(_02665__PTR13) );
  OR2_X1 U2522 ( .A1(_02663__PTR14), .A2(_02663__PTR46), .ZN(_01196__PTR0) );
  OR2_X1 U2523 ( .A1(_02663__PTR78), .A2(_02663__PTR110), .ZN(_01196__PTR1) );
  OR2_X1 U2524 ( .A1(_02663__PTR142), .A2(_02663__PTR174), .ZN(_01196__PTR2) );
  OR2_X1 U2525 ( .A1(_01196__PTR0), .A2(_01196__PTR1), .ZN(_01197__PTR0) );
  OR2_X1 U2526 ( .A1(_01196__PTR2), .A2(_02663__PTR206), .ZN(_01197__PTR1) );
  OR2_X1 U2527 ( .A1(_01197__PTR0), .A2(_01197__PTR1), .ZN(_02665__PTR14) );
  OR2_X1 U2528 ( .A1(_02663__PTR15), .A2(_02663__PTR47), .ZN(_01198__PTR0) );
  OR2_X1 U2529 ( .A1(_02663__PTR79), .A2(_02663__PTR111), .ZN(_01198__PTR1) );
  OR2_X1 U2530 ( .A1(_02663__PTR143), .A2(_02663__PTR175), .ZN(_01198__PTR2) );
  OR2_X1 U2531 ( .A1(_01198__PTR0), .A2(_01198__PTR1), .ZN(_01199__PTR0) );
  OR2_X1 U2532 ( .A1(_01198__PTR2), .A2(_02663__PTR207), .ZN(_01199__PTR1) );
  OR2_X1 U2533 ( .A1(_01199__PTR0), .A2(_01199__PTR1), .ZN(_02665__PTR15) );
  OR2_X1 U2534 ( .A1(_02663__PTR16), .A2(_02663__PTR48), .ZN(_01200__PTR0) );
  OR2_X1 U2535 ( .A1(_02663__PTR80), .A2(_02663__PTR112), .ZN(_01200__PTR1) );
  OR2_X1 U2536 ( .A1(_02663__PTR144), .A2(_02663__PTR176), .ZN(_01200__PTR2) );
  OR2_X1 U2537 ( .A1(_01200__PTR0), .A2(_01200__PTR1), .ZN(_01201__PTR0) );
  OR2_X1 U2538 ( .A1(_01200__PTR2), .A2(_02663__PTR208), .ZN(_01201__PTR1) );
  OR2_X1 U2539 ( .A1(_01201__PTR0), .A2(_01201__PTR1), .ZN(_02665__PTR16) );
  OR2_X1 U2540 ( .A1(_02663__PTR17), .A2(_02663__PTR49), .ZN(_01202__PTR0) );
  OR2_X1 U2541 ( .A1(_02663__PTR81), .A2(_02663__PTR113), .ZN(_01202__PTR1) );
  OR2_X1 U2542 ( .A1(_02663__PTR145), .A2(_02663__PTR177), .ZN(_01202__PTR2) );
  OR2_X1 U2543 ( .A1(_01202__PTR0), .A2(_01202__PTR1), .ZN(_01203__PTR0) );
  OR2_X1 U2544 ( .A1(_01202__PTR2), .A2(_02663__PTR209), .ZN(_01203__PTR1) );
  OR2_X1 U2545 ( .A1(_01203__PTR0), .A2(_01203__PTR1), .ZN(_02665__PTR17) );
  OR2_X1 U2546 ( .A1(_02663__PTR18), .A2(_02663__PTR50), .ZN(_01204__PTR0) );
  OR2_X1 U2547 ( .A1(_02663__PTR82), .A2(_02663__PTR114), .ZN(_01204__PTR1) );
  OR2_X1 U2548 ( .A1(_02663__PTR146), .A2(_02663__PTR178), .ZN(_01204__PTR2) );
  OR2_X1 U2549 ( .A1(_01204__PTR0), .A2(_01204__PTR1), .ZN(_01205__PTR0) );
  OR2_X1 U2550 ( .A1(_01204__PTR2), .A2(_02663__PTR210), .ZN(_01205__PTR1) );
  OR2_X1 U2551 ( .A1(_01205__PTR0), .A2(_01205__PTR1), .ZN(_02665__PTR18) );
  OR2_X1 U2552 ( .A1(_02663__PTR19), .A2(_02663__PTR51), .ZN(_01206__PTR0) );
  OR2_X1 U2553 ( .A1(_02663__PTR83), .A2(_02663__PTR115), .ZN(_01206__PTR1) );
  OR2_X1 U2554 ( .A1(_02663__PTR147), .A2(_02663__PTR179), .ZN(_01206__PTR2) );
  OR2_X1 U2555 ( .A1(_01206__PTR0), .A2(_01206__PTR1), .ZN(_01207__PTR0) );
  OR2_X1 U2556 ( .A1(_01206__PTR2), .A2(_02663__PTR211), .ZN(_01207__PTR1) );
  OR2_X1 U2557 ( .A1(_01207__PTR0), .A2(_01207__PTR1), .ZN(_02665__PTR19) );
  OR2_X1 U2558 ( .A1(_02663__PTR20), .A2(_02663__PTR52), .ZN(_01208__PTR0) );
  OR2_X1 U2559 ( .A1(_02663__PTR84), .A2(_02663__PTR116), .ZN(_01208__PTR1) );
  OR2_X1 U2560 ( .A1(_02663__PTR148), .A2(_02663__PTR180), .ZN(_01208__PTR2) );
  OR2_X1 U2561 ( .A1(_01208__PTR0), .A2(_01208__PTR1), .ZN(_01209__PTR0) );
  OR2_X1 U2562 ( .A1(_01208__PTR2), .A2(_02663__PTR212), .ZN(_01209__PTR1) );
  OR2_X1 U2563 ( .A1(_01209__PTR0), .A2(_01209__PTR1), .ZN(_02665__PTR20) );
  OR2_X1 U2564 ( .A1(_02663__PTR21), .A2(_02663__PTR53), .ZN(_01210__PTR0) );
  OR2_X1 U2565 ( .A1(_02663__PTR85), .A2(_02663__PTR117), .ZN(_01210__PTR1) );
  OR2_X1 U2566 ( .A1(_02663__PTR149), .A2(_02663__PTR181), .ZN(_01210__PTR2) );
  OR2_X1 U2567 ( .A1(_01210__PTR0), .A2(_01210__PTR1), .ZN(_01211__PTR0) );
  OR2_X1 U2568 ( .A1(_01210__PTR2), .A2(_02663__PTR213), .ZN(_01211__PTR1) );
  OR2_X1 U2569 ( .A1(_01211__PTR0), .A2(_01211__PTR1), .ZN(_02665__PTR21) );
  OR2_X1 U2570 ( .A1(_02663__PTR22), .A2(_02663__PTR54), .ZN(_01212__PTR0) );
  OR2_X1 U2571 ( .A1(_02663__PTR86), .A2(_02663__PTR118), .ZN(_01212__PTR1) );
  OR2_X1 U2572 ( .A1(_02663__PTR150), .A2(_02663__PTR182), .ZN(_01212__PTR2) );
  OR2_X1 U2573 ( .A1(_01212__PTR0), .A2(_01212__PTR1), .ZN(_01213__PTR0) );
  OR2_X1 U2574 ( .A1(_01212__PTR2), .A2(_02663__PTR214), .ZN(_01213__PTR1) );
  OR2_X1 U2575 ( .A1(_01213__PTR0), .A2(_01213__PTR1), .ZN(_02665__PTR22) );
  OR2_X1 U2576 ( .A1(_02663__PTR23), .A2(_02663__PTR55), .ZN(_01214__PTR0) );
  OR2_X1 U2577 ( .A1(_02663__PTR87), .A2(_02663__PTR119), .ZN(_01214__PTR1) );
  OR2_X1 U2578 ( .A1(_02663__PTR151), .A2(_02663__PTR183), .ZN(_01214__PTR2) );
  OR2_X1 U2579 ( .A1(_01214__PTR0), .A2(_01214__PTR1), .ZN(_01215__PTR0) );
  OR2_X1 U2580 ( .A1(_01214__PTR2), .A2(_02663__PTR215), .ZN(_01215__PTR1) );
  OR2_X1 U2581 ( .A1(_01215__PTR0), .A2(_01215__PTR1), .ZN(_02665__PTR23) );
  OR2_X1 U2582 ( .A1(_02663__PTR24), .A2(_02663__PTR56), .ZN(_01216__PTR0) );
  OR2_X1 U2583 ( .A1(_02663__PTR88), .A2(_02663__PTR120), .ZN(_01216__PTR1) );
  OR2_X1 U2584 ( .A1(_02663__PTR152), .A2(_02663__PTR184), .ZN(_01216__PTR2) );
  OR2_X1 U2585 ( .A1(_01216__PTR0), .A2(_01216__PTR1), .ZN(_01217__PTR0) );
  OR2_X1 U2586 ( .A1(_01216__PTR2), .A2(_02663__PTR216), .ZN(_01217__PTR1) );
  OR2_X1 U2587 ( .A1(_01217__PTR0), .A2(_01217__PTR1), .ZN(_02665__PTR24) );
  OR2_X1 U2588 ( .A1(_02663__PTR25), .A2(_02663__PTR57), .ZN(_01218__PTR0) );
  OR2_X1 U2589 ( .A1(_02663__PTR89), .A2(_02663__PTR121), .ZN(_01218__PTR1) );
  OR2_X1 U2590 ( .A1(_02663__PTR153), .A2(_02663__PTR185), .ZN(_01218__PTR2) );
  OR2_X1 U2591 ( .A1(_01218__PTR0), .A2(_01218__PTR1), .ZN(_01219__PTR0) );
  OR2_X1 U2592 ( .A1(_01218__PTR2), .A2(_02663__PTR217), .ZN(_01219__PTR1) );
  OR2_X1 U2593 ( .A1(_01219__PTR0), .A2(_01219__PTR1), .ZN(_02665__PTR25) );
  OR2_X1 U2594 ( .A1(_02663__PTR26), .A2(_02663__PTR58), .ZN(_01220__PTR0) );
  OR2_X1 U2595 ( .A1(_02663__PTR90), .A2(_02663__PTR122), .ZN(_01220__PTR1) );
  OR2_X1 U2596 ( .A1(_02663__PTR154), .A2(_02663__PTR186), .ZN(_01220__PTR2) );
  OR2_X1 U2597 ( .A1(_01220__PTR0), .A2(_01220__PTR1), .ZN(_01221__PTR0) );
  OR2_X1 U2598 ( .A1(_01220__PTR2), .A2(_02663__PTR218), .ZN(_01221__PTR1) );
  OR2_X1 U2599 ( .A1(_01221__PTR0), .A2(_01221__PTR1), .ZN(_02665__PTR26) );
  OR2_X1 U2600 ( .A1(_02663__PTR27), .A2(_02663__PTR59), .ZN(_01222__PTR0) );
  OR2_X1 U2601 ( .A1(_02663__PTR91), .A2(_02663__PTR123), .ZN(_01222__PTR1) );
  OR2_X1 U2602 ( .A1(_02663__PTR155), .A2(_02663__PTR187), .ZN(_01222__PTR2) );
  OR2_X1 U2603 ( .A1(_01222__PTR0), .A2(_01222__PTR1), .ZN(_01223__PTR0) );
  OR2_X1 U2604 ( .A1(_01222__PTR2), .A2(_02663__PTR219), .ZN(_01223__PTR1) );
  OR2_X1 U2605 ( .A1(_01223__PTR0), .A2(_01223__PTR1), .ZN(_02665__PTR27) );
  OR2_X1 U2606 ( .A1(_02663__PTR28), .A2(_02663__PTR60), .ZN(_01224__PTR0) );
  OR2_X1 U2607 ( .A1(_02663__PTR92), .A2(_02663__PTR124), .ZN(_01224__PTR1) );
  OR2_X1 U2608 ( .A1(_02663__PTR156), .A2(_02663__PTR188), .ZN(_01224__PTR2) );
  OR2_X1 U2609 ( .A1(_01224__PTR0), .A2(_01224__PTR1), .ZN(_01225__PTR0) );
  OR2_X1 U2610 ( .A1(_01224__PTR2), .A2(_02663__PTR220), .ZN(_01225__PTR1) );
  OR2_X1 U2611 ( .A1(_01225__PTR0), .A2(_01225__PTR1), .ZN(_02665__PTR28) );
  OR2_X1 U2612 ( .A1(_02663__PTR29), .A2(_02663__PTR61), .ZN(_01226__PTR0) );
  OR2_X1 U2613 ( .A1(_02663__PTR93), .A2(_02663__PTR125), .ZN(_01226__PTR1) );
  OR2_X1 U2614 ( .A1(_02663__PTR157), .A2(_02663__PTR189), .ZN(_01226__PTR2) );
  OR2_X1 U2615 ( .A1(_01226__PTR0), .A2(_01226__PTR1), .ZN(_01227__PTR0) );
  OR2_X1 U2616 ( .A1(_01226__PTR2), .A2(_02663__PTR221), .ZN(_01227__PTR1) );
  OR2_X1 U2617 ( .A1(_01227__PTR0), .A2(_01227__PTR1), .ZN(_02665__PTR29) );
  OR2_X1 U2618 ( .A1(_02663__PTR30), .A2(_02663__PTR62), .ZN(_01228__PTR0) );
  OR2_X1 U2619 ( .A1(_02663__PTR94), .A2(_02663__PTR126), .ZN(_01228__PTR1) );
  OR2_X1 U2620 ( .A1(_02663__PTR158), .A2(_02663__PTR190), .ZN(_01228__PTR2) );
  OR2_X1 U2621 ( .A1(_01228__PTR0), .A2(_01228__PTR1), .ZN(_01229__PTR0) );
  OR2_X1 U2622 ( .A1(_01228__PTR2), .A2(_02663__PTR222), .ZN(_01229__PTR1) );
  OR2_X1 U2623 ( .A1(_01229__PTR0), .A2(_01229__PTR1), .ZN(_02665__PTR30) );
  OR2_X1 U2624 ( .A1(_02663__PTR31), .A2(_02663__PTR63), .ZN(_01230__PTR0) );
  OR2_X1 U2625 ( .A1(_02663__PTR95), .A2(_02663__PTR127), .ZN(_01230__PTR1) );
  OR2_X1 U2626 ( .A1(_02663__PTR159), .A2(_02663__PTR191), .ZN(_01230__PTR2) );
  OR2_X1 U2627 ( .A1(_01230__PTR0), .A2(_01230__PTR1), .ZN(_01231__PTR0) );
  OR2_X1 U2628 ( .A1(_01230__PTR2), .A2(_02663__PTR223), .ZN(_01231__PTR1) );
  OR2_X1 U2629 ( .A1(_01231__PTR0), .A2(_01231__PTR1), .ZN(_02665__PTR31) );
  OR2_X1 U2630 ( .A1(_02664__PTR0), .A2(_02664__PTR1), .ZN(_01129__PTR0) );
  OR2_X1 U2631 ( .A1(_02437__PTR0), .A2(_02437__PTR1), .ZN(_01117__PTR0) );
  OR2_X1 U2632 ( .A1(_02664__PTR4), .A2(_02437__PTR2), .ZN(_02441__PTR2) );
  OR2_X1 U2633 ( .A1(_01129__PTR0), .A2(_01117__PTR0), .ZN(_01232__PTR0) );
  OR2_X1 U2634 ( .A1(_02441__PTR2), .A2(_02437__PTR3), .ZN(_01117__PTR1) );
  OR2_X1 U2635 ( .A1(_01232__PTR0), .A2(_01117__PTR1), .ZN(_03410_) );
  OR2_X1 U2636 ( .A1(_02671__PTR0), .A2(_02671__PTR32), .ZN(_01233_) );
  OR2_X1 U2637 ( .A1(_01233_), .A2(_02671__PTR64), .ZN(_02673__PTR0) );
  OR2_X1 U2638 ( .A1(_02671__PTR1), .A2(_02671__PTR33), .ZN(_01234_) );
  OR2_X1 U2639 ( .A1(_01234_), .A2(_02671__PTR65), .ZN(_02673__PTR1) );
  OR2_X1 U2640 ( .A1(_02671__PTR2), .A2(_02671__PTR34), .ZN(_01235_) );
  OR2_X1 U2641 ( .A1(_01235_), .A2(_02671__PTR66), .ZN(_02673__PTR2) );
  OR2_X1 U2642 ( .A1(_02671__PTR3), .A2(_02671__PTR35), .ZN(_01236_) );
  OR2_X1 U2643 ( .A1(_01236_), .A2(_02671__PTR67), .ZN(_02673__PTR3) );
  OR2_X1 U2644 ( .A1(_02671__PTR4), .A2(_02671__PTR36), .ZN(_01237_) );
  OR2_X1 U2645 ( .A1(_01237_), .A2(_02671__PTR68), .ZN(_02673__PTR4) );
  OR2_X1 U2646 ( .A1(_02671__PTR5), .A2(_02671__PTR37), .ZN(_01238_) );
  OR2_X1 U2647 ( .A1(_01238_), .A2(_02671__PTR69), .ZN(_02673__PTR5) );
  OR2_X1 U2648 ( .A1(_02671__PTR6), .A2(_02671__PTR38), .ZN(_01239_) );
  OR2_X1 U2649 ( .A1(_01239_), .A2(_02671__PTR70), .ZN(_02673__PTR6) );
  OR2_X1 U2650 ( .A1(_02671__PTR7), .A2(_02671__PTR39), .ZN(_01240_) );
  OR2_X1 U2651 ( .A1(_01240_), .A2(_02671__PTR71), .ZN(_02673__PTR7) );
  OR2_X1 U2652 ( .A1(_02671__PTR8), .A2(_02671__PTR40), .ZN(_01241_) );
  OR2_X1 U2653 ( .A1(_01241_), .A2(_02671__PTR72), .ZN(_02673__PTR8) );
  OR2_X1 U2654 ( .A1(_02671__PTR9), .A2(_02671__PTR41), .ZN(_01242_) );
  OR2_X1 U2655 ( .A1(_01242_), .A2(_02671__PTR73), .ZN(_02673__PTR9) );
  OR2_X1 U2656 ( .A1(_02671__PTR10), .A2(_02671__PTR42), .ZN(_01243_) );
  OR2_X1 U2657 ( .A1(_01243_), .A2(_02671__PTR74), .ZN(_02673__PTR10) );
  OR2_X1 U2658 ( .A1(_02671__PTR11), .A2(_02671__PTR43), .ZN(_01244_) );
  OR2_X1 U2659 ( .A1(_01244_), .A2(_02671__PTR75), .ZN(_02673__PTR11) );
  OR2_X1 U2660 ( .A1(_02671__PTR12), .A2(_02671__PTR44), .ZN(_01245_) );
  OR2_X1 U2661 ( .A1(_01245_), .A2(_02671__PTR76), .ZN(_02673__PTR12) );
  OR2_X1 U2662 ( .A1(_02671__PTR13), .A2(_02671__PTR45), .ZN(_01246_) );
  OR2_X1 U2663 ( .A1(_01246_), .A2(_02671__PTR77), .ZN(_02673__PTR13) );
  OR2_X1 U2664 ( .A1(_02671__PTR14), .A2(_02671__PTR46), .ZN(_01247_) );
  OR2_X1 U2665 ( .A1(_01247_), .A2(_02671__PTR78), .ZN(_02673__PTR14) );
  OR2_X1 U2666 ( .A1(_02671__PTR15), .A2(_02671__PTR47), .ZN(_01248_) );
  OR2_X1 U2667 ( .A1(_01248_), .A2(_02671__PTR79), .ZN(_02673__PTR15) );
  OR2_X1 U2668 ( .A1(_02671__PTR16), .A2(_02671__PTR48), .ZN(_01249_) );
  OR2_X1 U2669 ( .A1(_01249_), .A2(_02671__PTR80), .ZN(_02673__PTR16) );
  OR2_X1 U2670 ( .A1(_02671__PTR17), .A2(_02671__PTR49), .ZN(_01250_) );
  OR2_X1 U2671 ( .A1(_01250_), .A2(_02671__PTR81), .ZN(_02673__PTR17) );
  OR2_X1 U2672 ( .A1(_02671__PTR18), .A2(_02671__PTR50), .ZN(_01251_) );
  OR2_X1 U2673 ( .A1(_01251_), .A2(_02671__PTR82), .ZN(_02673__PTR18) );
  OR2_X1 U2674 ( .A1(_02671__PTR19), .A2(_02671__PTR51), .ZN(_01252_) );
  OR2_X1 U2675 ( .A1(_01252_), .A2(_02671__PTR83), .ZN(_02673__PTR19) );
  OR2_X1 U2676 ( .A1(_02671__PTR20), .A2(_02671__PTR52), .ZN(_01253_) );
  OR2_X1 U2677 ( .A1(_01253_), .A2(_02671__PTR84), .ZN(_02673__PTR20) );
  OR2_X1 U2678 ( .A1(_02671__PTR21), .A2(_02671__PTR53), .ZN(_01254_) );
  OR2_X1 U2679 ( .A1(_01254_), .A2(_02671__PTR85), .ZN(_02673__PTR21) );
  OR2_X1 U2680 ( .A1(_02671__PTR22), .A2(_02671__PTR54), .ZN(_01255_) );
  OR2_X1 U2681 ( .A1(_01255_), .A2(_02671__PTR86), .ZN(_02673__PTR22) );
  OR2_X1 U2682 ( .A1(_02671__PTR23), .A2(_02671__PTR55), .ZN(_01256_) );
  OR2_X1 U2683 ( .A1(_01256_), .A2(_02671__PTR87), .ZN(_02673__PTR23) );
  OR2_X1 U2684 ( .A1(_02671__PTR24), .A2(_02671__PTR56), .ZN(_01257_) );
  OR2_X1 U2685 ( .A1(_01257_), .A2(_02671__PTR88), .ZN(_02673__PTR24) );
  OR2_X1 U2686 ( .A1(_02671__PTR25), .A2(_02671__PTR57), .ZN(_01258_) );
  OR2_X1 U2687 ( .A1(_01258_), .A2(_02671__PTR89), .ZN(_02673__PTR25) );
  OR2_X1 U2688 ( .A1(_02671__PTR26), .A2(_02671__PTR58), .ZN(_01259_) );
  OR2_X1 U2689 ( .A1(_01259_), .A2(_02671__PTR90), .ZN(_02673__PTR26) );
  OR2_X1 U2690 ( .A1(_02671__PTR27), .A2(_02671__PTR59), .ZN(_01260_) );
  OR2_X1 U2691 ( .A1(_01260_), .A2(_02671__PTR91), .ZN(_02673__PTR27) );
  OR2_X1 U2692 ( .A1(_02671__PTR28), .A2(_02671__PTR60), .ZN(_01261_) );
  OR2_X1 U2693 ( .A1(_01261_), .A2(_02671__PTR92), .ZN(_02673__PTR28) );
  OR2_X1 U2694 ( .A1(_02671__PTR29), .A2(_02671__PTR61), .ZN(_01262_) );
  OR2_X1 U2695 ( .A1(_01262_), .A2(_02671__PTR93), .ZN(_02673__PTR29) );
  OR2_X1 U2696 ( .A1(_02671__PTR30), .A2(_02671__PTR62), .ZN(_01263_) );
  OR2_X1 U2697 ( .A1(_01263_), .A2(_02671__PTR94), .ZN(_02673__PTR30) );
  OR2_X1 U2698 ( .A1(_02671__PTR31), .A2(_02671__PTR63), .ZN(_01264_) );
  OR2_X1 U2699 ( .A1(_01264_), .A2(_02671__PTR95), .ZN(_02673__PTR31) );
  OR2_X1 U2700 ( .A1(_02672__PTR0), .A2(_02437__PTR2), .ZN(_01265_) );
  OR2_X1 U2701 ( .A1(_01265_), .A2(_02437__PTR3), .ZN(_03412_) );
  OR2_X1 U2702 ( .A1(_03242_), .A2(_03243_), .ZN(_01766__PTR2) );
  AND2_X1 U2703 ( .A1(_03240__PTR1), .A2(_03302__PTR1), .ZN(_03240__PTR3) );
  OR2_X1 U2704 ( .A1(_02697__PTR0), .A2(_02697__PTR4), .ZN(_02700__PTR0) );
  OR2_X1 U2705 ( .A1(_02697__PTR1), .A2(_02697__PTR5), .ZN(_02700__PTR1) );
  OR2_X1 U2706 ( .A1(_02697__PTR2), .A2(_02697__PTR6), .ZN(_02700__PTR2) );
  OR2_X1 U2707 ( .A1(_02697__PTR3), .A2(_02697__PTR7), .ZN(_02700__PTR3) );
  OR2_X1 U2708 ( .A1(_02698__PTR0), .A2(_02445__PTR2), .ZN(_03418_) );
  OR2_X1 U2709 ( .A1(_03220_), .A2(_03221_), .ZN(_02585_) );
  AND2_X1 U2710 ( .A1(_01266__PTR0), .A2(_03209__PTR3), .ZN(_01267_) );
  AND2_X1 U2711 ( .A1(_01267_), .A2(_01266__PTR2), .ZN(_03221_) );
  OR2_X1 U2712 ( .A1(_03217_), .A2(_03218_), .ZN(_02435__PTR2) );
  AND2_X1 U2713 ( .A1(_03207__PTR0), .A2(_03208__PTR1), .ZN(_01268__PTR0) );
  AND2_X1 U2714 ( .A1(_01268__PTR0), .A2(_01268__PTR1), .ZN(_01269_) );
  AND2_X1 U2715 ( .A1(_01269_), .A2(_01266__PTR2), .ZN(_03218_) );
  OR2_X1 U2716 ( .A1(_03211_), .A2(_03212_), .ZN(_02435__PTR3) );
  AND2_X1 U2717 ( .A1(_03207__PTR0), .A2(_03207__PTR1), .ZN(_01270__PTR0) );
  AND2_X1 U2718 ( .A1(_01270__PTR0), .A2(_03209__PTR3), .ZN(_01271_) );
  AND2_X1 U2719 ( .A1(_01271_), .A2(_01266__PTR2), .ZN(_03212_) );
  OR2_X1 U2720 ( .A1(_00306_), .A2(_00288_), .ZN(_01272__PTR0) );
  OR2_X1 U2721 ( .A1(P3_State_PTR2), .A2(_00307_), .ZN(_01272__PTR1) );
  OR2_X1 U2722 ( .A1(_01272__PTR0), .A2(_01272__PTR1), .ZN(_01273_) );
  OR2_X1 U2723 ( .A1(_01273_), .A2(_01765__PTR4), .ZN(_00000_) );
  OR2_X1 U2724 ( .A1(_01275_), .A2(_00287_), .ZN(_00003_) );
  OR2_X1 U2725 ( .A1(_00288_), .A2(_00287_), .ZN(_00004_) );
  AND2_X1 U2726 ( .A1(_00001_), .A2(_00002_), .ZN(_01276__PTR0) );
  AND2_X1 U2727 ( .A1(_00003_), .A2(_00004_), .ZN(_01276__PTR1) );
  AND2_X1 U2728 ( .A1(_01276__PTR0), .A2(_01276__PTR1), .ZN(_00154_) );
  OR2_X1 U2729 ( .A1(_00299_), .A2(_02475__PTR14), .ZN(_01277__PTR1) );
  OR2_X1 U2730 ( .A1(_01277__PTR0), .A2(_01277__PTR1), .ZN(_00005_) );
  OR2_X1 U2731 ( .A1(_00151_), .A2(_00299_), .ZN(_00006_) );
  AND2_X1 U2732 ( .A1(_00005_), .A2(_00006_), .ZN(_01278_) );
  AND2_X1 U2733 ( .A1(_01278_), .A2(_00292_), .ZN(_00155_) );
  OR2_X1 U2734 ( .A1(_00151_), .A2(P3_P1_State2_PTR2), .ZN(_00011_) );
  AND2_X1 U2735 ( .A1(_00011_), .A2(_00009_), .ZN(_01282_) );
  AND2_X1 U2736 ( .A1(_01282_), .A2(_00292_), .ZN(_00158_) );
  AND2_X1 U2737 ( .A1(_01280__PTR0), .A2(P3_P1_State2_PTR2), .ZN(_00159_) );
  OR2_X1 U2738 ( .A1(_01310__PTR0), .A2(_01283__PTR1), .ZN(_00026_) );
  AND2_X1 U2739 ( .A1(_00026_), .A2(_00013_), .ZN(_01311__PTR0) );
  AND2_X1 U2740 ( .A1(_01311__PTR0), .A2(_01287__PTR1), .ZN(_01312__PTR0) );
  AND2_X1 U2741 ( .A1(_01312__PTR0), .A2(_01288__PTR1), .ZN(_00168_) );
  OR2_X1 U2742 ( .A1(_01313__PTR0), .A2(_01283__PTR1), .ZN(_00027_) );
  AND2_X1 U2743 ( .A1(_00027_), .A2(_00013_), .ZN(_01314__PTR0) );
  AND2_X1 U2744 ( .A1(_01314__PTR0), .A2(_01287__PTR1), .ZN(_01315__PTR0) );
  AND2_X1 U2745 ( .A1(_01315__PTR0), .A2(_01288__PTR1), .ZN(_00169_) );
  OR2_X1 U2746 ( .A1(_01316__PTR0), .A2(_01283__PTR1), .ZN(_00028_) );
  AND2_X1 U2747 ( .A1(_00028_), .A2(_00013_), .ZN(_01317__PTR0) );
  AND2_X1 U2748 ( .A1(_01317__PTR0), .A2(_01287__PTR1), .ZN(_01318__PTR0) );
  AND2_X1 U2749 ( .A1(_01318__PTR0), .A2(_01288__PTR1), .ZN(_00170_) );
  OR2_X1 U2750 ( .A1(_01319__PTR0), .A2(_01283__PTR1), .ZN(_00029_) );
  AND2_X1 U2751 ( .A1(_00029_), .A2(_00013_), .ZN(_01320__PTR0) );
  AND2_X1 U2752 ( .A1(_01320__PTR0), .A2(_01287__PTR1), .ZN(_01321__PTR0) );
  AND2_X1 U2753 ( .A1(_01321__PTR0), .A2(_01288__PTR1), .ZN(_00171_) );
  OR2_X1 U2754 ( .A1(_01322__PTR0), .A2(_01283__PTR1), .ZN(_00030_) );
  AND2_X1 U2755 ( .A1(_00030_), .A2(_00013_), .ZN(_01323__PTR0) );
  AND2_X1 U2756 ( .A1(_01323__PTR0), .A2(_01287__PTR1), .ZN(_01324__PTR0) );
  AND2_X1 U2757 ( .A1(_01324__PTR0), .A2(_01288__PTR1), .ZN(_00172_) );
  OR2_X1 U2758 ( .A1(_01325__PTR0), .A2(_01283__PTR1), .ZN(_00031_) );
  AND2_X1 U2759 ( .A1(_00031_), .A2(_00013_), .ZN(_01326__PTR0) );
  AND2_X1 U2760 ( .A1(_01326__PTR0), .A2(_01287__PTR1), .ZN(_01327__PTR0) );
  AND2_X1 U2761 ( .A1(_01327__PTR0), .A2(_01288__PTR1), .ZN(_00173_) );
  OR2_X1 U2762 ( .A1(_01328__PTR0), .A2(_01283__PTR1), .ZN(_00032_) );
  AND2_X1 U2763 ( .A1(_00032_), .A2(_00013_), .ZN(_01329__PTR0) );
  AND2_X1 U2764 ( .A1(_01329__PTR0), .A2(_01287__PTR1), .ZN(_01330__PTR0) );
  AND2_X1 U2765 ( .A1(_01330__PTR0), .A2(_01288__PTR1), .ZN(_00174_) );
  OR2_X1 U2766 ( .A1(_01331__PTR0), .A2(_01283__PTR1), .ZN(_00033_) );
  AND2_X1 U2767 ( .A1(_00033_), .A2(_00013_), .ZN(_01332__PTR0) );
  AND2_X1 U2768 ( .A1(_01332__PTR0), .A2(_01287__PTR1), .ZN(_01333__PTR0) );
  AND2_X1 U2769 ( .A1(_01333__PTR0), .A2(_01288__PTR1), .ZN(_00175_) );
  OR2_X1 U2770 ( .A1(P3_P1_Flush), .A2(_00308_), .ZN(_01334__PTR2) );
  OR2_X1 U2771 ( .A1(_00151_), .A2(_01281__PTR1), .ZN(_01335_) );
  OR2_X1 U2772 ( .A1(_01335_), .A2(_01334__PTR2), .ZN(_00035_) );
  AND2_X1 U2773 ( .A1(_00034_), .A2(_00013_), .ZN(_01336__PTR0) );
  AND2_X1 U2774 ( .A1(_00035_), .A2(_00016_), .ZN(_01336__PTR1) );
  AND2_X1 U2775 ( .A1(_01336__PTR0), .A2(_01336__PTR1), .ZN(_01337_) );
  AND2_X1 U2776 ( .A1(_01337_), .A2(_00017_), .ZN(_00176_) );
  AND2_X1 U2777 ( .A1(_00036_), .A2(_00034_), .ZN(_01338__PTR0) );
  AND2_X1 U2778 ( .A1(_00016_), .A2(_00037_), .ZN(_01338__PTR1) );
  AND2_X1 U2779 ( .A1(_01338__PTR0), .A2(_01338__PTR1), .ZN(_00177_) );
  OR2_X1 U2780 ( .A1(_01285__PTR0), .A2(P3_P1_State2_PTR2), .ZN(_00038_) );
  AND2_X1 U2781 ( .A1(_00007_), .A2(_00038_), .ZN(_01339__PTR0) );
  AND2_X1 U2782 ( .A1(_01339__PTR0), .A2(_01339__PTR1), .ZN(_01340_) );
  AND2_X1 U2783 ( .A1(_01340_), .A2(_00292_), .ZN(_00178_) );
  AND2_X1 U2784 ( .A1(_00007_), .A2(_00008_), .ZN(_01279__PTR0) );
  AND2_X1 U2785 ( .A1(_00009_), .A2(_00292_), .ZN(_01279__PTR1) );
  AND2_X1 U2786 ( .A1(_01279__PTR0), .A2(_01279__PTR1), .ZN(_00156_) );
  AND2_X1 U2787 ( .A1(P3_P1_State2_PTR0), .A2(_00293_), .ZN(_01280__PTR0) );
  AND2_X1 U2788 ( .A1(P3_P1_State2_PTR2), .A2(_00292_), .ZN(_01280__PTR1) );
  AND2_X1 U2789 ( .A1(_01280__PTR0), .A2(_01280__PTR1), .ZN(_00157_) );
  OR2_X1 U2790 ( .A1(_00306_), .A2(P3_State_PTR1), .ZN(_01275_) );
  OR2_X1 U2791 ( .A1(_01275_), .A2(P3_State_PTR2), .ZN(_00002_) );
  OR2_X1 U2792 ( .A1(P3_State_PTR1), .A2(_00287_), .ZN(_00039_) );
  AND2_X1 U2793 ( .A1(_00002_), .A2(_00039_), .ZN(_00179_) );
  OR2_X1 U2794 ( .A1(_00150_), .A2(P3_P1_State2_PTR2), .ZN(_00040_) );
  OR2_X1 U2795 ( .A1(_00150_), .A2(_00299_), .ZN(_00007_) );
  OR2_X1 U2796 ( .A1(_00293_), .A2(P3_P1_State2_PTR2), .ZN(_00008_) );
  AND2_X1 U2797 ( .A1(_00040_), .A2(_00007_), .ZN(_01341__PTR0) );
  AND2_X1 U2798 ( .A1(_00008_), .A2(_00009_), .ZN(_01339__PTR1) );
  AND2_X1 U2799 ( .A1(_01341__PTR0), .A2(_01339__PTR1), .ZN(_01342_) );
  AND2_X1 U2800 ( .A1(_01342_), .A2(_00292_), .ZN(_00180_) );
  OR2_X1 U2801 ( .A1(_00301_), .A2(_02186__PTR14), .ZN(_01349__PTR1) );
  OR2_X1 U2802 ( .A1(_01349__PTR0), .A2(_01349__PTR1), .ZN(_00049_) );
  OR2_X1 U2803 ( .A1(_00145_), .A2(_00301_), .ZN(_00050_) );
  AND2_X1 U2804 ( .A1(_00049_), .A2(_00050_), .ZN(_01350_) );
  AND2_X1 U2805 ( .A1(_01350_), .A2(_00294_), .ZN(_00183_) );
  AND2_X1 U2806 ( .A1(_01352__PTR0), .A2(_01352__PTR1), .ZN(_00185_) );
  AND2_X1 U2807 ( .A1(P2_P1_State2_PTR0), .A2(_00295_), .ZN(_01352__PTR0) );
  AND2_X1 U2808 ( .A1(P2_P1_State2_PTR2), .A2(_00294_), .ZN(_01352__PTR1) );
  OR2_X1 U2809 ( .A1(P2_P1_State2_PTR0), .A2(_00295_), .ZN(_01349__PTR0) );
  OR2_X1 U2810 ( .A1(_01349__PTR0), .A2(_01353__PTR1), .ZN(_00078_) );
  OR2_X1 U2811 ( .A1(_00078_), .A2(_02186__PTR14), .ZN(_00054_) );
  OR2_X1 U2812 ( .A1(_00145_), .A2(P2_P1_State2_PTR2), .ZN(_00055_) );
  OR2_X1 U2813 ( .A1(_00295_), .A2(_00301_), .ZN(_00053_) );
  AND2_X1 U2814 ( .A1(_00055_), .A2(_00053_), .ZN(_01354_) );
  AND2_X1 U2815 ( .A1(_01354_), .A2(_00294_), .ZN(_00186_) );
  AND2_X1 U2816 ( .A1(_01352__PTR0), .A2(P2_P1_State2_PTR2), .ZN(_00187_) );
  OR2_X1 U2817 ( .A1(_01355__PTR0), .A2(_01355__PTR1), .ZN(_00056_) );
  OR2_X1 U2818 ( .A1(_01357__PTR0), .A2(_01353__PTR1), .ZN(_00058_) );
  AND2_X1 U2819 ( .A1(_00056_), .A2(_00057_), .ZN(_01359__PTR0) );
  AND2_X1 U2820 ( .A1(_01359__PTR0), .A2(_01359__PTR1), .ZN(_01360__PTR0) );
  AND2_X1 U2821 ( .A1(_01360__PTR0), .A2(_01360__PTR1), .ZN(_00188_) );
  OR2_X1 U2822 ( .A1(_00294_), .A2(_02186__PTR32), .ZN(_01355__PTR1) );
  OR2_X1 U2823 ( .A1(_01361__PTR0), .A2(_01355__PTR1), .ZN(_00063_) );
  OR2_X1 U2824 ( .A1(_00145_), .A2(_00081_), .ZN(_00059_) );
  OR2_X1 U2825 ( .A1(_00300_), .A2(_00294_), .ZN(_00060_) );
  OR2_X1 U2826 ( .A1(_00053_), .A2(P2_P1_State2_PTR3), .ZN(_00062_) );
  AND2_X1 U2827 ( .A1(_00063_), .A2(_00057_), .ZN(_01362__PTR0) );
  AND2_X1 U2828 ( .A1(_01362__PTR0), .A2(_01359__PTR1), .ZN(_01363__PTR0) );
  AND2_X1 U2829 ( .A1(_01363__PTR0), .A2(_01360__PTR1), .ZN(_00189_) );
  OR2_X1 U2830 ( .A1(_01364__PTR0), .A2(_01355__PTR1), .ZN(_00064_) );
  OR2_X1 U2831 ( .A1(_00300_), .A2(_00295_), .ZN(_00145_) );
  AND2_X1 U2832 ( .A1(_00064_), .A2(_00057_), .ZN(_01365__PTR0) );
  AND2_X1 U2833 ( .A1(_01365__PTR0), .A2(_01359__PTR1), .ZN(_01366__PTR0) );
  AND2_X1 U2834 ( .A1(_01366__PTR0), .A2(_01360__PTR1), .ZN(_00190_) );
  OR2_X1 U2835 ( .A1(_01367__PTR0), .A2(_01355__PTR1), .ZN(_00065_) );
  AND2_X1 U2836 ( .A1(_00065_), .A2(_00057_), .ZN(_01368__PTR0) );
  AND2_X1 U2837 ( .A1(_01369__PTR0), .A2(_01360__PTR1), .ZN(_00191_) );
  OR2_X1 U2838 ( .A1(_01370__PTR0), .A2(_01355__PTR1), .ZN(_00066_) );
  AND2_X1 U2839 ( .A1(_00066_), .A2(_00057_), .ZN(_01371__PTR0) );
  AND2_X1 U2840 ( .A1(_01371__PTR0), .A2(_01359__PTR1), .ZN(_01372__PTR0) );
  AND2_X1 U2841 ( .A1(_01359__PTR2), .A2(_00062_), .ZN(_01360__PTR1) );
  AND2_X1 U2842 ( .A1(_01372__PTR0), .A2(_01360__PTR1), .ZN(_00192_) );
  OR2_X1 U2843 ( .A1(_01373__PTR0), .A2(_01355__PTR1), .ZN(_00067_) );
  OR2_X1 U2844 ( .A1(_01356_), .A2(_01768__PTR2), .ZN(_00057_) );
  OR2_X1 U2845 ( .A1(_00300_), .A2(P2_P1_State2_PTR1), .ZN(_01357__PTR0) );
  OR2_X1 U2846 ( .A1(_00301_), .A2(P2_P1_State2_PTR3), .ZN(_01353__PTR1) );
  AND2_X1 U2847 ( .A1(_01374__PTR0), .A2(_01359__PTR1), .ZN(_01375__PTR0) );
  AND2_X1 U2848 ( .A1(_01375__PTR0), .A2(_01360__PTR1), .ZN(_00193_) );
  OR2_X1 U2849 ( .A1(_01376__PTR0), .A2(_01355__PTR1), .ZN(_00068_) );
  OR2_X1 U2850 ( .A1(_01358_), .A2(P2_P1_State2_PTR3), .ZN(_00061_) );
  AND2_X1 U2851 ( .A1(_00068_), .A2(_00057_), .ZN(_01377__PTR0) );
  AND2_X1 U2852 ( .A1(_00058_), .A2(_00059_), .ZN(_01359__PTR1) );
  AND2_X1 U2853 ( .A1(_00060_), .A2(_00061_), .ZN(_01359__PTR2) );
  AND2_X1 U2854 ( .A1(_01377__PTR0), .A2(_01359__PTR1), .ZN(_01378__PTR0) );
  AND2_X1 U2855 ( .A1(_01378__PTR0), .A2(_01360__PTR1), .ZN(_00194_) );
  OR2_X1 U2856 ( .A1(_01379__PTR0), .A2(_01355__PTR1), .ZN(_00069_) );
  AND2_X1 U2857 ( .A1(_00069_), .A2(_00057_), .ZN(_01380__PTR0) );
  AND2_X1 U2858 ( .A1(_01380__PTR0), .A2(_01359__PTR1), .ZN(_01381__PTR0) );
  AND2_X1 U2859 ( .A1(_01381__PTR0), .A2(_01360__PTR1), .ZN(_00195_) );
  OR2_X1 U2860 ( .A1(_01382__PTR0), .A2(_01355__PTR1), .ZN(_00070_) );
  OR2_X1 U2861 ( .A1(P2_P1_State2_PTR0), .A2(_00294_), .ZN(_01356_) );
  AND2_X1 U2862 ( .A1(_00070_), .A2(_00057_), .ZN(_01383__PTR0) );
  AND2_X1 U2863 ( .A1(_01383__PTR0), .A2(_01359__PTR1), .ZN(_01384__PTR0) );
  AND2_X1 U2864 ( .A1(_01384__PTR0), .A2(_01360__PTR1), .ZN(_00196_) );
  OR2_X1 U2865 ( .A1(_01385__PTR0), .A2(_01355__PTR1), .ZN(_00071_) );
  AND2_X1 U2866 ( .A1(_00071_), .A2(_00057_), .ZN(_01386__PTR0) );
  AND2_X1 U2867 ( .A1(_01386__PTR0), .A2(_01359__PTR1), .ZN(_01387__PTR0) );
  AND2_X1 U2868 ( .A1(_01387__PTR0), .A2(_01360__PTR1), .ZN(_00197_) );
  AND2_X1 U2869 ( .A1(_00072_), .A2(_00057_), .ZN(_01389__PTR0) );
  AND2_X1 U2870 ( .A1(_01389__PTR0), .A2(_01359__PTR1), .ZN(_01390__PTR0) );
  AND2_X1 U2871 ( .A1(_01390__PTR0), .A2(_01360__PTR1), .ZN(_00198_) );
  OR2_X1 U2872 ( .A1(_01391__PTR0), .A2(_01355__PTR1), .ZN(_00073_) );
  AND2_X1 U2873 ( .A1(_00073_), .A2(_00057_), .ZN(_01392__PTR0) );
  AND2_X1 U2874 ( .A1(_01392__PTR0), .A2(_01359__PTR1), .ZN(_01393__PTR0) );
  AND2_X1 U2875 ( .A1(_01393__PTR0), .A2(_01360__PTR1), .ZN(_00199_) );
  OR2_X1 U2876 ( .A1(_01394__PTR0), .A2(_01355__PTR1), .ZN(_00074_) );
  AND2_X1 U2877 ( .A1(_00074_), .A2(_00057_), .ZN(_01395__PTR0) );
  AND2_X1 U2878 ( .A1(_01395__PTR0), .A2(_01359__PTR1), .ZN(_01396__PTR0) );
  AND2_X1 U2879 ( .A1(_01396__PTR0), .A2(_01360__PTR1), .ZN(_00200_) );
  OR2_X1 U2880 ( .A1(_01397__PTR0), .A2(_01355__PTR1), .ZN(_00075_) );
  AND2_X1 U2881 ( .A1(_00075_), .A2(_00057_), .ZN(_01398__PTR0) );
  AND2_X1 U2882 ( .A1(_01398__PTR0), .A2(_01359__PTR1), .ZN(_01399__PTR0) );
  AND2_X1 U2883 ( .A1(_01399__PTR0), .A2(_01360__PTR1), .ZN(_00201_) );
  OR2_X1 U2884 ( .A1(_01400__PTR0), .A2(_01355__PTR1), .ZN(_00076_) );
  AND2_X1 U2885 ( .A1(_00076_), .A2(_00057_), .ZN(_01401__PTR0) );
  AND2_X1 U2886 ( .A1(_01401__PTR0), .A2(_01359__PTR1), .ZN(_01402__PTR0) );
  AND2_X1 U2887 ( .A1(_01402__PTR0), .A2(_01360__PTR1), .ZN(_00202_) );
  OR2_X1 U2888 ( .A1(_01403__PTR0), .A2(_01355__PTR1), .ZN(_00077_) );
  AND2_X1 U2889 ( .A1(_00077_), .A2(_00057_), .ZN(_01404__PTR0) );
  AND2_X1 U2890 ( .A1(_01404__PTR0), .A2(_01359__PTR1), .ZN(_01405__PTR0) );
  AND2_X1 U2891 ( .A1(_01405__PTR0), .A2(_01360__PTR1), .ZN(_00203_) );
  OR2_X1 U2892 ( .A1(P2_P1_Flush), .A2(_00304_), .ZN(_01406__PTR2) );
  OR2_X1 U2893 ( .A1(_00145_), .A2(_01353__PTR1), .ZN(_01407_) );
  OR2_X1 U2894 ( .A1(_01407_), .A2(_01406__PTR2), .ZN(_00079_) );
  AND2_X1 U2895 ( .A1(_00078_), .A2(_00057_), .ZN(_01408__PTR0) );
  AND2_X1 U2896 ( .A1(_00079_), .A2(_00060_), .ZN(_01408__PTR1) );
  AND2_X1 U2897 ( .A1(_01408__PTR0), .A2(_01408__PTR1), .ZN(_01409_) );
  AND2_X1 U2898 ( .A1(_01409_), .A2(_00061_), .ZN(_00204_) );
  AND2_X1 U2899 ( .A1(_00080_), .A2(_00078_), .ZN(_01410__PTR0) );
  AND2_X1 U2900 ( .A1(_00060_), .A2(_00081_), .ZN(_01410__PTR1) );
  AND2_X1 U2901 ( .A1(_01410__PTR0), .A2(_01410__PTR1), .ZN(_00205_) );
  OR2_X1 U2902 ( .A1(_01357__PTR0), .A2(P2_P1_State2_PTR2), .ZN(_00082_) );
  AND2_X1 U2903 ( .A1(_01411__PTR0), .A2(_01411__PTR1), .ZN(_01412_) );
  AND2_X1 U2904 ( .A1(_01412_), .A2(_00294_), .ZN(_00206_) );
  OR2_X1 U2905 ( .A1(_00144_), .A2(_00301_), .ZN(_00051_) );
  OR2_X1 U2906 ( .A1(_00295_), .A2(P2_P1_State2_PTR2), .ZN(_00052_) );
  AND2_X1 U2907 ( .A1(_00051_), .A2(_00052_), .ZN(_01351__PTR0) );
  AND2_X1 U2908 ( .A1(_00053_), .A2(_00294_), .ZN(_01351__PTR1) );
  AND2_X1 U2909 ( .A1(_01351__PTR0), .A2(_01351__PTR1), .ZN(_00184_) );
  AND2_X1 U2910 ( .A1(_00046_), .A2(_00083_), .ZN(_00207_) );
  OR2_X1 U2911 ( .A1(_00144_), .A2(P2_P1_State2_PTR2), .ZN(_00084_) );
  AND2_X1 U2912 ( .A1(_00084_), .A2(_00051_), .ZN(_01413__PTR0) );
  AND2_X1 U2913 ( .A1(_00052_), .A2(_00053_), .ZN(_01411__PTR1) );
  AND2_X1 U2914 ( .A1(_01413__PTR0), .A2(_01411__PTR1), .ZN(_01414_) );
  AND2_X1 U2915 ( .A1(_01414_), .A2(_00294_), .ZN(_00208_) );
  OR2_X1 U2916 ( .A1(_01344__PTR0), .A2(P2_State_PTR2), .ZN(_00085_) );
  OR2_X1 U2917 ( .A1(_01344__PTR0), .A2(_00285_), .ZN(_00086_) );
  OR2_X1 U2918 ( .A1(P2_State_PTR1), .A2(_00285_), .ZN(_00083_) );
  AND2_X1 U2919 ( .A1(_00085_), .A2(_00086_), .ZN(_01415__PTR0) );
  AND2_X1 U2920 ( .A1(_00087_), .A2(_00083_), .ZN(_01415__PTR1) );
  AND2_X1 U2921 ( .A1(_01415__PTR0), .A2(_01415__PTR1), .ZN(_00209_) );
  OR2_X1 U2922 ( .A1(_00305_), .A2(_00286_), .ZN(_01344__PTR0) );
  OR2_X1 U2923 ( .A1(P1_State_PTR2), .A2(_00312_), .ZN(_01416__PTR1) );
  OR2_X1 U2924 ( .A1(_01416__PTR0), .A2(_01416__PTR1), .ZN(_01417_) );
  OR2_X1 U2925 ( .A1(_00303_), .A2(_01894__PTR14), .ZN(_01421__PTR1) );
  OR2_X1 U2926 ( .A1(_01421__PTR0), .A2(_01421__PTR1), .ZN(_00093_) );
  OR2_X1 U2927 ( .A1(_00139_), .A2(_00303_), .ZN(_00094_) );
  AND2_X1 U2928 ( .A1(_00093_), .A2(_00094_), .ZN(_01422_) );
  AND2_X1 U2929 ( .A1(_01422_), .A2(_00296_), .ZN(_00211_) );
  AND2_X1 U2930 ( .A1(_00097_), .A2(_00296_), .ZN(_01423__PTR1) );
  AND2_X1 U2931 ( .A1(_01423__PTR0), .A2(_01423__PTR1), .ZN(_00212_) );
  AND2_X1 U2932 ( .A1(P1_P1_State2_PTR0), .A2(_00297_), .ZN(_01424__PTR0) );
  AND2_X1 U2933 ( .A1(P1_P1_State2_PTR2), .A2(_00296_), .ZN(_01424__PTR1) );
  AND2_X1 U2934 ( .A1(_01424__PTR0), .A2(P1_P1_State2_PTR2), .ZN(_00215_) );
  OR2_X1 U2935 ( .A1(_01433__PTR0), .A2(_01427__PTR1), .ZN(_00107_) );
  AND2_X1 U2936 ( .A1(_01438__PTR0), .A2(_01432__PTR1), .ZN(_00218_) );
  AND2_X1 U2937 ( .A1(_00109_), .A2(_00101_), .ZN(_01440__PTR0) );
  AND2_X1 U2938 ( .A1(_01440__PTR0), .A2(_01431__PTR1), .ZN(_01441__PTR0) );
  AND2_X1 U2939 ( .A1(_00110_), .A2(_00101_), .ZN(_01443__PTR0) );
  AND2_X1 U2940 ( .A1(_01443__PTR0), .A2(_01431__PTR1), .ZN(_01444__PTR0) );
  AND2_X1 U2941 ( .A1(_01444__PTR0), .A2(_01432__PTR1), .ZN(_00220_) );
  AND2_X1 U2942 ( .A1(_00113_), .A2(_00101_), .ZN(_01452__PTR0) );
  AND2_X1 U2943 ( .A1(_01452__PTR0), .A2(_01431__PTR1), .ZN(_01453__PTR0) );
  AND2_X1 U2944 ( .A1(_01453__PTR0), .A2(_01432__PTR1), .ZN(_00223_) );
  OR2_X1 U2945 ( .A1(_01454__PTR0), .A2(_01427__PTR1), .ZN(_00114_) );
  AND2_X1 U2946 ( .A1(_00114_), .A2(_00101_), .ZN(_01455__PTR0) );
  AND2_X1 U2947 ( .A1(_01455__PTR0), .A2(_01431__PTR1), .ZN(_01456__PTR0) );
  AND2_X1 U2948 ( .A1(_01456__PTR0), .A2(_01432__PTR1), .ZN(_00224_) );
  OR2_X1 U2949 ( .A1(_01457__PTR0), .A2(_01427__PTR1), .ZN(_00115_) );
  AND2_X1 U2950 ( .A1(_00115_), .A2(_00101_), .ZN(_01458__PTR0) );
  AND2_X1 U2951 ( .A1(_01458__PTR0), .A2(_01431__PTR1), .ZN(_01459__PTR0) );
  AND2_X1 U2952 ( .A1(_01459__PTR0), .A2(_01432__PTR1), .ZN(_00225_) );
  OR2_X1 U2953 ( .A1(_01460__PTR0), .A2(_01427__PTR1), .ZN(_00116_) );
  AND2_X1 U2954 ( .A1(_00116_), .A2(_00101_), .ZN(_01461__PTR0) );
  AND2_X1 U2955 ( .A1(_01461__PTR0), .A2(_01431__PTR1), .ZN(_01462__PTR0) );
  AND2_X1 U2956 ( .A1(_01462__PTR0), .A2(_01432__PTR1), .ZN(_00226_) );
  OR2_X1 U2957 ( .A1(_01463__PTR0), .A2(_01427__PTR1), .ZN(_00117_) );
  AND2_X1 U2958 ( .A1(_00117_), .A2(_00101_), .ZN(_01464__PTR0) );
  AND2_X1 U2959 ( .A1(_01464__PTR0), .A2(_01431__PTR1), .ZN(_01465__PTR0) );
  AND2_X1 U2960 ( .A1(_01465__PTR0), .A2(_01432__PTR1), .ZN(_00227_) );
  AND2_X1 U2961 ( .A1(_00119_), .A2(_00101_), .ZN(_01470__PTR0) );
  OR2_X1 U2962 ( .A1(_01475__PTR0), .A2(_01427__PTR1), .ZN(_00121_) );
  OR2_X1 U2963 ( .A1(_01428_), .A2(_01770__PTR2), .ZN(_00101_) );
  OR2_X1 U2964 ( .A1(_01429__PTR0), .A2(_01425__PTR1), .ZN(_00102_) );
  AND2_X1 U2965 ( .A1(_00121_), .A2(_00101_), .ZN(_01476__PTR0) );
  AND2_X1 U2966 ( .A1(_01476__PTR0), .A2(_01431__PTR1), .ZN(_01477__PTR0) );
  AND2_X1 U2967 ( .A1(_01477__PTR0), .A2(_01432__PTR1), .ZN(_00231_) );
  OR2_X1 U2968 ( .A1(_01430_), .A2(P1_P1_State2_PTR3), .ZN(_00105_) );
  AND2_X1 U2969 ( .A1(_00122_), .A2(_00101_), .ZN(_01480__PTR0) );
  AND2_X1 U2970 ( .A1(_00123_), .A2(_00104_), .ZN(_01480__PTR1) );
  AND2_X1 U2971 ( .A1(_01481_), .A2(_00105_), .ZN(_00232_) );
  AND2_X1 U2972 ( .A1(_00124_), .A2(_00122_), .ZN(_01482__PTR0) );
  AND2_X1 U2973 ( .A1(_00104_), .A2(_00125_), .ZN(_01482__PTR1) );
  AND2_X1 U2974 ( .A1(_01482__PTR0), .A2(_01482__PTR1), .ZN(_00233_) );
  AND2_X1 U2975 ( .A1(_00095_), .A2(_00096_), .ZN(_01423__PTR0) );
  AND2_X1 U2976 ( .A1(_00090_), .A2(_00127_), .ZN(_00235_) );
  OR2_X1 U2977 ( .A1(_00138_), .A2(P1_P1_State2_PTR2), .ZN(_00128_) );
  AND2_X1 U2978 ( .A1(_00128_), .A2(_00095_), .ZN(_01485__PTR0) );
  AND2_X1 U2979 ( .A1(_01485__PTR0), .A2(_01483__PTR1), .ZN(_01486_) );
  AND2_X1 U2980 ( .A1(_01486_), .A2(_00296_), .ZN(_00236_) );
  AND2_X1 U2981 ( .A1(_00124_), .A2(_00132_), .ZN(_01489__PTR0) );
  AND2_X1 U2982 ( .A1(_00133_), .A2(_00103_), .ZN(_01489__PTR1) );
  AND2_X1 U2983 ( .A1(_01489__PTR0), .A2(_01489__PTR1), .ZN(_01490_) );
  AND2_X1 U2984 ( .A1(_01490_), .A2(_00106_), .ZN(_00238_) );
  OR2_X1 U2985 ( .A1(_00138_), .A2(_01425__PTR1), .ZN(_00124_) );
  OR2_X1 U2986 ( .A1(_01488_), .A2(_01894__PTR9), .ZN(_00132_) );
  OR2_X1 U2987 ( .A1(_01429__PTR0), .A2(_00125_), .ZN(_00133_) );
  OR2_X1 U2988 ( .A1(P1_P1_State2_PTR0), .A2(_00297_), .ZN(_01421__PTR0) );
  OR2_X1 U2989 ( .A1(_01421__PTR0), .A2(_00125_), .ZN(_01488_) );
  AND2_X1 U2990 ( .A1(_01424__PTR0), .A2(_01424__PTR1), .ZN(_00213_) );
  AND2_X1 U2991 ( .A1(_00138_), .A2(_00139_), .ZN(_01491__PTR0) );
  AND2_X1 U2992 ( .A1(_01491__PTR0), .A2(_01424__PTR1), .ZN(_00239_) );
  OR2_X1 U2993 ( .A1(_01419_), .A2(P1_State_PTR2), .ZN(_00090_) );
  OR2_X1 U2994 ( .A1(_00311_), .A2(P1_State_PTR1), .ZN(_01419_) );
  OR2_X1 U2995 ( .A1(_01419_), .A2(_00275_), .ZN(_00091_) );
  AND2_X1 U2996 ( .A1(_00089_), .A2(_00090_), .ZN(_01420__PTR0) );
  AND2_X1 U2997 ( .A1(_00091_), .A2(_00092_), .ZN(_01420__PTR1) );
  AND2_X1 U2998 ( .A1(_01420__PTR0), .A2(_01420__PTR1), .ZN(_00210_) );
  OR2_X1 U2999 ( .A1(_00276_), .A2(_00275_), .ZN(_00092_) );
  AND2_X1 U3000 ( .A1(_00089_), .A2(_00092_), .ZN(_00240_) );
  OR2_X1 U3001 ( .A1(_01417_), .A2(_01769__PTR4), .ZN(_00088_) );
  OR2_X1 U3002 ( .A1(_00311_), .A2(_00276_), .ZN(_01416__PTR0) );
  OR2_X1 U3003 ( .A1(_01416__PTR0), .A2(P1_State_PTR2), .ZN(_00129_) );
  OR2_X1 U3004 ( .A1(_01416__PTR0), .A2(_00275_), .ZN(_00130_) );
  OR2_X1 U3005 ( .A1(P1_State_PTR1), .A2(_00275_), .ZN(_00127_) );
  AND2_X1 U3006 ( .A1(_00129_), .A2(_00130_), .ZN(_01487__PTR0) );
  OR2_X1 U3007 ( .A1(P1_State_PTR1), .A2(P1_State_PTR2), .ZN(_00131_) );
  AND2_X1 U3008 ( .A1(_00131_), .A2(_00127_), .ZN(_01487__PTR1) );
  AND2_X1 U3009 ( .A1(_01487__PTR0), .A2(_01487__PTR1), .ZN(_00237_) );
  OR2_X1 U3010 ( .A1(P1_P1_State2_PTR0), .A2(P1_P1_State2_PTR1), .ZN(_00138_) );
  OR2_X1 U3011 ( .A1(P1_P1_State2_PTR2), .A2(_01894__PTR9), .ZN(_01492__PTR1) );
  OR2_X1 U3012 ( .A1(_01421__PTR0), .A2(_01492__PTR1), .ZN(_00140_) );
  AND2_X1 U3013 ( .A1(_00140_), .A2(_00099_), .ZN(_01493__PTR0) );
  AND2_X1 U3014 ( .A1(_01493__PTR0), .A2(_01423__PTR1), .ZN(_00241_) );
  AND2_X1 U3015 ( .A1(_01426_), .A2(_00296_), .ZN(_00214_) );
  OR2_X1 U3016 ( .A1(_00139_), .A2(P1_P1_State2_PTR2), .ZN(_00099_) );
  AND2_X1 U3017 ( .A1(_00099_), .A2(_00097_), .ZN(_01426_) );
  OR2_X1 U3018 ( .A1(_00138_), .A2(_00303_), .ZN(_00095_) );
  OR2_X1 U3019 ( .A1(_01429__PTR0), .A2(P1_P1_State2_PTR2), .ZN(_00126_) );
  OR2_X1 U3020 ( .A1(_00297_), .A2(P1_P1_State2_PTR2), .ZN(_00096_) );
  AND2_X1 U3021 ( .A1(_00095_), .A2(_00126_), .ZN(_01483__PTR0) );
  AND2_X1 U3022 ( .A1(_00096_), .A2(_00097_), .ZN(_01483__PTR1) );
  AND2_X1 U3023 ( .A1(_01483__PTR0), .A2(_01483__PTR1), .ZN(_01484_) );
  AND2_X1 U3024 ( .A1(_01484_), .A2(_00296_), .ZN(_00234_) );
  OR2_X1 U3025 ( .A1(P1_P1_Flush), .A2(_00310_), .ZN(_01478__PTR2) );
  OR2_X1 U3026 ( .A1(_00139_), .A2(_01425__PTR1), .ZN(_01479_) );
  OR2_X1 U3027 ( .A1(_01479_), .A2(_01478__PTR2), .ZN(_00123_) );
  OR2_X1 U3028 ( .A1(P1_P1_State2_PTR1), .A2(_00303_), .ZN(_01494_) );
  OR2_X1 U3029 ( .A1(_01494_), .A2(P1_P1_State2_PTR3), .ZN(_00141_) );
  OR2_X1 U3030 ( .A1(P1_P1_State2_PTR2), .A2(P1_P1_State2_PTR3), .ZN(_00125_) );
  AND2_X1 U3031 ( .A1(_00141_), .A2(_00125_), .ZN(_01495__PTR2) );
  AND2_X1 U3032 ( .A1(_01480__PTR0), .A2(_01480__PTR1), .ZN(_01481_) );
  AND2_X1 U3033 ( .A1(_01481_), .A2(_01495__PTR2), .ZN(_00242_) );
  OR2_X1 U3034 ( .A1(P1_P1_State2_PTR1), .A2(P1_P1_State2_PTR2), .ZN(_01430_) );
  AND2_X1 U3035 ( .A1(_01480__PTR0), .A2(_01431__PTR1), .ZN(_01496__PTR0) );
  AND2_X1 U3036 ( .A1(_01480__PTR1), .A2(_00105_), .ZN(_01496__PTR1) );
  AND2_X1 U3037 ( .A1(_01496__PTR0), .A2(_01496__PTR1), .ZN(_00243_) );
  OR2_X1 U3038 ( .A1(_01835__PTR0), .A2(P1_P1_State2_PTR0), .ZN(_01475__PTR0) );
  OR2_X1 U3039 ( .A1(_01835__PTR1), .A2(P1_P1_State2_PTR0), .ZN(_01454__PTR0) );
  OR2_X1 U3040 ( .A1(_01835__PTR2), .A2(P1_P1_State2_PTR0), .ZN(_01457__PTR0) );
  OR2_X1 U3041 ( .A1(_01835__PTR3), .A2(P1_P1_State2_PTR0), .ZN(_01460__PTR0) );
  OR2_X1 U3042 ( .A1(_01835__PTR4), .A2(P1_P1_State2_PTR0), .ZN(_01463__PTR0) );
  OR2_X1 U3043 ( .A1(_01835__PTR5), .A2(P1_P1_State2_PTR0), .ZN(_01466__PTR0) );
  OR2_X1 U3044 ( .A1(_00297_), .A2(_00303_), .ZN(_00097_) );
  OR2_X1 U3045 ( .A1(_00097_), .A2(P1_P1_State2_PTR3), .ZN(_00106_) );
  AND2_X1 U3046 ( .A1(_00118_), .A2(_00101_), .ZN(_01467__PTR0) );
  AND2_X1 U3047 ( .A1(_01467__PTR0), .A2(_01431__PTR1), .ZN(_01468__PTR0) );
  AND2_X1 U3048 ( .A1(_01431__PTR2), .A2(_00106_), .ZN(_01432__PTR1) );
  AND2_X1 U3049 ( .A1(_01468__PTR0), .A2(_01432__PTR1), .ZN(_00228_) );
  OR2_X1 U3050 ( .A1(_00296_), .A2(_01894__PTR32), .ZN(_01427__PTR1) );
  OR2_X1 U3051 ( .A1(_01466__PTR0), .A2(_01427__PTR1), .ZN(_00118_) );
  OR2_X1 U3052 ( .A1(P1_P1_State2_PTR0), .A2(_00296_), .ZN(_01428_) );
  OR2_X1 U3053 ( .A1(_00302_), .A2(P1_P1_State2_PTR1), .ZN(_01429__PTR0) );
  OR2_X1 U3054 ( .A1(_00303_), .A2(P1_P1_State2_PTR3), .ZN(_01425__PTR1) );
  OR2_X1 U3055 ( .A1(_00302_), .A2(_00297_), .ZN(_00139_) );
  OR2_X1 U3056 ( .A1(_00139_), .A2(_00125_), .ZN(_00103_) );
  OR2_X1 U3057 ( .A1(_00302_), .A2(_00296_), .ZN(_00104_) );
  AND2_X1 U3058 ( .A1(_00102_), .A2(_00103_), .ZN(_01431__PTR1) );
  AND2_X1 U3059 ( .A1(_00104_), .A2(_00105_), .ZN(_01431__PTR2) );
  OR2_X1 U3060 ( .A1(_01835__PTR6), .A2(P1_P1_State2_PTR0), .ZN(_01469__PTR0) );
  OR2_X1 U3061 ( .A1(_01469__PTR0), .A2(_01427__PTR1), .ZN(_00119_) );
  AND2_X1 U3062 ( .A1(_01470__PTR0), .A2(_01431__PTR1), .ZN(_01471__PTR0) );
  AND2_X1 U3063 ( .A1(_01471__PTR0), .A2(_01432__PTR1), .ZN(_00229_) );
  OR2_X1 U3064 ( .A1(_01835__PTR7), .A2(P1_P1_State2_PTR0), .ZN(_01472__PTR0) );
  OR2_X1 U3065 ( .A1(_01472__PTR0), .A2(_01427__PTR1), .ZN(_00120_) );
  AND2_X1 U3066 ( .A1(_00120_), .A2(_00101_), .ZN(_01473__PTR0) );
  AND2_X1 U3067 ( .A1(_01473__PTR0), .A2(_01431__PTR1), .ZN(_01474__PTR0) );
  AND2_X1 U3068 ( .A1(_01474__PTR0), .A2(_01432__PTR1), .ZN(_00230_) );
  OR2_X1 U3069 ( .A1(_01835__PTR8), .A2(P1_P1_State2_PTR0), .ZN(_01427__PTR0) );
  OR2_X1 U3070 ( .A1(_01427__PTR0), .A2(_01427__PTR1), .ZN(_00100_) );
  AND2_X1 U3071 ( .A1(_00100_), .A2(_00101_), .ZN(_01431__PTR0) );
  AND2_X1 U3072 ( .A1(_01431__PTR0), .A2(_01431__PTR1), .ZN(_01432__PTR0) );
  AND2_X1 U3073 ( .A1(_01432__PTR0), .A2(_01432__PTR1), .ZN(_00216_) );
  OR2_X1 U3074 ( .A1(_01835__PTR9), .A2(P1_P1_State2_PTR0), .ZN(_01433__PTR0) );
  AND2_X1 U3075 ( .A1(_00107_), .A2(_00101_), .ZN(_01434__PTR0) );
  AND2_X1 U3076 ( .A1(_01434__PTR0), .A2(_01431__PTR1), .ZN(_01435__PTR0) );
  AND2_X1 U3077 ( .A1(_01435__PTR0), .A2(_01432__PTR1), .ZN(_00217_) );
  OR2_X1 U3078 ( .A1(_01835__PTR10), .A2(P1_P1_State2_PTR0), .ZN(_01436__PTR0) );
  OR2_X1 U3079 ( .A1(_01436__PTR0), .A2(_01427__PTR1), .ZN(_00108_) );
  AND2_X1 U3080 ( .A1(_00108_), .A2(_00101_), .ZN(_01437__PTR0) );
  AND2_X1 U3081 ( .A1(_01437__PTR0), .A2(_01431__PTR1), .ZN(_01438__PTR0) );
  OR2_X1 U3082 ( .A1(_01835__PTR11), .A2(P1_P1_State2_PTR0), .ZN(_01439__PTR0) );
  OR2_X1 U3083 ( .A1(_01439__PTR0), .A2(_01427__PTR1), .ZN(_00109_) );
  AND2_X1 U3084 ( .A1(_01441__PTR0), .A2(_01432__PTR1), .ZN(_00219_) );
  OR2_X1 U3085 ( .A1(_01835__PTR12), .A2(P1_P1_State2_PTR0), .ZN(_01442__PTR0) );
  OR2_X1 U3086 ( .A1(_01442__PTR0), .A2(_01427__PTR1), .ZN(_00110_) );
  OR2_X1 U3087 ( .A1(_01835__PTR13), .A2(P1_P1_State2_PTR0), .ZN(_01445__PTR0) );
  OR2_X1 U3088 ( .A1(_01445__PTR0), .A2(_01427__PTR1), .ZN(_00111_) );
  AND2_X1 U3089 ( .A1(_00111_), .A2(_00101_), .ZN(_01446__PTR0) );
  AND2_X1 U3090 ( .A1(_01446__PTR0), .A2(_01431__PTR1), .ZN(_01447__PTR0) );
  AND2_X1 U3091 ( .A1(_01447__PTR0), .A2(_01432__PTR1), .ZN(_00221_) );
  OR2_X1 U3092 ( .A1(_01835__PTR14), .A2(P1_P1_State2_PTR0), .ZN(_01448__PTR0) );
  OR2_X1 U3093 ( .A1(_01448__PTR0), .A2(_01427__PTR1), .ZN(_00112_) );
  AND2_X1 U3094 ( .A1(_00112_), .A2(_00101_), .ZN(_01449__PTR0) );
  AND2_X1 U3095 ( .A1(_01449__PTR0), .A2(_01431__PTR1), .ZN(_01450__PTR0) );
  AND2_X1 U3096 ( .A1(_01450__PTR0), .A2(_01432__PTR1), .ZN(_00222_) );
  OR2_X1 U3097 ( .A1(_01835__PTR15), .A2(P1_P1_State2_PTR0), .ZN(_01451__PTR0) );
  OR2_X1 U3098 ( .A1(_01451__PTR0), .A2(_01427__PTR1), .ZN(_00113_) );
  OR2_X1 U3099 ( .A1(_01421__PTR0), .A2(_01425__PTR1), .ZN(_00122_) );
  OR2_X1 U3100 ( .A1(_00122_), .A2(_01894__PTR14), .ZN(_00098_) );
  OR2_X1 U3101 ( .A1(P2_P1_State2_PTR0), .A2(P2_P1_State2_PTR1), .ZN(_00144_) );
  OR2_X1 U3102 ( .A1(_00144_), .A2(_01353__PTR1), .ZN(_00080_) );
  OR2_X1 U3103 ( .A1(P2_P1_State2_PTR2), .A2(P2_P1_State2_PTR3), .ZN(_00081_) );
  OR2_X1 U3104 ( .A1(_01349__PTR0), .A2(_00081_), .ZN(_01497_) );
  OR2_X1 U3105 ( .A1(_01497_), .A2(_02186__PTR9), .ZN(_00142_) );
  OR2_X1 U3106 ( .A1(_01357__PTR0), .A2(_00081_), .ZN(_00143_) );
  AND2_X1 U3107 ( .A1(_00080_), .A2(_00142_), .ZN(_01498__PTR0) );
  AND2_X1 U3108 ( .A1(_00143_), .A2(_00059_), .ZN(_01498__PTR1) );
  AND2_X1 U3109 ( .A1(_01498__PTR0), .A2(_01498__PTR1), .ZN(_01499_) );
  AND2_X1 U3110 ( .A1(_01499_), .A2(_00062_), .ZN(_00244_) );
  AND2_X1 U3111 ( .A1(_00144_), .A2(_00145_), .ZN(_01500__PTR0) );
  AND2_X1 U3112 ( .A1(_01500__PTR0), .A2(_01352__PTR1), .ZN(_00245_) );
  OR2_X1 U3113 ( .A1(_00305_), .A2(P2_State_PTR1), .ZN(_01347_) );
  OR2_X1 U3114 ( .A1(_01347_), .A2(P2_State_PTR2), .ZN(_00046_) );
  OR2_X1 U3115 ( .A1(_01347_), .A2(_00285_), .ZN(_00047_) );
  OR2_X1 U3116 ( .A1(_00286_), .A2(_00285_), .ZN(_00048_) );
  AND2_X1 U3117 ( .A1(_00045_), .A2(_00046_), .ZN(_01348__PTR0) );
  AND2_X1 U3118 ( .A1(_00047_), .A2(_00048_), .ZN(_01348__PTR1) );
  AND2_X1 U3119 ( .A1(_01348__PTR0), .A2(_01348__PTR1), .ZN(_00182_) );
  AND2_X1 U3120 ( .A1(_00045_), .A2(_00048_), .ZN(_00246_) );
  OR2_X1 U3121 ( .A1(P2_State_PTR2), .A2(_00309_), .ZN(_01344__PTR1) );
  OR2_X1 U3122 ( .A1(_01344__PTR0), .A2(_01344__PTR1), .ZN(_01345_) );
  OR2_X1 U3123 ( .A1(_01345_), .A2(_01767__PTR4), .ZN(_00044_) );
  OR2_X1 U3124 ( .A1(P2_State_PTR1), .A2(P2_State_PTR2), .ZN(_00087_) );
  OR2_X1 U3125 ( .A1(P2_P1_State2_PTR2), .A2(_02186__PTR9), .ZN(_01501__PTR1) );
  OR2_X1 U3126 ( .A1(_01349__PTR0), .A2(_01501__PTR1), .ZN(_00146_) );
  AND2_X1 U3127 ( .A1(_00146_), .A2(_00055_), .ZN(_01502__PTR0) );
  AND2_X1 U3128 ( .A1(_01502__PTR0), .A2(_01351__PTR1), .ZN(_00247_) );
  AND2_X1 U3129 ( .A1(_00051_), .A2(_00082_), .ZN(_01411__PTR0) );
  OR2_X1 U3130 ( .A1(P2_P1_State2_PTR1), .A2(_00301_), .ZN(_01503_) );
  OR2_X1 U3131 ( .A1(_01503_), .A2(P2_P1_State2_PTR3), .ZN(_00147_) );
  AND2_X1 U3132 ( .A1(_00147_), .A2(_00081_), .ZN(_01504__PTR2) );
  AND2_X1 U3133 ( .A1(_01409_), .A2(_01504__PTR2), .ZN(_00248_) );
  OR2_X1 U3134 ( .A1(P2_P1_State2_PTR1), .A2(P2_P1_State2_PTR2), .ZN(_01358_) );
  AND2_X1 U3135 ( .A1(_01408__PTR0), .A2(_01359__PTR1), .ZN(_01505__PTR0) );
  AND2_X1 U3136 ( .A1(_01408__PTR1), .A2(_00061_), .ZN(_01505__PTR1) );
  AND2_X1 U3137 ( .A1(_01505__PTR0), .A2(_01505__PTR1), .ZN(_00249_) );
  OR2_X1 U3138 ( .A1(_02128__PTR0), .A2(P2_P1_State2_PTR0), .ZN(_01403__PTR0) );
  OR2_X1 U3139 ( .A1(_02128__PTR1), .A2(P2_P1_State2_PTR0), .ZN(_01382__PTR0) );
  OR2_X1 U3140 ( .A1(_02128__PTR2), .A2(P2_P1_State2_PTR0), .ZN(_01385__PTR0) );
  OR2_X1 U3141 ( .A1(_02128__PTR3), .A2(P2_P1_State2_PTR0), .ZN(_01388__PTR0) );
  OR2_X1 U3142 ( .A1(_01388__PTR0), .A2(_01355__PTR1), .ZN(_00072_) );
  OR2_X1 U3143 ( .A1(_02128__PTR4), .A2(P2_P1_State2_PTR0), .ZN(_01391__PTR0) );
  OR2_X1 U3144 ( .A1(_02128__PTR5), .A2(P2_P1_State2_PTR0), .ZN(_01394__PTR0) );
  OR2_X1 U3145 ( .A1(_02128__PTR6), .A2(P2_P1_State2_PTR0), .ZN(_01397__PTR0) );
  OR2_X1 U3146 ( .A1(_02128__PTR7), .A2(P2_P1_State2_PTR0), .ZN(_01400__PTR0) );
  OR2_X1 U3147 ( .A1(_02128__PTR8), .A2(P2_P1_State2_PTR0), .ZN(_01355__PTR0) );
  OR2_X1 U3148 ( .A1(_02128__PTR9), .A2(P2_P1_State2_PTR0), .ZN(_01361__PTR0) );
  OR2_X1 U3149 ( .A1(_02128__PTR10), .A2(P2_P1_State2_PTR0), .ZN(_01364__PTR0) );
  OR2_X1 U3150 ( .A1(_02128__PTR11), .A2(P2_P1_State2_PTR0), .ZN(_01367__PTR0) );
  AND2_X1 U3151 ( .A1(_01368__PTR0), .A2(_01359__PTR1), .ZN(_01369__PTR0) );
  OR2_X1 U3152 ( .A1(_02128__PTR12), .A2(P2_P1_State2_PTR0), .ZN(_01370__PTR0) );
  OR2_X1 U3153 ( .A1(_02128__PTR13), .A2(P2_P1_State2_PTR0), .ZN(_01373__PTR0) );
  OR2_X1 U3154 ( .A1(_01855__PTR1), .A2(_02086__PTR4), .ZN(_01507__PTR2) );
  AND2_X1 U3155 ( .A1(_00067_), .A2(_00057_), .ZN(_01374__PTR0) );
  OR2_X1 U3156 ( .A1(_01507__PTR2), .A2(_01507__PTR3), .ZN(_01508__PTR1) );
  OR2_X1 U3157 ( .A1(_01508__PTR0), .A2(_01508__PTR1), .ZN(_01509_) );
  OR2_X1 U3158 ( .A1(_02128__PTR14), .A2(P2_P1_State2_PTR0), .ZN(_01376__PTR0) );
  OR2_X1 U3159 ( .A1(_01509_), .A2(_01506__PTR8), .ZN(_02120__PTR0) );
  OR2_X1 U3160 ( .A1(_02054_), .A2(_02090__PTR3), .ZN(_01510__PTR3) );
  OR2_X1 U3161 ( .A1(_02128__PTR15), .A2(P2_P1_State2_PTR0), .ZN(_01379__PTR0) );
  OR2_X1 U3162 ( .A1(_01506__PTR2), .A2(_01510__PTR3), .ZN(_01511__PTR1) );
  OR2_X1 U3163 ( .A1(P3_P1_State2_PTR0), .A2(P3_P1_State2_PTR1), .ZN(_00150_) );
  OR2_X1 U3164 ( .A1(_00150_), .A2(_01281__PTR1), .ZN(_00036_) );
  OR2_X1 U3165 ( .A1(P3_P1_State2_PTR2), .A2(P3_P1_State2_PTR3), .ZN(_00037_) );
  OR2_X1 U3166 ( .A1(_01277__PTR0), .A2(_00037_), .ZN(_01512_) );
  OR2_X1 U3167 ( .A1(_01512_), .A2(_02475__PTR9), .ZN(_00148_) );
  OR2_X1 U3168 ( .A1(_01285__PTR0), .A2(_00037_), .ZN(_00149_) );
  OR2_X1 U3169 ( .A1(_01510__PTR4), .A2(_01510__PTR5), .ZN(_01511__PTR2) );
  AND2_X1 U3170 ( .A1(_00036_), .A2(_00148_), .ZN(_01513__PTR0) );
  AND2_X1 U3171 ( .A1(_00149_), .A2(_00015_), .ZN(_01513__PTR1) );
  AND2_X1 U3172 ( .A1(_01513__PTR0), .A2(_01513__PTR1), .ZN(_01514_) );
  AND2_X1 U3173 ( .A1(_01514_), .A2(_00018_), .ZN(_00250_) );
  OR2_X1 U3174 ( .A1(_01507__PTR0), .A2(_01511__PTR1), .ZN(_01515__PTR0) );
  OR2_X1 U3175 ( .A1(_01511__PTR2), .A2(_01511__PTR3), .ZN(_01515__PTR1) );
  OR2_X1 U3176 ( .A1(_01515__PTR0), .A2(_01515__PTR1), .ZN(_01516_) );
  OR2_X1 U3177 ( .A1(_01516_), .A2(_02050_), .ZN(_02116__PTR0) );
  OR2_X1 U3178 ( .A1(_02387__PTR1), .A2(_02344_), .ZN(_01517__PTR1) );
  OR2_X1 U3179 ( .A1(_02343_), .A2(_02342_), .ZN(_01517__PTR2) );
  OR2_X1 U3180 ( .A1(_01517__PTR0), .A2(_01517__PTR1), .ZN(_01518__PTR0) );
  OR2_X1 U3181 ( .A1(_01517__PTR2), .A2(_01517__PTR3), .ZN(_01518__PTR1) );
  OR2_X1 U3182 ( .A1(_01518__PTR0), .A2(_01518__PTR1), .ZN(_01519_) );
  OR2_X1 U3183 ( .A1(_01519_), .A2(_02339_), .ZN(_02375__PTR0) );
  OR2_X1 U3184 ( .A1(_02090__PTR3), .A2(_02102__PTR2), .ZN(_01520__PTR4) );
  AND2_X1 U3185 ( .A1(_00150_), .A2(_00151_), .ZN(_01522__PTR0) );
  AND2_X1 U3186 ( .A1(_01522__PTR0), .A2(_01280__PTR1), .ZN(_00251_) );
  OR2_X1 U3187 ( .A1(_01520__PTR4), .A2(_01510__PTR5), .ZN(_01521__PTR2) );
  OR2_X1 U3188 ( .A1(_01521__PTR2), .A2(_01511__PTR3), .ZN(_01523__PTR1) );
  OR2_X1 U3189 ( .A1(_01508__PTR0), .A2(_01523__PTR1), .ZN(_01524_) );
  OR2_X1 U3190 ( .A1(_01524_), .A2(_02050_), .ZN(_02109__PTR0) );
  AND2_X1 U3191 ( .A1(_00001_), .A2(_00004_), .ZN(_00252_) );
  OR2_X1 U3192 ( .A1(_01272__PTR0), .A2(P3_State_PTR2), .ZN(_00041_) );
  OR2_X1 U3193 ( .A1(_01272__PTR0), .A2(_00287_), .ZN(_00042_) );
  OR2_X1 U3194 ( .A1(P3_State_PTR1), .A2(P3_State_PTR2), .ZN(_00043_) );
  AND2_X1 U3195 ( .A1(_00041_), .A2(_00042_), .ZN(_01343__PTR0) );
  AND2_X1 U3196 ( .A1(_00043_), .A2(_00039_), .ZN(_01343__PTR1) );
  AND2_X1 U3197 ( .A1(_01343__PTR0), .A2(_01343__PTR1), .ZN(_00181_) );
  OR2_X1 U3198 ( .A1(_02054_), .A2(_02102__PTR2), .ZN(_01525__PTR3) );
  OR2_X1 U3199 ( .A1(_01506__PTR2), .A2(_01525__PTR3), .ZN(_01526__PTR1) );
  OR2_X1 U3200 ( .A1(_01510__PTR5), .A2(_01510__PTR6), .ZN(_01526__PTR2) );
  OR2_X1 U3201 ( .A1(P3_P1_State2_PTR2), .A2(_02475__PTR9), .ZN(_01527__PTR1) );
  OR2_X1 U3202 ( .A1(_01277__PTR0), .A2(_01527__PTR1), .ZN(_00152_) );
  AND2_X1 U3203 ( .A1(_00152_), .A2(_00011_), .ZN(_01528__PTR0) );
  AND2_X1 U3204 ( .A1(_01528__PTR0), .A2(_01279__PTR1), .ZN(_00253_) );
  OR2_X1 U3205 ( .A1(_01507__PTR0), .A2(_01526__PTR1), .ZN(_01529__PTR0) );
  OR2_X1 U3206 ( .A1(_01526__PTR2), .A2(_01526__PTR3), .ZN(_01529__PTR1) );
  OR2_X1 U3207 ( .A1(_01529__PTR0), .A2(_01529__PTR1), .ZN(_01863__PTR3) );
  OR2_X1 U3208 ( .A1(_02058_), .A2(_02098__PTR1), .ZN(_01530__PTR0) );
  OR2_X1 U3209 ( .A1(_01530__PTR0), .A2(_02086__PTR1), .ZN(_01531__PTR0) );
  OR2_X1 U3210 ( .A1(_01870__PTR1), .A2(_01510__PTR5), .ZN(_01531__PTR2) );
  OR2_X1 U3211 ( .A1(_01510__PTR6), .A2(_01510__PTR7), .ZN(_01511__PTR3) );
  OR2_X1 U3212 ( .A1(_01531__PTR0), .A2(_01531__PTR1), .ZN(_01532__PTR0) );
  OR2_X1 U3213 ( .A1(_01531__PTR2), .A2(_01511__PTR3), .ZN(_01532__PTR1) );
  OR2_X1 U3214 ( .A1(_01532__PTR0), .A2(_01532__PTR1), .ZN(_01533_) );
  OR2_X1 U3215 ( .A1(P3_P1_State2_PTR1), .A2(_00299_), .ZN(_01534_) );
  OR2_X1 U3216 ( .A1(_01534_), .A2(P3_P1_State2_PTR3), .ZN(_00153_) );
  AND2_X1 U3217 ( .A1(_00153_), .A2(_00037_), .ZN(_01535__PTR2) );
  AND2_X1 U3218 ( .A1(_01337_), .A2(_01535__PTR2), .ZN(_00254_) );
  OR2_X1 U3219 ( .A1(_01533_), .A2(_02050_), .ZN(_02102__PTR0) );
  OR2_X1 U3220 ( .A1(P3_P1_State2_PTR1), .A2(P3_P1_State2_PTR2), .ZN(_01286_) );
  OR2_X1 U3221 ( .A1(_01286_), .A2(P3_P1_State2_PTR3), .ZN(_00017_) );
  AND2_X1 U3222 ( .A1(_01336__PTR0), .A2(_01287__PTR1), .ZN(_01536__PTR0) );
  AND2_X1 U3223 ( .A1(_01336__PTR1), .A2(_00017_), .ZN(_01536__PTR1) );
  AND2_X1 U3224 ( .A1(_01536__PTR0), .A2(_01536__PTR1), .ZN(_00255_) );
  OR2_X1 U3225 ( .A1(_01863__PTR0), .A2(_01863__PTR2), .ZN(_01855__PTR0) );
  OR2_X1 U3226 ( .A1(_02417__PTR0), .A2(P3_P1_State2_PTR0), .ZN(_01331__PTR0) );
  OR2_X1 U3227 ( .A1(_02102__PTR2), .A2(_02053_), .ZN(_01537__PTR4) );
  OR2_X1 U3228 ( .A1(_02052_), .A2(_01855__PTR2), .ZN(_01510__PTR6) );
  OR2_X1 U3229 ( .A1(_01855__PTR3), .A2(_02051_), .ZN(_01510__PTR7) );
  OR2_X1 U3230 ( .A1(_01506__PTR0), .A2(_02086__PTR1), .ZN(_01538__PTR0) );
  OR2_X1 U3231 ( .A1(_01530__PTR2), .A2(_01855__PTR0), .ZN(_01538__PTR1) );
  OR2_X1 U3232 ( .A1(_01537__PTR4), .A2(_01510__PTR6), .ZN(_01538__PTR2) );
  OR2_X1 U3233 ( .A1(_02417__PTR1), .A2(P3_P1_State2_PTR0), .ZN(_01310__PTR0) );
  OR2_X1 U3234 ( .A1(_01510__PTR7), .A2(_02050_), .ZN(_01526__PTR3) );
  OR2_X1 U3235 ( .A1(_01538__PTR0), .A2(_01538__PTR1), .ZN(_01539__PTR0) );
  OR2_X1 U3236 ( .A1(_01538__PTR2), .A2(_01526__PTR3), .ZN(_01539__PTR1) );
  OR2_X1 U3237 ( .A1(_01539__PTR0), .A2(_01539__PTR1), .ZN(_02098__PTR0) );
  OR2_X1 U3238 ( .A1(_02417__PTR2), .A2(P3_P1_State2_PTR0), .ZN(_01313__PTR0) );
  OR2_X1 U3239 ( .A1(_02098__PTR1), .A2(_02057_), .ZN(_01506__PTR1) );
  OR2_X1 U3240 ( .A1(_02056_), .A2(_02055_), .ZN(_01506__PTR2) );
  OR2_X1 U3241 ( .A1(_02054_), .A2(_01863__PTR0), .ZN(_01506__PTR3) );
  OR2_X1 U3242 ( .A1(_02090__PTR3), .A2(_01863__PTR2), .ZN(_01540__PTR4) );
  OR2_X1 U3243 ( .A1(_02090__PTR4), .A2(_02102__PTR2), .ZN(_01510__PTR4) );
  OR2_X1 U3244 ( .A1(_02098__PTR4), .A2(_02053_), .ZN(_01510__PTR5) );
  OR2_X1 U3245 ( .A1(_02417__PTR3), .A2(P3_P1_State2_PTR0), .ZN(_01316__PTR0) );
  OR2_X1 U3246 ( .A1(_01506__PTR0), .A2(_01506__PTR1), .ZN(_01507__PTR0) );
  OR2_X1 U3247 ( .A1(_01506__PTR2), .A2(_01506__PTR3), .ZN(_01507__PTR1) );
  OR2_X1 U3248 ( .A1(_01540__PTR4), .A2(_01510__PTR4), .ZN(_01541__PTR2) );
  OR2_X1 U3249 ( .A1(_01510__PTR5), .A2(_01540__PTR7), .ZN(_01541__PTR3) );
  OR2_X1 U3250 ( .A1(_02417__PTR4), .A2(P3_P1_State2_PTR0), .ZN(_01319__PTR0) );
  OR2_X1 U3251 ( .A1(_01507__PTR0), .A2(_01507__PTR1), .ZN(_01508__PTR0) );
  OR2_X1 U3252 ( .A1(_01541__PTR2), .A2(_01541__PTR3), .ZN(_01542__PTR1) );
  OR2_X1 U3253 ( .A1(_01508__PTR0), .A2(_01542__PTR1), .ZN(_01543_) );
  OR2_X1 U3254 ( .A1(_01543_), .A2(_02050_), .ZN(_02094__PTR0) );
  OR2_X1 U3255 ( .A1(_02417__PTR5), .A2(P3_P1_State2_PTR0), .ZN(_01322__PTR0) );
  OR2_X1 U3256 ( .A1(_02676__PTR1), .A2(_02633_), .ZN(_01544__PTR1) );
  OR2_X1 U3257 ( .A1(_02417__PTR6), .A2(P3_P1_State2_PTR0), .ZN(_01325__PTR0) );
  OR2_X1 U3258 ( .A1(_02632_), .A2(_02631_), .ZN(_01544__PTR2) );
  OR2_X1 U3259 ( .A1(_01544__PTR0), .A2(_01544__PTR1), .ZN(_01545__PTR0) );
  OR2_X1 U3260 ( .A1(_01544__PTR2), .A2(_01544__PTR3), .ZN(_01545__PTR1) );
  OR2_X1 U3261 ( .A1(_01545__PTR0), .A2(_01545__PTR1), .ZN(_01546_) );
  OR2_X1 U3262 ( .A1(_02417__PTR7), .A2(P3_P1_State2_PTR0), .ZN(_01328__PTR0) );
  OR2_X1 U3263 ( .A1(_01546_), .A2(_02628_), .ZN(_02664__PTR0) );
  OR2_X1 U3264 ( .A1(_02417__PTR8), .A2(P3_P1_State2_PTR0), .ZN(_01283__PTR0) );
  OR2_X1 U3265 ( .A1(_00292_), .A2(_02475__PTR32), .ZN(_01283__PTR1) );
  OR2_X1 U3266 ( .A1(_01283__PTR0), .A2(_01283__PTR1), .ZN(_00012_) );
  OR2_X1 U3267 ( .A1(P3_P1_State2_PTR0), .A2(_00292_), .ZN(_01284_) );
  OR2_X1 U3268 ( .A1(_01284_), .A2(_01766__PTR2), .ZN(_00013_) );
  OR2_X1 U3269 ( .A1(_00298_), .A2(P3_P1_State2_PTR1), .ZN(_01285__PTR0) );
  OR2_X1 U3270 ( .A1(_00299_), .A2(P3_P1_State2_PTR3), .ZN(_01281__PTR1) );
  OR2_X1 U3271 ( .A1(_01285__PTR0), .A2(_01281__PTR1), .ZN(_00014_) );
  OR2_X1 U3272 ( .A1(_00298_), .A2(_00293_), .ZN(_00151_) );
  OR2_X1 U3273 ( .A1(_00151_), .A2(_00037_), .ZN(_00015_) );
  OR2_X1 U3274 ( .A1(_00298_), .A2(_00292_), .ZN(_00016_) );
  OR2_X1 U3275 ( .A1(_00293_), .A2(_00299_), .ZN(_00009_) );
  OR2_X1 U3276 ( .A1(_00009_), .A2(P3_P1_State2_PTR3), .ZN(_00018_) );
  AND2_X1 U3277 ( .A1(_00012_), .A2(_00013_), .ZN(_01287__PTR0) );
  AND2_X1 U3278 ( .A1(_00014_), .A2(_00015_), .ZN(_01287__PTR1) );
  AND2_X1 U3279 ( .A1(_00016_), .A2(_00017_), .ZN(_01287__PTR2) );
  AND2_X1 U3280 ( .A1(_01287__PTR0), .A2(_01287__PTR1), .ZN(_01288__PTR0) );
  AND2_X1 U3281 ( .A1(_01287__PTR2), .A2(_00018_), .ZN(_01288__PTR1) );
  AND2_X1 U3282 ( .A1(_01288__PTR0), .A2(_01288__PTR1), .ZN(_00160_) );
  OR2_X1 U3283 ( .A1(_02417__PTR9), .A2(P3_P1_State2_PTR0), .ZN(_01289__PTR0) );
  OR2_X1 U3284 ( .A1(_01289__PTR0), .A2(_01283__PTR1), .ZN(_00019_) );
  AND2_X1 U3285 ( .A1(_00019_), .A2(_00013_), .ZN(_01290__PTR0) );
  AND2_X1 U3286 ( .A1(_01290__PTR0), .A2(_01287__PTR1), .ZN(_01291__PTR0) );
  AND2_X1 U3287 ( .A1(_01291__PTR0), .A2(_01288__PTR1), .ZN(_00161_) );
  OR2_X1 U3288 ( .A1(_02417__PTR10), .A2(P3_P1_State2_PTR0), .ZN(_01292__PTR0) );
  OR2_X1 U3289 ( .A1(_01292__PTR0), .A2(_01283__PTR1), .ZN(_00020_) );
  OR2_X1 U3290 ( .A1(_02148__PTR1), .A2(_02375__PTR4), .ZN(_01548__PTR2) );
  AND2_X1 U3291 ( .A1(_00020_), .A2(_00013_), .ZN(_01293__PTR0) );
  AND2_X1 U3292 ( .A1(_01293__PTR0), .A2(_01287__PTR1), .ZN(_01294__PTR0) );
  AND2_X1 U3293 ( .A1(_01294__PTR0), .A2(_01288__PTR1), .ZN(_00162_) );
  OR2_X1 U3294 ( .A1(_01548__PTR2), .A2(_01548__PTR3), .ZN(_01549__PTR1) );
  OR2_X1 U3295 ( .A1(_01549__PTR0), .A2(_01549__PTR1), .ZN(_01550_) );
  OR2_X1 U3296 ( .A1(_02417__PTR11), .A2(P3_P1_State2_PTR0), .ZN(_01295__PTR0) );
  OR2_X1 U3297 ( .A1(_01295__PTR0), .A2(_01283__PTR1), .ZN(_00021_) );
  AND2_X1 U3298 ( .A1(_00021_), .A2(_00013_), .ZN(_01296__PTR0) );
  AND2_X1 U3299 ( .A1(_01296__PTR0), .A2(_01287__PTR1), .ZN(_01297__PTR0) );
  AND2_X1 U3300 ( .A1(_01297__PTR0), .A2(_01288__PTR1), .ZN(_00163_) );
  OR2_X1 U3301 ( .A1(_01550_), .A2(_01547__PTR8), .ZN(_02409__PTR0) );
  OR2_X1 U3302 ( .A1(_02343_), .A2(_02379__PTR3), .ZN(_01551__PTR3) );
  OR2_X1 U3303 ( .A1(_02417__PTR12), .A2(P3_P1_State2_PTR0), .ZN(_01298__PTR0) );
  OR2_X1 U3304 ( .A1(_01298__PTR0), .A2(_01283__PTR1), .ZN(_00022_) );
  AND2_X1 U3305 ( .A1(_00022_), .A2(_00013_), .ZN(_01299__PTR0) );
  AND2_X1 U3306 ( .A1(_01299__PTR0), .A2(_01287__PTR1), .ZN(_01300__PTR0) );
  AND2_X1 U3307 ( .A1(_01300__PTR0), .A2(_01288__PTR1), .ZN(_00164_) );
  OR2_X1 U3308 ( .A1(_01547__PTR2), .A2(_01551__PTR3), .ZN(_01552__PTR1) );
  OR2_X1 U3309 ( .A1(_02417__PTR13), .A2(P3_P1_State2_PTR0), .ZN(_01301__PTR0) );
  OR2_X1 U3310 ( .A1(_01301__PTR0), .A2(_01283__PTR1), .ZN(_00023_) );
  OR2_X1 U3311 ( .A1(_01551__PTR4), .A2(_01551__PTR5), .ZN(_01552__PTR2) );
  AND2_X1 U3312 ( .A1(_00023_), .A2(_00013_), .ZN(_01302__PTR0) );
  AND2_X1 U3313 ( .A1(_01302__PTR0), .A2(_01287__PTR1), .ZN(_01303__PTR0) );
  AND2_X1 U3314 ( .A1(_01303__PTR0), .A2(_01288__PTR1), .ZN(_00165_) );
  OR2_X1 U3315 ( .A1(_01548__PTR0), .A2(_01552__PTR1), .ZN(_01553__PTR0) );
  OR2_X1 U3316 ( .A1(_01552__PTR2), .A2(_01552__PTR3), .ZN(_01553__PTR1) );
  OR2_X1 U3317 ( .A1(_01553__PTR0), .A2(_01553__PTR1), .ZN(_01554_) );
  OR2_X1 U3318 ( .A1(_02417__PTR14), .A2(P3_P1_State2_PTR0), .ZN(_01304__PTR0) );
  OR2_X1 U3319 ( .A1(_01304__PTR0), .A2(_01283__PTR1), .ZN(_00024_) );
  AND2_X1 U3320 ( .A1(_00024_), .A2(_00013_), .ZN(_01305__PTR0) );
  AND2_X1 U3321 ( .A1(_01305__PTR0), .A2(_01287__PTR1), .ZN(_01306__PTR0) );
  AND2_X1 U3322 ( .A1(_01306__PTR0), .A2(_01288__PTR1), .ZN(_00166_) );
  OR2_X1 U3323 ( .A1(_01554_), .A2(_02339_), .ZN(_02405__PTR0) );
  OR2_X1 U3324 ( .A1(_02417__PTR15), .A2(P3_P1_State2_PTR0), .ZN(_01307__PTR0) );
  OR2_X1 U3325 ( .A1(_01307__PTR0), .A2(_01283__PTR1), .ZN(_00025_) );
  OR2_X1 U3326 ( .A1(_02379__PTR3), .A2(_02391__PTR2), .ZN(_01555__PTR4) );
  AND2_X1 U3327 ( .A1(_00025_), .A2(_00013_), .ZN(_01308__PTR0) );
  AND2_X1 U3328 ( .A1(_01308__PTR0), .A2(_01287__PTR1), .ZN(_01309__PTR0) );
  AND2_X1 U3329 ( .A1(_01309__PTR0), .A2(_01288__PTR1), .ZN(_00167_) );
  OR2_X1 U3330 ( .A1(P3_P1_State2_PTR0), .A2(_00293_), .ZN(_01277__PTR0) );
  OR2_X1 U3331 ( .A1(_01277__PTR0), .A2(_01281__PTR1), .ZN(_00034_) );
  OR2_X1 U3332 ( .A1(_00034_), .A2(_02475__PTR14), .ZN(_00010_) );
  OR2_X1 U3333 ( .A1(_01555__PTR4), .A2(_01551__PTR5), .ZN(_01556__PTR2) );
  OR2_X1 U3334 ( .A1(_01556__PTR2), .A2(_01552__PTR3), .ZN(_01557__PTR1) );
  OR2_X1 U3335 ( .A1(_01549__PTR0), .A2(_01557__PTR1), .ZN(_01558_) );
  OR2_X1 U3336 ( .A1(_01558_), .A2(_02339_), .ZN(_02398__PTR0) );
  OR2_X1 U3337 ( .A1(_02343_), .A2(_02391__PTR2), .ZN(_01559__PTR3) );
  OR2_X1 U3338 ( .A1(_01547__PTR2), .A2(_01559__PTR3), .ZN(_01560__PTR1) );
  OR2_X1 U3339 ( .A1(_01551__PTR5), .A2(_01551__PTR6), .ZN(_01560__PTR2) );
  OR2_X1 U3340 ( .A1(_01548__PTR0), .A2(_01560__PTR1), .ZN(_01561__PTR0) );
  OR2_X1 U3341 ( .A1(_01560__PTR2), .A2(_01560__PTR3), .ZN(_01561__PTR1) );
  OR2_X1 U3342 ( .A1(_01561__PTR0), .A2(_01561__PTR1), .ZN(_02156__PTR3) );
  OR2_X1 U3343 ( .A1(_02347_), .A2(_02387__PTR1), .ZN(_01562__PTR0) );
  OR2_X1 U3344 ( .A1(_01562__PTR0), .A2(_02375__PTR1), .ZN(_01563__PTR0) );
  OR2_X1 U3345 ( .A1(_02163__PTR1), .A2(_01551__PTR5), .ZN(_01563__PTR2) );
  OR2_X1 U3346 ( .A1(_01551__PTR6), .A2(_01551__PTR7), .ZN(_01552__PTR3) );
  OR2_X1 U3347 ( .A1(_01563__PTR0), .A2(_01563__PTR1), .ZN(_01564__PTR0) );
  OR2_X1 U3348 ( .A1(_01563__PTR2), .A2(_01552__PTR3), .ZN(_01564__PTR1) );
  OR2_X1 U3349 ( .A1(_01564__PTR0), .A2(_01564__PTR1), .ZN(_01565_) );
  OR2_X1 U3350 ( .A1(_01565_), .A2(_02339_), .ZN(_02391__PTR0) );
  OR2_X1 U3351 ( .A1(_02156__PTR0), .A2(_02156__PTR2), .ZN(_02148__PTR0) );
  OR2_X1 U3352 ( .A1(_02391__PTR2), .A2(_02342_), .ZN(_01566__PTR4) );
  OR2_X1 U3353 ( .A1(_02341_), .A2(_02148__PTR2), .ZN(_01551__PTR6) );
  OR2_X1 U3354 ( .A1(_02148__PTR3), .A2(_02340_), .ZN(_01551__PTR7) );
  OR2_X1 U3355 ( .A1(_01517__PTR0), .A2(_02375__PTR1), .ZN(_01567__PTR0) );
  OR2_X1 U3356 ( .A1(_01562__PTR2), .A2(_02148__PTR0), .ZN(_01567__PTR1) );
  OR2_X1 U3357 ( .A1(_01566__PTR4), .A2(_01551__PTR6), .ZN(_01567__PTR2) );
  OR2_X1 U3358 ( .A1(_01551__PTR7), .A2(_02339_), .ZN(_01560__PTR3) );
  OR2_X1 U3359 ( .A1(_01567__PTR0), .A2(_01567__PTR1), .ZN(_01568__PTR0) );
  OR2_X1 U3360 ( .A1(_01567__PTR2), .A2(_01560__PTR3), .ZN(_01568__PTR1) );
  OR2_X1 U3361 ( .A1(_01568__PTR0), .A2(_01568__PTR1), .ZN(_02387__PTR0) );
  OR2_X1 U3362 ( .A1(_02347_), .A2(_02391__PTR1), .ZN(_01517__PTR0) );
  OR2_X1 U3363 ( .A1(_02387__PTR1), .A2(_02346_), .ZN(_01547__PTR1) );
  OR2_X1 U3364 ( .A1(_02345_), .A2(_02344_), .ZN(_01547__PTR2) );
  OR2_X1 U3365 ( .A1(_02343_), .A2(_02156__PTR0), .ZN(_01547__PTR3) );
  OR2_X1 U3366 ( .A1(_02379__PTR3), .A2(_02156__PTR2), .ZN(_01569__PTR4) );
  OR2_X1 U3367 ( .A1(_02379__PTR4), .A2(_02391__PTR2), .ZN(_01551__PTR4) );
  OR2_X1 U3368 ( .A1(_02387__PTR4), .A2(_02342_), .ZN(_01551__PTR5) );
  OR2_X1 U3369 ( .A1(_02341_), .A2(_02340_), .ZN(_01517__PTR3) );
  OR2_X1 U3370 ( .A1(_01517__PTR0), .A2(_01547__PTR1), .ZN(_01548__PTR0) );
  OR2_X1 U3371 ( .A1(_01547__PTR2), .A2(_01547__PTR3), .ZN(_01548__PTR1) );
  OR2_X1 U3372 ( .A1(_01569__PTR4), .A2(_01551__PTR4), .ZN(_01570__PTR2) );
  OR2_X1 U3373 ( .A1(_01551__PTR5), .A2(_01517__PTR3), .ZN(_01570__PTR3) );
  OR2_X1 U3374 ( .A1(_01548__PTR0), .A2(_01548__PTR1), .ZN(_01549__PTR0) );
  OR2_X1 U3375 ( .A1(_01570__PTR2), .A2(_01570__PTR3), .ZN(_01571__PTR1) );
  OR2_X1 U3376 ( .A1(_01549__PTR0), .A2(_01571__PTR1), .ZN(_01572_) );
  OR2_X1 U3377 ( .A1(_01572_), .A2(_02339_), .ZN(_02383__PTR0) );
  OR2_X1 U3378 ( .A1(P3_State_PTR0), .A2(_00288_), .ZN(_01274_) );
  OR2_X1 U3379 ( .A1(_01274_), .A2(P3_State_PTR2), .ZN(_00001_) );
  OR2_X1 U3380 ( .A1(P2_State_PTR0), .A2(_00286_), .ZN(_01346_) );
  OR2_X1 U3381 ( .A1(_01346_), .A2(P2_State_PTR2), .ZN(_00045_) );
  OR2_X1 U3382 ( .A1(P1_State_PTR0), .A2(_00276_), .ZN(_01418_) );
  OR2_X1 U3383 ( .A1(_01418_), .A2(P1_State_PTR2), .ZN(_00089_) );
  AND2_X1 U3384 ( .A1(_00306_), .A2(P3_State_PTR1), .ZN(_00256_) );
  AND2_X1 U3385 ( .A1(_00305_), .A2(P2_State_PTR1), .ZN(_00257_) );
  AND2_X1 U3386 ( .A1(_00311_), .A2(P1_State_PTR1), .ZN(_00258_) );
  OR2_X1 U3387 ( .A1(_02124__PTR1), .A2(_02124__PTR2), .ZN(_01573_) );
  OR2_X1 U3388 ( .A1(_01573_), .A2(_02124__PTR3), .ZN(_00135_) );
  OR2_X1 U3389 ( .A1(P1_DataWidth_PTR0), .A2(_01894__PTR9), .ZN(_01574__PTR0) );
  OR2_X1 U3390 ( .A1(_01574__PTR0), .A2(_01574__PTR1), .ZN(_01575__PTR0) );
  OR2_X1 U3391 ( .A1(_01575__PTR0), .A2(_01575__PTR1), .ZN(_01576__PTR0) );
  OR2_X1 U3392 ( .A1(_01576__PTR0), .A2(_01576__PTR1), .ZN(_01577__PTR0) );
  OR2_X1 U3393 ( .A1(_01577__PTR0), .A2(_01577__PTR1), .ZN(_01771_) );
  OR2_X1 U3394 ( .A1(_00289_), .A2(P1_StateBS16), .ZN(_01578__PTR0) );
  OR2_X1 U3395 ( .A1(_01578__PTR0), .A2(_01574__PTR1), .ZN(_01579__PTR0) );
  OR2_X1 U3396 ( .A1(_01579__PTR0), .A2(_01575__PTR1), .ZN(_01580__PTR0) );
  OR2_X1 U3397 ( .A1(_01580__PTR0), .A2(_01576__PTR1), .ZN(_01581__PTR0) );
  OR2_X1 U3398 ( .A1(_01581__PTR0), .A2(_01577__PTR1), .ZN(_01772_) );
  OR2_X1 U3399 ( .A1(_05760_), .A2(_05770_), .ZN(_00134_) );
  OR2_X1 U3400 ( .A1(_02102__PTR1), .A2(_02098__PTR1), .ZN(_01582__PTR0) );
  OR2_X1 U3401 ( .A1(_02057_), .A2(_02056_), .ZN(_02086__PTR1) );
  OR2_X1 U3402 ( .A1(_02055_), .A2(_02054_), .ZN(_01530__PTR2) );
  OR2_X1 U3403 ( .A1(_01863__PTR0), .A2(_02090__PTR3), .ZN(_01870__PTR0) );
  OR2_X1 U3404 ( .A1(_02102__PTR2), .A2(_02098__PTR4), .ZN(_02086__PTR4) );
  OR2_X1 U3405 ( .A1(_02053_), .A2(_02052_), .ZN(_01506__PTR6) );
  OR2_X1 U3406 ( .A1(_02051_), .A2(_02050_), .ZN(_01506__PTR8) );
  OR2_X1 U3407 ( .A1(_01582__PTR0), .A2(_02086__PTR1), .ZN(_01583__PTR0) );
  OR2_X1 U3408 ( .A1(_01530__PTR2), .A2(_01870__PTR0), .ZN(_01531__PTR1) );
  OR2_X1 U3409 ( .A1(_01870__PTR1), .A2(_02086__PTR4), .ZN(_01583__PTR2) );
  OR2_X1 U3410 ( .A1(_01506__PTR6), .A2(_02090__PTR6), .ZN(_01507__PTR3) );
  OR2_X1 U3411 ( .A1(_01583__PTR0), .A2(_01531__PTR1), .ZN(_01584__PTR0) );
  OR2_X1 U3412 ( .A1(_01583__PTR2), .A2(_01507__PTR3), .ZN(_01584__PTR1) );
  OR2_X1 U3413 ( .A1(_01584__PTR0), .A2(_01584__PTR1), .ZN(_01585_) );
  OR2_X1 U3414 ( .A1(_01585_), .A2(_01506__PTR8), .ZN(_01834_) );
  OR2_X1 U3415 ( .A1(_01586__PTR0), .A2(_01586__PTR1), .ZN(_01587__PTR0) );
  OR2_X1 U3416 ( .A1(_01587__PTR0), .A2(_01587__PTR1), .ZN(_01773_) );
  OR2_X1 U3417 ( .A1(_01586__PTR2), .A2(_01586__PTR3), .ZN(_01587__PTR1) );
  OR2_X1 U3418 ( .A1(_01589__PTR0), .A2(_01587__PTR1), .ZN(_01774_) );
  OR2_X1 U3419 ( .A1(_01586__PTR2), .A2(_01590__PTR3), .ZN(_01591__PTR1) );
  OR2_X1 U3420 ( .A1(_01589__PTR0), .A2(_01591__PTR1), .ZN(_01775_) );
  OR2_X1 U3421 ( .A1(_01592__PTR2), .A2(_01590__PTR3), .ZN(_01593__PTR1) );
  OR2_X1 U3422 ( .A1(_01589__PTR0), .A2(_01593__PTR1), .ZN(_01776_) );
  OR2_X1 U3423 ( .A1(_01594__PTR0), .A2(_01594__PTR1), .ZN(_01595__PTR0) );
  OR2_X1 U3424 ( .A1(_01595__PTR0), .A2(_01595__PTR1), .ZN(_01777_) );
  OR2_X1 U3425 ( .A1(_01883__PTR6), .A2(_01883__PTR7), .ZN(_01594__PTR3) );
  OR2_X1 U3426 ( .A1(_01586__PTR2), .A2(_01594__PTR3), .ZN(_01595__PTR1) );
  OR2_X1 U3427 ( .A1(_01596__PTR0), .A2(_01595__PTR1), .ZN(_01778_) );
  OR2_X1 U3428 ( .A1(_01598__PTR0), .A2(_01598__PTR1), .ZN(_01779_) );
  OR2_X1 U3429 ( .A1(_01588__PTR0), .A2(_01594__PTR1), .ZN(_01596__PTR0) );
  OR2_X1 U3430 ( .A1(_01596__PTR0), .A2(_01598__PTR1), .ZN(_01780_) );
  OR2_X1 U3431 ( .A1(_01600__PTR0), .A2(_01600__PTR1), .ZN(_01781_) );
  OR2_X1 U3432 ( .A1(_01883__PTR4), .A2(_01883__PTR5), .ZN(_01586__PTR2) );
  OR2_X1 U3433 ( .A1(_01586__PTR2), .A2(_01599__PTR3), .ZN(_01600__PTR1) );
  OR2_X1 U3434 ( .A1(_01601__PTR0), .A2(_01600__PTR1), .ZN(_01782_) );
  OR2_X1 U3435 ( .A1(_01601__PTR0), .A2(_01603__PTR1), .ZN(_01783_) );
  OR2_X1 U3436 ( .A1(_01588__PTR0), .A2(_01599__PTR1), .ZN(_01604__PTR0) );
  OR2_X1 U3437 ( .A1(_01604__PTR0), .A2(_01603__PTR1), .ZN(_01784_) );
  OR2_X1 U3438 ( .A1(_00269_), .A2(_00264_), .ZN(_01602__PTR2) );
  OR2_X1 U3439 ( .A1(_01602__PTR2), .A2(_01599__PTR3), .ZN(_01603__PTR1) );
  OR2_X1 U3440 ( .A1(_01589__PTR0), .A2(_01603__PTR1), .ZN(_01785_) );
  OR2_X1 U3441 ( .A1(_01597__PTR0), .A2(_01599__PTR1), .ZN(_01605__PTR0) );
  OR2_X1 U3442 ( .A1(_01605__PTR0), .A2(_01598__PTR1), .ZN(_01786_) );
  OR2_X1 U3443 ( .A1(_00267_), .A2(_01883__PTR1), .ZN(_01594__PTR0) );
  OR2_X1 U3444 ( .A1(_01594__PTR0), .A2(_01599__PTR1), .ZN(_01600__PTR0) );
  OR2_X1 U3445 ( .A1(_01600__PTR0), .A2(_01598__PTR1), .ZN(_01787_) );
  OR2_X1 U3446 ( .A1(_00267_), .A2(_00262_), .ZN(_01586__PTR0) );
  OR2_X1 U3447 ( .A1(_01883__PTR2), .A2(_00268_), .ZN(_01599__PTR1) );
  OR2_X1 U3448 ( .A1(_00265_), .A2(_00266_), .ZN(_01590__PTR3) );
  OR2_X1 U3449 ( .A1(_01586__PTR0), .A2(_01599__PTR1), .ZN(_01601__PTR0) );
  OR2_X1 U3450 ( .A1(_01597__PTR2), .A2(_01590__PTR3), .ZN(_01598__PTR1) );
  OR2_X1 U3451 ( .A1(_01601__PTR0), .A2(_01598__PTR1), .ZN(_01788_) );
  OR2_X1 U3452 ( .A1(_01883__PTR0), .A2(_00262_), .ZN(_01597__PTR0) );
  OR2_X1 U3453 ( .A1(_00263_), .A2(_01883__PTR3), .ZN(_01594__PTR1) );
  OR2_X1 U3454 ( .A1(_01883__PTR4), .A2(_00264_), .ZN(_01597__PTR2) );
  OR2_X1 U3455 ( .A1(_00265_), .A2(_01883__PTR7), .ZN(_01586__PTR3) );
  OR2_X1 U3456 ( .A1(_01597__PTR0), .A2(_01594__PTR1), .ZN(_01598__PTR0) );
  OR2_X1 U3457 ( .A1(_01597__PTR2), .A2(_01586__PTR3), .ZN(_01606__PTR1) );
  OR2_X1 U3458 ( .A1(_01598__PTR0), .A2(_01606__PTR1), .ZN(_01789_) );
  OR2_X1 U3459 ( .A1(_01883__PTR0), .A2(_01883__PTR1), .ZN(_01588__PTR0) );
  OR2_X1 U3460 ( .A1(_01883__PTR2), .A2(_01883__PTR3), .ZN(_01586__PTR1) );
  OR2_X1 U3461 ( .A1(_00269_), .A2(_01883__PTR5), .ZN(_01592__PTR2) );
  OR2_X1 U3462 ( .A1(_01883__PTR6), .A2(_00266_), .ZN(_01599__PTR3) );
  OR2_X1 U3463 ( .A1(_01588__PTR0), .A2(_01586__PTR1), .ZN(_01589__PTR0) );
  OR2_X1 U3464 ( .A1(_01592__PTR2), .A2(_01599__PTR3), .ZN(_01607__PTR1) );
  OR2_X1 U3465 ( .A1(_01589__PTR0), .A2(_01607__PTR1), .ZN(_01790_) );
  OR2_X1 U3466 ( .A1(P1_State_PTR0), .A2(P1_State_PTR1), .ZN(_01608_) );
  OR2_X1 U3467 ( .A1(_01608_), .A2(_00275_), .ZN(_01791_) );
  OR2_X1 U3468 ( .A1(P1_EAX_PTR0), .A2(P1_EAX_PTR1), .ZN(_01609__PTR0) );
  OR2_X1 U3469 ( .A1(P1_EAX_PTR2), .A2(P1_EAX_PTR3), .ZN(_01609__PTR1) );
  OR2_X1 U3470 ( .A1(P1_EAX_PTR4), .A2(P1_EAX_PTR5), .ZN(_01609__PTR2) );
  OR2_X1 U3471 ( .A1(P1_EAX_PTR6), .A2(P1_EAX_PTR7), .ZN(_01609__PTR3) );
  OR2_X1 U3472 ( .A1(P1_EAX_PTR8), .A2(P1_EAX_PTR9), .ZN(_01609__PTR4) );
  OR2_X1 U3473 ( .A1(P1_EAX_PTR10), .A2(P1_EAX_PTR11), .ZN(_01609__PTR5) );
  OR2_X1 U3474 ( .A1(P1_EAX_PTR12), .A2(P1_EAX_PTR13), .ZN(_01609__PTR6) );
  OR2_X1 U3475 ( .A1(P1_EAX_PTR14), .A2(P1_EAX_PTR15), .ZN(_01609__PTR7) );
  OR2_X1 U3476 ( .A1(_01609__PTR0), .A2(_01609__PTR1), .ZN(_01610__PTR0) );
  OR2_X1 U3477 ( .A1(_01609__PTR2), .A2(_01609__PTR3), .ZN(_01610__PTR1) );
  OR2_X1 U3478 ( .A1(_01609__PTR4), .A2(_01609__PTR5), .ZN(_01610__PTR2) );
  OR2_X1 U3479 ( .A1(_01609__PTR6), .A2(_01609__PTR7), .ZN(_01610__PTR3) );
  OR2_X1 U3480 ( .A1(_01610__PTR0), .A2(_01610__PTR1), .ZN(_01611__PTR0) );
  OR2_X1 U3481 ( .A1(_01610__PTR2), .A2(_01610__PTR3), .ZN(_01611__PTR1) );
  OR2_X1 U3482 ( .A1(_01611__PTR0), .A2(_01611__PTR1), .ZN(_02022_) );
  OR2_X1 U3483 ( .A1(di1_PTR16), .A2(di1_PTR17), .ZN(_01612__PTR8) );
  OR2_X1 U3484 ( .A1(di1_PTR18), .A2(di1_PTR19), .ZN(_01612__PTR9) );
  OR2_X1 U3485 ( .A1(di1_PTR20), .A2(di1_PTR21), .ZN(_01612__PTR10) );
  OR2_X1 U3486 ( .A1(di1_PTR22), .A2(di1_PTR23), .ZN(_01612__PTR11) );
  OR2_X1 U3487 ( .A1(_01612__PTR8), .A2(_01612__PTR9), .ZN(_01613__PTR4) );
  OR2_X1 U3488 ( .A1(_01612__PTR10), .A2(_01612__PTR11), .ZN(_01613__PTR5) );
  OR2_X1 U3489 ( .A1(_01613__PTR4), .A2(_01613__PTR5), .ZN(_01614__PTR2) );
  OR2_X1 U3490 ( .A1(_01614__PTR0), .A2(_01614__PTR1), .ZN(_01615_) );
  OR2_X1 U3491 ( .A1(_01615_), .A2(_01614__PTR2), .ZN(_01979_) );
  OR2_X1 U3492 ( .A1(di1_PTR0), .A2(di1_PTR1), .ZN(_01612__PTR0) );
  OR2_X1 U3493 ( .A1(di1_PTR2), .A2(di1_PTR3), .ZN(_01612__PTR1) );
  OR2_X1 U3494 ( .A1(di1_PTR4), .A2(di1_PTR5), .ZN(_01612__PTR2) );
  OR2_X1 U3495 ( .A1(di1_PTR6), .A2(di1_PTR7), .ZN(_01612__PTR3) );
  OR2_X1 U3496 ( .A1(di1_PTR8), .A2(di1_PTR9), .ZN(_01612__PTR4) );
  OR2_X1 U3497 ( .A1(di1_PTR10), .A2(di1_PTR11), .ZN(_01612__PTR5) );
  OR2_X1 U3498 ( .A1(di1_PTR12), .A2(di1_PTR13), .ZN(_01612__PTR6) );
  OR2_X1 U3499 ( .A1(di1_PTR14), .A2(di1_PTR15), .ZN(_01612__PTR7) );
  OR2_X1 U3500 ( .A1(_01612__PTR0), .A2(_01612__PTR1), .ZN(_01613__PTR0) );
  OR2_X1 U3501 ( .A1(_01612__PTR2), .A2(_01612__PTR3), .ZN(_01613__PTR1) );
  OR2_X1 U3502 ( .A1(_01612__PTR4), .A2(_01612__PTR5), .ZN(_01613__PTR2) );
  OR2_X1 U3503 ( .A1(_01612__PTR6), .A2(_01612__PTR7), .ZN(_01613__PTR3) );
  OR2_X1 U3504 ( .A1(_01613__PTR0), .A2(_01613__PTR1), .ZN(_01614__PTR0) );
  OR2_X1 U3505 ( .A1(_01613__PTR2), .A2(_01613__PTR3), .ZN(_01614__PTR1) );
  OR2_X1 U3506 ( .A1(_02668__PTR3), .A2(_02680__PTR2), .ZN(_01616__PTR4) );
  OR2_X1 U3507 ( .A1(_01616__PTR4), .A2(_01616__PTR5), .ZN(_01617__PTR2) );
  OR2_X1 U3508 ( .A1(_01617__PTR2), .A2(_01617__PTR3), .ZN(_01618__PTR1) );
  OR2_X1 U3509 ( .A1(_01618__PTR0), .A2(_01618__PTR1), .ZN(_01619_) );
  OR2_X1 U3510 ( .A1(_01619_), .A2(_02628_), .ZN(_02687__PTR0) );
  OR2_X1 U3511 ( .A1(_02437__PTR1), .A2(_02664__PTR4), .ZN(_01621__PTR2) );
  OR2_X1 U3512 ( .A1(_01621__PTR2), .A2(_01621__PTR3), .ZN(_01622__PTR1) );
  OR2_X1 U3513 ( .A1(_01618__PTR0), .A2(_01622__PTR1), .ZN(_01623_) );
  OR2_X1 U3514 ( .A1(_01623_), .A2(_01620__PTR8), .ZN(_02698__PTR0) );
  OR2_X1 U3515 ( .A1(_02632_), .A2(_02668__PTR3), .ZN(_01624__PTR3) );
  OR2_X1 U3516 ( .A1(_01616__PTR2), .A2(_01624__PTR3), .ZN(_01625__PTR1) );
  OR2_X1 U3517 ( .A1(_01624__PTR4), .A2(_01616__PTR5), .ZN(_01625__PTR2) );
  OR2_X1 U3518 ( .A1(_01617__PTR0), .A2(_01625__PTR1), .ZN(_01626__PTR0) );
  OR2_X1 U3519 ( .A1(_01625__PTR2), .A2(_01617__PTR3), .ZN(_01626__PTR1) );
  OR2_X1 U3520 ( .A1(_01626__PTR0), .A2(_01626__PTR1), .ZN(_01627_) );
  OR2_X1 U3521 ( .A1(_01627_), .A2(_02628_), .ZN(_02694__PTR0) );
  OR2_X1 U3522 ( .A1(P1_rEIP_PTR0), .A2(P1_rEIP_PTR1), .ZN(_01997_) );
  OR2_X1 U3523 ( .A1(_02413__PTR1), .A2(_02413__PTR2), .ZN(_01628_) );
  OR2_X1 U3524 ( .A1(_01628_), .A2(_02413__PTR3), .ZN(_00136_) );
  OR2_X1 U3525 ( .A1(P2_DataWidth_PTR0), .A2(_02186__PTR9), .ZN(_01629__PTR0) );
  OR2_X1 U3526 ( .A1(_01629__PTR0), .A2(_01629__PTR1), .ZN(_01630__PTR0) );
  OR2_X1 U3527 ( .A1(_01630__PTR0), .A2(_01630__PTR1), .ZN(_01631__PTR0) );
  OR2_X1 U3528 ( .A1(_01631__PTR0), .A2(_01631__PTR1), .ZN(_01632__PTR0) );
  OR2_X1 U3529 ( .A1(_01632__PTR0), .A2(_01632__PTR1), .ZN(_01792_) );
  OR2_X1 U3530 ( .A1(_00290_), .A2(P2_StateBS16), .ZN(_01633__PTR0) );
  OR2_X1 U3531 ( .A1(_01633__PTR0), .A2(_01629__PTR1), .ZN(_01634__PTR0) );
  OR2_X1 U3532 ( .A1(_01634__PTR0), .A2(_01630__PTR1), .ZN(_01635__PTR0) );
  OR2_X1 U3533 ( .A1(_01635__PTR0), .A2(_01631__PTR1), .ZN(_01636__PTR0) );
  OR2_X1 U3534 ( .A1(_01636__PTR0), .A2(_01632__PTR1), .ZN(_01793_) );
  OR2_X1 U3535 ( .A1(_02391__PTR1), .A2(_02387__PTR1), .ZN(_01637__PTR0) );
  OR2_X1 U3536 ( .A1(_02346_), .A2(_02345_), .ZN(_02375__PTR1) );
  OR2_X1 U3537 ( .A1(_02344_), .A2(_02343_), .ZN(_01562__PTR2) );
  OR2_X1 U3538 ( .A1(_02156__PTR0), .A2(_02379__PTR3), .ZN(_02163__PTR0) );
  OR2_X1 U3539 ( .A1(_02391__PTR2), .A2(_02387__PTR4), .ZN(_02375__PTR4) );
  OR2_X1 U3540 ( .A1(_02342_), .A2(_02341_), .ZN(_01547__PTR6) );
  OR2_X1 U3541 ( .A1(_02340_), .A2(_02339_), .ZN(_01547__PTR8) );
  OR2_X1 U3542 ( .A1(_01637__PTR0), .A2(_02375__PTR1), .ZN(_01638__PTR0) );
  OR2_X1 U3543 ( .A1(_01562__PTR2), .A2(_02163__PTR0), .ZN(_01563__PTR1) );
  OR2_X1 U3544 ( .A1(_02163__PTR1), .A2(_02375__PTR4), .ZN(_01638__PTR2) );
  OR2_X1 U3545 ( .A1(_01547__PTR6), .A2(_02379__PTR6), .ZN(_01548__PTR3) );
  OR2_X1 U3546 ( .A1(_01638__PTR0), .A2(_01563__PTR1), .ZN(_01639__PTR0) );
  OR2_X1 U3547 ( .A1(_01638__PTR2), .A2(_01548__PTR3), .ZN(_01639__PTR1) );
  OR2_X1 U3548 ( .A1(_01639__PTR0), .A2(_01639__PTR1), .ZN(_01640_) );
  OR2_X1 U3549 ( .A1(_01640_), .A2(_01547__PTR8), .ZN(_02127_) );
  OR2_X1 U3550 ( .A1(_01641__PTR0), .A2(_01641__PTR1), .ZN(_01642__PTR0) );
  OR2_X1 U3551 ( .A1(_01642__PTR0), .A2(_01642__PTR1), .ZN(_01794_) );
  OR2_X1 U3552 ( .A1(_01641__PTR2), .A2(_01641__PTR3), .ZN(_01642__PTR1) );
  OR2_X1 U3553 ( .A1(_01644__PTR0), .A2(_01642__PTR1), .ZN(_01795_) );
  OR2_X1 U3554 ( .A1(_01641__PTR2), .A2(_01645__PTR3), .ZN(_01646__PTR1) );
  OR2_X1 U3555 ( .A1(_01644__PTR0), .A2(_01646__PTR1), .ZN(_01796_) );
  OR2_X1 U3556 ( .A1(_01647__PTR2), .A2(_01645__PTR3), .ZN(_01648__PTR1) );
  OR2_X1 U3557 ( .A1(_01644__PTR0), .A2(_01648__PTR1), .ZN(_01797_) );
  OR2_X1 U3558 ( .A1(_01649__PTR0), .A2(_01649__PTR1), .ZN(_01650__PTR0) );
  OR2_X1 U3559 ( .A1(_01650__PTR0), .A2(_01650__PTR1), .ZN(_01798_) );
  OR2_X1 U3560 ( .A1(_02175__PTR6), .A2(_02175__PTR7), .ZN(_01649__PTR3) );
  OR2_X1 U3561 ( .A1(_01641__PTR2), .A2(_01649__PTR3), .ZN(_01650__PTR1) );
  OR2_X1 U3562 ( .A1(_01651__PTR0), .A2(_01650__PTR1), .ZN(_01799_) );
  OR2_X1 U3563 ( .A1(_01653__PTR0), .A2(_01653__PTR1), .ZN(_01800_) );
  OR2_X1 U3564 ( .A1(_01643__PTR0), .A2(_01649__PTR1), .ZN(_01651__PTR0) );
  OR2_X1 U3565 ( .A1(_01651__PTR0), .A2(_01653__PTR1), .ZN(_01801_) );
  OR2_X1 U3566 ( .A1(_01655__PTR0), .A2(_01655__PTR1), .ZN(_01802_) );
  OR2_X1 U3567 ( .A1(_02175__PTR4), .A2(_02175__PTR5), .ZN(_01641__PTR2) );
  OR2_X1 U3568 ( .A1(_01641__PTR2), .A2(_01654__PTR3), .ZN(_01655__PTR1) );
  OR2_X1 U3569 ( .A1(_01656__PTR0), .A2(_01655__PTR1), .ZN(_01803_) );
  OR2_X1 U3570 ( .A1(_01656__PTR0), .A2(_01658__PTR1), .ZN(_01804_) );
  OR2_X1 U3571 ( .A1(_01643__PTR0), .A2(_01654__PTR1), .ZN(_01659__PTR0) );
  OR2_X1 U3572 ( .A1(_01659__PTR0), .A2(_01658__PTR1), .ZN(_01805_) );
  OR2_X1 U3573 ( .A1(_00261_), .A2(_00272_), .ZN(_01657__PTR2) );
  OR2_X1 U3574 ( .A1(_01657__PTR2), .A2(_01654__PTR3), .ZN(_01658__PTR1) );
  OR2_X1 U3575 ( .A1(_01644__PTR0), .A2(_01658__PTR1), .ZN(_01806_) );
  OR2_X1 U3576 ( .A1(_01652__PTR0), .A2(_01654__PTR1), .ZN(_01660__PTR0) );
  OR2_X1 U3577 ( .A1(_01660__PTR0), .A2(_01653__PTR1), .ZN(_01807_) );
  OR2_X1 U3578 ( .A1(_00274_), .A2(_02175__PTR1), .ZN(_01649__PTR0) );
  OR2_X1 U3579 ( .A1(_01649__PTR0), .A2(_01654__PTR1), .ZN(_01655__PTR0) );
  OR2_X1 U3580 ( .A1(_01655__PTR0), .A2(_01653__PTR1), .ZN(_01808_) );
  OR2_X1 U3581 ( .A1(_00274_), .A2(_00270_), .ZN(_01641__PTR0) );
  OR2_X1 U3582 ( .A1(_02175__PTR2), .A2(_00271_), .ZN(_01654__PTR1) );
  OR2_X1 U3583 ( .A1(_00259_), .A2(_00260_), .ZN(_01645__PTR3) );
  OR2_X1 U3584 ( .A1(_01641__PTR0), .A2(_01654__PTR1), .ZN(_01656__PTR0) );
  OR2_X1 U3585 ( .A1(_01652__PTR2), .A2(_01645__PTR3), .ZN(_01653__PTR1) );
  OR2_X1 U3586 ( .A1(_01656__PTR0), .A2(_01653__PTR1), .ZN(_01809_) );
  OR2_X1 U3587 ( .A1(_02175__PTR0), .A2(_00270_), .ZN(_01652__PTR0) );
  OR2_X1 U3588 ( .A1(_00273_), .A2(_02175__PTR3), .ZN(_01649__PTR1) );
  OR2_X1 U3589 ( .A1(_02175__PTR4), .A2(_00272_), .ZN(_01652__PTR2) );
  OR2_X1 U3590 ( .A1(_00259_), .A2(_02175__PTR7), .ZN(_01641__PTR3) );
  OR2_X1 U3591 ( .A1(_01652__PTR0), .A2(_01649__PTR1), .ZN(_01653__PTR0) );
  OR2_X1 U3592 ( .A1(_01652__PTR2), .A2(_01641__PTR3), .ZN(_01661__PTR1) );
  OR2_X1 U3593 ( .A1(_01653__PTR0), .A2(_01661__PTR1), .ZN(_01810_) );
  OR2_X1 U3594 ( .A1(_02175__PTR0), .A2(_02175__PTR1), .ZN(_01643__PTR0) );
  OR2_X1 U3595 ( .A1(_02175__PTR2), .A2(_02175__PTR3), .ZN(_01641__PTR1) );
  OR2_X1 U3596 ( .A1(_00261_), .A2(_02175__PTR5), .ZN(_01647__PTR2) );
  OR2_X1 U3597 ( .A1(_02175__PTR6), .A2(_00260_), .ZN(_01654__PTR3) );
  OR2_X1 U3598 ( .A1(_01643__PTR0), .A2(_01641__PTR1), .ZN(_01644__PTR0) );
  OR2_X1 U3599 ( .A1(_01647__PTR2), .A2(_01654__PTR3), .ZN(_01662__PTR1) );
  OR2_X1 U3600 ( .A1(_01644__PTR0), .A2(_01662__PTR1), .ZN(_01811_) );
  OR2_X1 U3601 ( .A1(P2_State_PTR0), .A2(P2_State_PTR1), .ZN(_01663_) );
  OR2_X1 U3602 ( .A1(_01663_), .A2(_00285_), .ZN(_01812_) );
  OR2_X1 U3603 ( .A1(P2_EAX_PTR0), .A2(P2_EAX_PTR1), .ZN(_01664__PTR0) );
  OR2_X1 U3604 ( .A1(P2_EAX_PTR2), .A2(P2_EAX_PTR3), .ZN(_01664__PTR1) );
  OR2_X1 U3605 ( .A1(P2_EAX_PTR4), .A2(P2_EAX_PTR5), .ZN(_01664__PTR2) );
  OR2_X1 U3606 ( .A1(P2_EAX_PTR6), .A2(P2_EAX_PTR7), .ZN(_01664__PTR3) );
  OR2_X1 U3607 ( .A1(P2_EAX_PTR8), .A2(P2_EAX_PTR9), .ZN(_01664__PTR4) );
  OR2_X1 U3608 ( .A1(P2_EAX_PTR10), .A2(P2_EAX_PTR11), .ZN(_01664__PTR5) );
  OR2_X1 U3609 ( .A1(P2_EAX_PTR12), .A2(P2_EAX_PTR13), .ZN(_01664__PTR6) );
  OR2_X1 U3610 ( .A1(P2_EAX_PTR14), .A2(P2_EAX_PTR15), .ZN(_01664__PTR7) );
  OR2_X1 U3611 ( .A1(_01664__PTR0), .A2(_01664__PTR1), .ZN(_01665__PTR0) );
  OR2_X1 U3612 ( .A1(_01664__PTR2), .A2(_01664__PTR3), .ZN(_01665__PTR1) );
  OR2_X1 U3613 ( .A1(_01664__PTR4), .A2(_01664__PTR5), .ZN(_01665__PTR2) );
  OR2_X1 U3614 ( .A1(_01664__PTR6), .A2(_01664__PTR7), .ZN(_01665__PTR3) );
  OR2_X1 U3615 ( .A1(_01665__PTR0), .A2(_01665__PTR1), .ZN(_01666__PTR0) );
  OR2_X1 U3616 ( .A1(_01665__PTR2), .A2(_01665__PTR3), .ZN(_01666__PTR1) );
  OR2_X1 U3617 ( .A1(_01666__PTR0), .A2(_01666__PTR1), .ZN(_02312_) );
  OR2_X1 U3618 ( .A1(di2_PTR16), .A2(di2_PTR17), .ZN(_01667__PTR8) );
  OR2_X1 U3619 ( .A1(di2_PTR18), .A2(di2_PTR19), .ZN(_01667__PTR9) );
  OR2_X1 U3620 ( .A1(di2_PTR20), .A2(di2_PTR21), .ZN(_01667__PTR10) );
  OR2_X1 U3621 ( .A1(di2_PTR22), .A2(di2_PTR23), .ZN(_01667__PTR11) );
  OR2_X1 U3622 ( .A1(_01667__PTR8), .A2(_01667__PTR9), .ZN(_01668__PTR4) );
  OR2_X1 U3623 ( .A1(_01667__PTR10), .A2(_01667__PTR11), .ZN(_01668__PTR5) );
  OR2_X1 U3624 ( .A1(_01668__PTR4), .A2(_01668__PTR5), .ZN(_01669__PTR2) );
  OR2_X1 U3625 ( .A1(_01669__PTR0), .A2(_01669__PTR1), .ZN(_01670_) );
  OR2_X1 U3626 ( .A1(_01670_), .A2(_01669__PTR2), .ZN(_02271_) );
  OR2_X1 U3627 ( .A1(di2_PTR0), .A2(di2_PTR1), .ZN(_01667__PTR0) );
  OR2_X1 U3628 ( .A1(di2_PTR2), .A2(di2_PTR3), .ZN(_01667__PTR1) );
  OR2_X1 U3629 ( .A1(di2_PTR4), .A2(di2_PTR5), .ZN(_01667__PTR2) );
  OR2_X1 U3630 ( .A1(di2_PTR6), .A2(di2_PTR7), .ZN(_01667__PTR3) );
  OR2_X1 U3631 ( .A1(di2_PTR8), .A2(di2_PTR9), .ZN(_01667__PTR4) );
  OR2_X1 U3632 ( .A1(di2_PTR10), .A2(di2_PTR11), .ZN(_01667__PTR5) );
  OR2_X1 U3633 ( .A1(di2_PTR12), .A2(di2_PTR13), .ZN(_01667__PTR6) );
  OR2_X1 U3634 ( .A1(di2_PTR14), .A2(di2_PTR15), .ZN(_01667__PTR7) );
  OR2_X1 U3635 ( .A1(_01667__PTR0), .A2(_01667__PTR1), .ZN(_01668__PTR0) );
  OR2_X1 U3636 ( .A1(_01667__PTR2), .A2(_01667__PTR3), .ZN(_01668__PTR1) );
  OR2_X1 U3637 ( .A1(_01667__PTR4), .A2(_01667__PTR5), .ZN(_01668__PTR2) );
  OR2_X1 U3638 ( .A1(_01667__PTR6), .A2(_01667__PTR7), .ZN(_01668__PTR3) );
  OR2_X1 U3639 ( .A1(_01668__PTR0), .A2(_01668__PTR1), .ZN(_01669__PTR0) );
  OR2_X1 U3640 ( .A1(_01668__PTR2), .A2(_01668__PTR3), .ZN(_01669__PTR1) );
  OR2_X1 U3641 ( .A1(P2_rEIP_PTR0), .A2(P2_rEIP_PTR1), .ZN(_02289_) );
  OR2_X1 U3642 ( .A1(_02702__PTR1), .A2(_02702__PTR2), .ZN(_01671_) );
  OR2_X1 U3643 ( .A1(_01671_), .A2(_02702__PTR3), .ZN(_00137_) );
  OR2_X1 U3644 ( .A1(P3_DataWidth_PTR0), .A2(_02475__PTR9), .ZN(_01672__PTR0) );
  OR2_X1 U3645 ( .A1(_01672__PTR0), .A2(_01672__PTR1), .ZN(_01673__PTR0) );
  OR2_X1 U3646 ( .A1(_01673__PTR0), .A2(_01673__PTR1), .ZN(_01674__PTR0) );
  OR2_X1 U3647 ( .A1(_01674__PTR0), .A2(_01674__PTR1), .ZN(_01675__PTR0) );
  OR2_X1 U3648 ( .A1(_01675__PTR0), .A2(_01675__PTR1), .ZN(_01813_) );
  OR2_X1 U3649 ( .A1(_00291_), .A2(P3_StateBS16), .ZN(_01676__PTR0) );
  OR2_X1 U3650 ( .A1(_01676__PTR0), .A2(_01672__PTR1), .ZN(_01677__PTR0) );
  OR2_X1 U3651 ( .A1(_01677__PTR0), .A2(_01673__PTR1), .ZN(_01678__PTR0) );
  OR2_X1 U3652 ( .A1(_01678__PTR0), .A2(_01674__PTR1), .ZN(_01679__PTR0) );
  OR2_X1 U3653 ( .A1(_01679__PTR0), .A2(_01675__PTR1), .ZN(_01814_) );
  OR2_X1 U3654 ( .A1(_02632_), .A2(_02680__PTR2), .ZN(_01680__PTR3) );
  OR2_X1 U3655 ( .A1(_01616__PTR2), .A2(_01680__PTR3), .ZN(_01681__PTR1) );
  OR2_X1 U3656 ( .A1(_01616__PTR5), .A2(_01616__PTR6), .ZN(_01681__PTR2) );
  OR2_X1 U3657 ( .A1(_01617__PTR0), .A2(_01681__PTR1), .ZN(_01682__PTR0) );
  OR2_X1 U3658 ( .A1(_01681__PTR2), .A2(_01681__PTR3), .ZN(_01682__PTR1) );
  OR2_X1 U3659 ( .A1(_01682__PTR0), .A2(_01682__PTR1), .ZN(_02445__PTR3) );
  OR2_X1 U3660 ( .A1(_02636_), .A2(_02676__PTR1), .ZN(_01683__PTR0) );
  OR2_X1 U3661 ( .A1(_01683__PTR0), .A2(_02664__PTR1), .ZN(_01684__PTR0) );
  OR2_X1 U3662 ( .A1(_02452__PTR1), .A2(_01616__PTR5), .ZN(_01684__PTR2) );
  OR2_X1 U3663 ( .A1(_01616__PTR6), .A2(_01616__PTR7), .ZN(_01617__PTR3) );
  OR2_X1 U3664 ( .A1(_01684__PTR0), .A2(_01684__PTR1), .ZN(_01685__PTR0) );
  OR2_X1 U3665 ( .A1(_01684__PTR2), .A2(_01617__PTR3), .ZN(_01685__PTR1) );
  OR2_X1 U3666 ( .A1(_01685__PTR0), .A2(_01685__PTR1), .ZN(_01686_) );
  OR2_X1 U3667 ( .A1(_01686_), .A2(_02628_), .ZN(_02680__PTR0) );
  OR2_X1 U3668 ( .A1(_02680__PTR1), .A2(_02676__PTR1), .ZN(_01687__PTR0) );
  OR2_X1 U3669 ( .A1(_02445__PTR0), .A2(_02668__PTR3), .ZN(_02452__PTR0) );
  OR2_X1 U3670 ( .A1(_02631_), .A2(_02630_), .ZN(_01620__PTR6) );
  OR2_X1 U3671 ( .A1(_02629_), .A2(_02628_), .ZN(_01620__PTR8) );
  OR2_X1 U3672 ( .A1(_01687__PTR0), .A2(_02664__PTR1), .ZN(_01688__PTR0) );
  OR2_X1 U3673 ( .A1(_01683__PTR2), .A2(_02452__PTR0), .ZN(_01684__PTR1) );
  OR2_X1 U3674 ( .A1(_02452__PTR1), .A2(_02664__PTR4), .ZN(_01688__PTR2) );
  OR2_X1 U3675 ( .A1(_01620__PTR6), .A2(_02668__PTR6), .ZN(_01621__PTR3) );
  OR2_X1 U3676 ( .A1(_01688__PTR0), .A2(_01684__PTR1), .ZN(_01689__PTR0) );
  OR2_X1 U3677 ( .A1(_01688__PTR2), .A2(_01621__PTR3), .ZN(_01689__PTR1) );
  OR2_X1 U3678 ( .A1(_01689__PTR0), .A2(_01689__PTR1), .ZN(_01690_) );
  OR2_X1 U3679 ( .A1(_01690_), .A2(_01620__PTR8), .ZN(_02416_) );
  OR2_X1 U3680 ( .A1(_01691__PTR0), .A2(_01691__PTR1), .ZN(_01692__PTR0) );
  OR2_X1 U3681 ( .A1(_01692__PTR0), .A2(_01692__PTR1), .ZN(_01815_) );
  OR2_X1 U3682 ( .A1(_01691__PTR2), .A2(_01691__PTR3), .ZN(_01692__PTR1) );
  OR2_X1 U3683 ( .A1(_01694__PTR0), .A2(_01692__PTR1), .ZN(_01816_) );
  OR2_X1 U3684 ( .A1(_01691__PTR2), .A2(_01695__PTR3), .ZN(_01696__PTR1) );
  OR2_X1 U3685 ( .A1(_01694__PTR0), .A2(_01696__PTR1), .ZN(_01817_) );
  OR2_X1 U3686 ( .A1(_01697__PTR2), .A2(_01695__PTR3), .ZN(_01698__PTR1) );
  OR2_X1 U3687 ( .A1(_01694__PTR0), .A2(_01698__PTR1), .ZN(_01818_) );
  OR2_X1 U3688 ( .A1(_01699__PTR0), .A2(_01699__PTR1), .ZN(_01700__PTR0) );
  OR2_X1 U3689 ( .A1(_01700__PTR0), .A2(_01700__PTR1), .ZN(_01819_) );
  OR2_X1 U3690 ( .A1(_02464__PTR6), .A2(_02464__PTR7), .ZN(_01699__PTR3) );
  OR2_X1 U3691 ( .A1(_01691__PTR2), .A2(_01699__PTR3), .ZN(_01700__PTR1) );
  OR2_X1 U3692 ( .A1(_01701__PTR0), .A2(_01700__PTR1), .ZN(_01820_) );
  OR2_X1 U3693 ( .A1(_01703__PTR0), .A2(_01703__PTR1), .ZN(_01821_) );
  OR2_X1 U3694 ( .A1(_01693__PTR0), .A2(_01699__PTR1), .ZN(_01701__PTR0) );
  OR2_X1 U3695 ( .A1(_01701__PTR0), .A2(_01703__PTR1), .ZN(_01822_) );
  OR2_X1 U3696 ( .A1(_01705__PTR0), .A2(_01705__PTR1), .ZN(_01823_) );
  OR2_X1 U3697 ( .A1(_02464__PTR4), .A2(_02464__PTR5), .ZN(_01691__PTR2) );
  OR2_X1 U3698 ( .A1(_01691__PTR2), .A2(_01704__PTR3), .ZN(_01705__PTR1) );
  OR2_X1 U3699 ( .A1(_01706__PTR0), .A2(_01705__PTR1), .ZN(_01824_) );
  OR2_X1 U3700 ( .A1(_01706__PTR0), .A2(_01708__PTR1), .ZN(_01825_) );
  OR2_X1 U3701 ( .A1(_01693__PTR0), .A2(_01704__PTR1), .ZN(_01709__PTR0) );
  OR2_X1 U3702 ( .A1(_01709__PTR0), .A2(_01708__PTR1), .ZN(_01826_) );
  OR2_X1 U3703 ( .A1(_00281_), .A2(_00279_), .ZN(_01707__PTR2) );
  OR2_X1 U3704 ( .A1(_01707__PTR2), .A2(_01704__PTR3), .ZN(_01708__PTR1) );
  OR2_X1 U3705 ( .A1(_01694__PTR0), .A2(_01708__PTR1), .ZN(_01827_) );
  OR2_X1 U3706 ( .A1(_01702__PTR0), .A2(_01704__PTR1), .ZN(_01710__PTR0) );
  OR2_X1 U3707 ( .A1(_01710__PTR0), .A2(_01703__PTR1), .ZN(_01828_) );
  OR2_X1 U3708 ( .A1(_00283_), .A2(_02464__PTR1), .ZN(_01699__PTR0) );
  OR2_X1 U3709 ( .A1(_01699__PTR0), .A2(_01704__PTR1), .ZN(_01705__PTR0) );
  OR2_X1 U3710 ( .A1(_01705__PTR0), .A2(_01703__PTR1), .ZN(_01829_) );
  OR2_X1 U3711 ( .A1(_00283_), .A2(_00277_), .ZN(_01691__PTR0) );
  OR2_X1 U3712 ( .A1(_02464__PTR2), .A2(_00284_), .ZN(_01704__PTR1) );
  OR2_X1 U3713 ( .A1(_00280_), .A2(_00282_), .ZN(_01695__PTR3) );
  OR2_X1 U3714 ( .A1(_01691__PTR0), .A2(_01704__PTR1), .ZN(_01706__PTR0) );
  OR2_X1 U3715 ( .A1(_01702__PTR2), .A2(_01695__PTR3), .ZN(_01703__PTR1) );
  OR2_X1 U3716 ( .A1(_01706__PTR0), .A2(_01703__PTR1), .ZN(_01830_) );
  OR2_X1 U3717 ( .A1(_02464__PTR0), .A2(_00277_), .ZN(_01702__PTR0) );
  OR2_X1 U3718 ( .A1(_00278_), .A2(_02464__PTR3), .ZN(_01699__PTR1) );
  OR2_X1 U3719 ( .A1(_02464__PTR4), .A2(_00279_), .ZN(_01702__PTR2) );
  OR2_X1 U3720 ( .A1(_00280_), .A2(_02464__PTR7), .ZN(_01691__PTR3) );
  OR2_X1 U3721 ( .A1(_01702__PTR0), .A2(_01699__PTR1), .ZN(_01703__PTR0) );
  OR2_X1 U3722 ( .A1(_01702__PTR2), .A2(_01691__PTR3), .ZN(_01711__PTR1) );
  OR2_X1 U3723 ( .A1(_01703__PTR0), .A2(_01711__PTR1), .ZN(_01831_) );
  OR2_X1 U3724 ( .A1(_02464__PTR0), .A2(_02464__PTR1), .ZN(_01693__PTR0) );
  OR2_X1 U3725 ( .A1(_02464__PTR2), .A2(_02464__PTR3), .ZN(_01691__PTR1) );
  OR2_X1 U3726 ( .A1(_00281_), .A2(_02464__PTR5), .ZN(_01697__PTR2) );
  OR2_X1 U3727 ( .A1(_02464__PTR6), .A2(_00282_), .ZN(_01704__PTR3) );
  OR2_X1 U3728 ( .A1(_01693__PTR0), .A2(_01691__PTR1), .ZN(_01694__PTR0) );
  OR2_X1 U3729 ( .A1(_01697__PTR2), .A2(_01704__PTR3), .ZN(_01712__PTR1) );
  OR2_X1 U3730 ( .A1(_01694__PTR0), .A2(_01712__PTR1), .ZN(_01832_) );
  OR2_X1 U3731 ( .A1(P3_State_PTR0), .A2(P3_State_PTR1), .ZN(_01713_) );
  OR2_X1 U3732 ( .A1(_01713_), .A2(_00287_), .ZN(_01833_) );
  OR2_X1 U3733 ( .A1(P3_EAX_PTR0), .A2(P3_EAX_PTR1), .ZN(_01714__PTR0) );
  OR2_X1 U3734 ( .A1(P3_EAX_PTR2), .A2(P3_EAX_PTR3), .ZN(_01714__PTR1) );
  OR2_X1 U3735 ( .A1(P3_EAX_PTR4), .A2(P3_EAX_PTR5), .ZN(_01714__PTR2) );
  OR2_X1 U3736 ( .A1(P3_EAX_PTR6), .A2(P3_EAX_PTR7), .ZN(_01714__PTR3) );
  OR2_X1 U3737 ( .A1(P3_EAX_PTR8), .A2(P3_EAX_PTR9), .ZN(_01714__PTR4) );
  OR2_X1 U3738 ( .A1(P3_EAX_PTR10), .A2(P3_EAX_PTR11), .ZN(_01714__PTR5) );
  OR2_X1 U3739 ( .A1(P3_EAX_PTR12), .A2(P3_EAX_PTR13), .ZN(_01714__PTR6) );
  OR2_X1 U3740 ( .A1(P3_EAX_PTR14), .A2(P3_EAX_PTR15), .ZN(_01714__PTR7) );
  OR2_X1 U3741 ( .A1(_01714__PTR0), .A2(_01714__PTR1), .ZN(_01715__PTR0) );
  OR2_X1 U3742 ( .A1(_01714__PTR2), .A2(_01714__PTR3), .ZN(_01715__PTR1) );
  OR2_X1 U3743 ( .A1(_01714__PTR4), .A2(_01714__PTR5), .ZN(_01715__PTR2) );
  OR2_X1 U3744 ( .A1(_01714__PTR6), .A2(_01714__PTR7), .ZN(_01715__PTR3) );
  OR2_X1 U3745 ( .A1(_01715__PTR0), .A2(_01715__PTR1), .ZN(_01716__PTR0) );
  OR2_X1 U3746 ( .A1(_01715__PTR2), .A2(_01715__PTR3), .ZN(_01716__PTR1) );
  OR2_X1 U3747 ( .A1(_01716__PTR0), .A2(_01716__PTR1), .ZN(_02601_) );
  OR2_X1 U3748 ( .A1(_02058_), .A2(_02102__PTR1), .ZN(_01506__PTR0) );
  OR2_X1 U3749 ( .A1(_02098__PTR1), .A2(_02055_), .ZN(_01717__PTR1) );
  OR2_X1 U3750 ( .A1(_02054_), .A2(_02053_), .ZN(_01717__PTR2) );
  OR2_X1 U3751 ( .A1(_02052_), .A2(_02051_), .ZN(_01540__PTR7) );
  OR2_X1 U3752 ( .A1(_01506__PTR0), .A2(_01717__PTR1), .ZN(_01718__PTR0) );
  OR2_X1 U3753 ( .A1(_01717__PTR2), .A2(_01540__PTR7), .ZN(_01718__PTR1) );
  OR2_X1 U3754 ( .A1(_01718__PTR0), .A2(_01718__PTR1), .ZN(_01719_) );
  OR2_X1 U3755 ( .A1(_01719_), .A2(_02050_), .ZN(_02086__PTR0) );
  OR2_X1 U3756 ( .A1(buf2_PTR16), .A2(buf2_PTR17), .ZN(_01720__PTR8) );
  OR2_X1 U3757 ( .A1(buf2_PTR18), .A2(buf2_PTR19), .ZN(_01720__PTR9) );
  OR2_X1 U3758 ( .A1(buf2_PTR20), .A2(buf2_PTR21), .ZN(_01720__PTR10) );
  OR2_X1 U3759 ( .A1(buf2_PTR22), .A2(buf2_PTR23), .ZN(_01720__PTR11) );
  OR2_X1 U3760 ( .A1(_01720__PTR8), .A2(_01720__PTR9), .ZN(_01721__PTR4) );
  OR2_X1 U3761 ( .A1(_01720__PTR10), .A2(_01720__PTR11), .ZN(_01721__PTR5) );
  OR2_X1 U3762 ( .A1(_01721__PTR4), .A2(_01721__PTR5), .ZN(_01722__PTR2) );
  OR2_X1 U3763 ( .A1(_01722__PTR0), .A2(_01722__PTR1), .ZN(_01723_) );
  OR2_X1 U3764 ( .A1(_01723_), .A2(_01722__PTR2), .ZN(_02560_) );
  OR2_X1 U3765 ( .A1(buf2_PTR0), .A2(buf2_PTR1), .ZN(_01720__PTR0) );
  OR2_X1 U3766 ( .A1(buf2_PTR2), .A2(buf2_PTR3), .ZN(_01720__PTR1) );
  OR2_X1 U3767 ( .A1(buf2_PTR4), .A2(buf2_PTR5), .ZN(_01720__PTR2) );
  OR2_X1 U3768 ( .A1(buf2_PTR6), .A2(buf2_PTR7), .ZN(_01720__PTR3) );
  OR2_X1 U3769 ( .A1(buf2_PTR8), .A2(buf2_PTR9), .ZN(_01720__PTR4) );
  OR2_X1 U3770 ( .A1(buf2_PTR10), .A2(buf2_PTR11), .ZN(_01720__PTR5) );
  OR2_X1 U3771 ( .A1(buf2_PTR12), .A2(buf2_PTR13), .ZN(_01720__PTR6) );
  OR2_X1 U3772 ( .A1(buf2_PTR14), .A2(buf2_PTR15), .ZN(_01720__PTR7) );
  OR2_X1 U3773 ( .A1(_01720__PTR0), .A2(_01720__PTR1), .ZN(_01721__PTR0) );
  OR2_X1 U3774 ( .A1(_01720__PTR2), .A2(_01720__PTR3), .ZN(_01721__PTR1) );
  OR2_X1 U3775 ( .A1(_01720__PTR4), .A2(_01720__PTR5), .ZN(_01721__PTR2) );
  OR2_X1 U3776 ( .A1(_01720__PTR6), .A2(_01720__PTR7), .ZN(_01721__PTR3) );
  OR2_X1 U3777 ( .A1(_01721__PTR0), .A2(_01721__PTR1), .ZN(_01722__PTR0) );
  OR2_X1 U3778 ( .A1(_01721__PTR2), .A2(_01721__PTR3), .ZN(_01722__PTR1) );
  OR2_X1 U3779 ( .A1(_02635_), .A2(_02634_), .ZN(_02664__PTR1) );
  OR2_X1 U3780 ( .A1(_02633_), .A2(_02632_), .ZN(_01683__PTR2) );
  OR2_X1 U3781 ( .A1(_02445__PTR0), .A2(_02445__PTR2), .ZN(_02437__PTR0) );
  OR2_X1 U3782 ( .A1(_02680__PTR2), .A2(_02631_), .ZN(_01724__PTR4) );
  OR2_X1 U3783 ( .A1(_02630_), .A2(_02437__PTR2), .ZN(_01616__PTR6) );
  OR2_X1 U3784 ( .A1(_02437__PTR3), .A2(_02629_), .ZN(_01616__PTR7) );
  OR2_X1 U3785 ( .A1(_01544__PTR0), .A2(_02664__PTR1), .ZN(_01725__PTR0) );
  OR2_X1 U3786 ( .A1(_01683__PTR2), .A2(_02437__PTR0), .ZN(_01725__PTR1) );
  OR2_X1 U3787 ( .A1(_01724__PTR4), .A2(_01616__PTR6), .ZN(_01725__PTR2) );
  OR2_X1 U3788 ( .A1(_01616__PTR7), .A2(_02628_), .ZN(_01681__PTR3) );
  OR2_X1 U3789 ( .A1(_01725__PTR0), .A2(_01725__PTR1), .ZN(_01726__PTR0) );
  OR2_X1 U3790 ( .A1(_01725__PTR2), .A2(_01681__PTR3), .ZN(_01726__PTR1) );
  OR2_X1 U3791 ( .A1(_01726__PTR0), .A2(_01726__PTR1), .ZN(_02676__PTR0) );
  OR2_X1 U3792 ( .A1(_02636_), .A2(_02680__PTR1), .ZN(_01544__PTR0) );
  OR2_X1 U3793 ( .A1(_02676__PTR1), .A2(_02635_), .ZN(_01616__PTR1) );
  OR2_X1 U3794 ( .A1(_02634_), .A2(_02633_), .ZN(_01616__PTR2) );
  OR2_X1 U3795 ( .A1(_02632_), .A2(_02445__PTR0), .ZN(_01616__PTR3) );
  OR2_X1 U3796 ( .A1(_02668__PTR3), .A2(_02445__PTR2), .ZN(_01727__PTR4) );
  OR2_X1 U3797 ( .A1(_02668__PTR4), .A2(_02680__PTR2), .ZN(_01624__PTR4) );
  OR2_X1 U3798 ( .A1(_02676__PTR4), .A2(_02631_), .ZN(_01616__PTR5) );
  OR2_X1 U3799 ( .A1(_02630_), .A2(_02629_), .ZN(_01544__PTR3) );
  OR2_X1 U3800 ( .A1(_01544__PTR0), .A2(_01616__PTR1), .ZN(_01617__PTR0) );
  OR2_X1 U3801 ( .A1(_01616__PTR2), .A2(_01616__PTR3), .ZN(_01617__PTR1) );
  OR2_X1 U3802 ( .A1(_01727__PTR4), .A2(_01624__PTR4), .ZN(_01728__PTR2) );
  OR2_X1 U3803 ( .A1(_01616__PTR5), .A2(_01544__PTR3), .ZN(_01728__PTR3) );
  OR2_X1 U3804 ( .A1(_01617__PTR0), .A2(_01617__PTR1), .ZN(_01618__PTR0) );
  OR2_X1 U3805 ( .A1(_01728__PTR2), .A2(_01728__PTR3), .ZN(_01729__PTR1) );
  OR2_X1 U3806 ( .A1(_01618__PTR0), .A2(_01729__PTR1), .ZN(_01730_) );
  OR2_X1 U3807 ( .A1(_01730_), .A2(_02628_), .ZN(_02672__PTR0) );
  OR2_X1 U3808 ( .A1(_02680__PTR2), .A2(_02676__PTR4), .ZN(_02664__PTR4) );
  OR2_X1 U3809 ( .A1(P3_rEIP_PTR0), .A2(P3_rEIP_PTR1), .ZN(_02578_) );
  OR2_X1 U3810 ( .A1(_02123__PTR11), .A2(_02123__PTR15), .ZN(_02126__PTR3) );
  OR2_X1 U3811 ( .A1(_02123__PTR10), .A2(_02123__PTR14), .ZN(_01731__PTR1) );
  OR2_X1 U3812 ( .A1(_02123__PTR6), .A2(_01731__PTR1), .ZN(_02126__PTR2) );
  OR2_X1 U3813 ( .A1(_02123__PTR9), .A2(_02123__PTR13), .ZN(_01732__PTR1) );
  OR2_X1 U3814 ( .A1(_02123__PTR5), .A2(_01732__PTR1), .ZN(_02126__PTR1) );
  OR2_X1 U3815 ( .A1(_02123__PTR8), .A2(_02123__PTR12), .ZN(_01733__PTR1) );
  OR2_X1 U3816 ( .A1(_02123__PTR4), .A2(_01733__PTR1), .ZN(_02126__PTR0) );
  OR2_X1 U3817 ( .A1(_02124__PTR0), .A2(_02124__PTR1), .ZN(_01734__PTR0) );
  OR2_X1 U3818 ( .A1(_02124__PTR2), .A2(_02124__PTR3), .ZN(_01734__PTR1) );
  OR2_X1 U3819 ( .A1(_01734__PTR0), .A2(_01734__PTR1), .ZN(_02929_) );
  OR2_X1 U3820 ( .A1(_02115__PTR31), .A2(_02115__PTR63), .ZN(_01735_) );
  OR2_X1 U3821 ( .A1(_01735_), .A2(_02115__PTR95), .ZN(_02117__PTR31) );
  OR2_X1 U3822 ( .A1(_02115__PTR30), .A2(_02115__PTR62), .ZN(_01736_) );
  OR2_X1 U3823 ( .A1(_01736_), .A2(_02115__PTR94), .ZN(_02117__PTR30) );
  OR2_X1 U3824 ( .A1(_02115__PTR29), .A2(_02115__PTR61), .ZN(_01737_) );
  OR2_X1 U3825 ( .A1(_01737_), .A2(_02115__PTR93), .ZN(_02117__PTR29) );
  OR2_X1 U3826 ( .A1(_02115__PTR28), .A2(_02115__PTR60), .ZN(_01738_) );
  OR2_X1 U3827 ( .A1(_01738_), .A2(_02115__PTR92), .ZN(_02117__PTR28) );
  OR2_X1 U3828 ( .A1(_02115__PTR27), .A2(_02115__PTR59), .ZN(_01739_) );
  OR2_X1 U3829 ( .A1(_01739_), .A2(_02115__PTR91), .ZN(_02117__PTR27) );
  OR2_X1 U3830 ( .A1(_02115__PTR26), .A2(_02115__PTR58), .ZN(_01740_) );
  OR2_X1 U3831 ( .A1(_01740_), .A2(_02115__PTR90), .ZN(_02117__PTR26) );
  OR2_X1 U3832 ( .A1(_02115__PTR25), .A2(_02115__PTR57), .ZN(_01741_) );
  OR2_X1 U3833 ( .A1(_01741_), .A2(_02115__PTR89), .ZN(_02117__PTR25) );
  OR2_X1 U3834 ( .A1(_02115__PTR24), .A2(_02115__PTR56), .ZN(_01742_) );
  OR2_X1 U3835 ( .A1(_01742_), .A2(_02115__PTR88), .ZN(_02117__PTR24) );
  OR2_X1 U3836 ( .A1(P1_BE_n_PTR0), .A2(P1_BE_n_PTR1), .ZN(_01744__PTR0) );
  OR2_X1 U3837 ( .A1(P1_BE_n_PTR2), .A2(P1_BE_n_PTR3), .ZN(_01744__PTR1) );
  OR2_X1 U3838 ( .A1(_01744__PTR0), .A2(_01744__PTR1), .ZN(_01745_) );
  OR2_X1 U3839 ( .A1(P2_BE_n_PTR0), .A2(P2_BE_n_PTR1), .ZN(_01746__PTR0) );
  OR2_X1 U3840 ( .A1(P2_BE_n_PTR2), .A2(P2_BE_n_PTR3), .ZN(_01746__PTR1) );
  OR2_X1 U3841 ( .A1(_01746__PTR0), .A2(_01746__PTR1), .ZN(_01747_) );
  OR2_X1 U3842 ( .A1(P3_BE_n_PTR0), .A2(P3_BE_n_PTR1), .ZN(_01748__PTR0) );
  OR2_X1 U3843 ( .A1(P3_BE_n_PTR2), .A2(P3_BE_n_PTR3), .ZN(_01748__PTR1) );
  OR2_X1 U3844 ( .A1(_01748__PTR0), .A2(_01748__PTR1), .ZN(_01749_) );
  OR2_X1 U3845 ( .A1(P1_DataWidth_PTR0), .A2(P1_StateBS16), .ZN(_01750__PTR0) );
  OR2_X1 U3846 ( .A1(P1_DataWidth_PTR2), .A2(P1_DataWidth_PTR3), .ZN(_01574__PTR1) );
  OR2_X1 U3847 ( .A1(P1_DataWidth_PTR4), .A2(P1_DataWidth_PTR5), .ZN(_01574__PTR2) );
  OR2_X1 U3848 ( .A1(P1_DataWidth_PTR6), .A2(P1_DataWidth_PTR7), .ZN(_01574__PTR3) );
  OR2_X1 U3849 ( .A1(P1_DataWidth_PTR8), .A2(P1_DataWidth_PTR9), .ZN(_01574__PTR4) );
  OR2_X1 U3850 ( .A1(P1_DataWidth_PTR10), .A2(P1_DataWidth_PTR11), .ZN(_01574__PTR5) );
  OR2_X1 U3851 ( .A1(P1_DataWidth_PTR12), .A2(P1_DataWidth_PTR13), .ZN(_01574__PTR6) );
  OR2_X1 U3852 ( .A1(P1_DataWidth_PTR14), .A2(P1_DataWidth_PTR15), .ZN(_01574__PTR7) );
  OR2_X1 U3853 ( .A1(P1_DataWidth_PTR16), .A2(P1_DataWidth_PTR17), .ZN(_01574__PTR8) );
  OR2_X1 U3854 ( .A1(P1_DataWidth_PTR18), .A2(P1_DataWidth_PTR19), .ZN(_01574__PTR9) );
  OR2_X1 U3855 ( .A1(P1_DataWidth_PTR20), .A2(P1_DataWidth_PTR21), .ZN(_01574__PTR10) );
  OR2_X1 U3856 ( .A1(P1_DataWidth_PTR22), .A2(P1_DataWidth_PTR23), .ZN(_01574__PTR11) );
  OR2_X1 U3857 ( .A1(P1_DataWidth_PTR24), .A2(P1_DataWidth_PTR25), .ZN(_01574__PTR12) );
  OR2_X1 U3858 ( .A1(P1_DataWidth_PTR26), .A2(P1_DataWidth_PTR27), .ZN(_01574__PTR13) );
  OR2_X1 U3859 ( .A1(P1_DataWidth_PTR28), .A2(P1_DataWidth_PTR29), .ZN(_01574__PTR14) );
  OR2_X1 U3860 ( .A1(P1_DataWidth_PTR30), .A2(P1_DataWidth_PTR31), .ZN(_01574__PTR15) );
  OR2_X1 U3861 ( .A1(_01750__PTR0), .A2(_01574__PTR1), .ZN(_01751__PTR0) );
  OR2_X1 U3862 ( .A1(_01574__PTR2), .A2(_01574__PTR3), .ZN(_01575__PTR1) );
  OR2_X1 U3863 ( .A1(_01574__PTR4), .A2(_01574__PTR5), .ZN(_01575__PTR2) );
  OR2_X1 U3864 ( .A1(_01574__PTR6), .A2(_01574__PTR7), .ZN(_01575__PTR3) );
  OR2_X1 U3865 ( .A1(_01574__PTR8), .A2(_01574__PTR9), .ZN(_01575__PTR4) );
  OR2_X1 U3866 ( .A1(_01574__PTR10), .A2(_01574__PTR11), .ZN(_01575__PTR5) );
  OR2_X1 U3867 ( .A1(_01574__PTR12), .A2(_01574__PTR13), .ZN(_01575__PTR6) );
  OR2_X1 U3868 ( .A1(_01574__PTR14), .A2(_01574__PTR15), .ZN(_01575__PTR7) );
  OR2_X1 U3869 ( .A1(_01751__PTR0), .A2(_01575__PTR1), .ZN(_01752__PTR0) );
  OR2_X1 U3870 ( .A1(_01575__PTR2), .A2(_01575__PTR3), .ZN(_01576__PTR1) );
  OR2_X1 U3871 ( .A1(_01575__PTR4), .A2(_01575__PTR5), .ZN(_01576__PTR2) );
  OR2_X1 U3872 ( .A1(_01575__PTR6), .A2(_01575__PTR7), .ZN(_01576__PTR3) );
  OR2_X1 U3873 ( .A1(_01752__PTR0), .A2(_01576__PTR1), .ZN(_01753__PTR0) );
  OR2_X1 U3874 ( .A1(_01576__PTR2), .A2(_01576__PTR3), .ZN(_01577__PTR1) );
  OR2_X1 U3875 ( .A1(_01753__PTR0), .A2(_01577__PTR1), .ZN(_01754_) );
  OR2_X1 U3876 ( .A1(P2_DataWidth_PTR0), .A2(P2_StateBS16), .ZN(_01755__PTR0) );
  OR2_X1 U3877 ( .A1(P2_DataWidth_PTR2), .A2(P2_DataWidth_PTR3), .ZN(_01629__PTR1) );
  OR2_X1 U3878 ( .A1(P2_DataWidth_PTR4), .A2(P2_DataWidth_PTR5), .ZN(_01629__PTR2) );
  OR2_X1 U3879 ( .A1(P2_DataWidth_PTR6), .A2(P2_DataWidth_PTR7), .ZN(_01629__PTR3) );
  OR2_X1 U3880 ( .A1(P2_DataWidth_PTR8), .A2(P2_DataWidth_PTR9), .ZN(_01629__PTR4) );
  OR2_X1 U3881 ( .A1(P2_DataWidth_PTR10), .A2(P2_DataWidth_PTR11), .ZN(_01629__PTR5) );
  OR2_X1 U3882 ( .A1(P2_DataWidth_PTR12), .A2(P2_DataWidth_PTR13), .ZN(_01629__PTR6) );
  OR2_X1 U3883 ( .A1(P2_DataWidth_PTR14), .A2(P2_DataWidth_PTR15), .ZN(_01629__PTR7) );
  OR2_X1 U3884 ( .A1(P2_DataWidth_PTR16), .A2(P2_DataWidth_PTR17), .ZN(_01629__PTR8) );
  OR2_X1 U3885 ( .A1(P2_DataWidth_PTR18), .A2(P2_DataWidth_PTR19), .ZN(_01629__PTR9) );
  OR2_X1 U3886 ( .A1(P2_DataWidth_PTR20), .A2(P2_DataWidth_PTR21), .ZN(_01629__PTR10) );
  OR2_X1 U3887 ( .A1(P2_DataWidth_PTR22), .A2(P2_DataWidth_PTR23), .ZN(_01629__PTR11) );
  OR2_X1 U3888 ( .A1(P2_DataWidth_PTR24), .A2(P2_DataWidth_PTR25), .ZN(_01629__PTR12) );
  OR2_X1 U3889 ( .A1(P2_DataWidth_PTR26), .A2(P2_DataWidth_PTR27), .ZN(_01629__PTR13) );
  OR2_X1 U3890 ( .A1(P2_DataWidth_PTR28), .A2(P2_DataWidth_PTR29), .ZN(_01629__PTR14) );
  OR2_X1 U3891 ( .A1(P2_DataWidth_PTR30), .A2(P2_DataWidth_PTR31), .ZN(_01629__PTR15) );
  OR2_X1 U3892 ( .A1(_01755__PTR0), .A2(_01629__PTR1), .ZN(_01756__PTR0) );
  OR2_X1 U3893 ( .A1(_01629__PTR2), .A2(_01629__PTR3), .ZN(_01630__PTR1) );
  OR2_X1 U3894 ( .A1(_01629__PTR4), .A2(_01629__PTR5), .ZN(_01630__PTR2) );
  OR2_X1 U3895 ( .A1(_01629__PTR6), .A2(_01629__PTR7), .ZN(_01630__PTR3) );
  OR2_X1 U3896 ( .A1(_01629__PTR8), .A2(_01629__PTR9), .ZN(_01630__PTR4) );
  OR2_X1 U3897 ( .A1(_01629__PTR10), .A2(_01629__PTR11), .ZN(_01630__PTR5) );
  OR2_X1 U3898 ( .A1(_01629__PTR12), .A2(_01629__PTR13), .ZN(_01630__PTR6) );
  OR2_X1 U3899 ( .A1(_01629__PTR14), .A2(_01629__PTR15), .ZN(_01630__PTR7) );
  OR2_X1 U3900 ( .A1(_01756__PTR0), .A2(_01630__PTR1), .ZN(_01757__PTR0) );
  OR2_X1 U3901 ( .A1(_01630__PTR2), .A2(_01630__PTR3), .ZN(_01631__PTR1) );
  OR2_X1 U3902 ( .A1(_01630__PTR4), .A2(_01630__PTR5), .ZN(_01631__PTR2) );
  OR2_X1 U3903 ( .A1(_01630__PTR6), .A2(_01630__PTR7), .ZN(_01631__PTR3) );
  OR2_X1 U3904 ( .A1(_01757__PTR0), .A2(_01631__PTR1), .ZN(_01758__PTR0) );
  OR2_X1 U3905 ( .A1(_01631__PTR2), .A2(_01631__PTR3), .ZN(_01632__PTR1) );
  OR2_X1 U3906 ( .A1(_01758__PTR0), .A2(_01632__PTR1), .ZN(_01759_) );
  OR2_X1 U3907 ( .A1(P3_DataWidth_PTR0), .A2(P3_StateBS16), .ZN(_01760__PTR0) );
  OR2_X1 U3908 ( .A1(P3_DataWidth_PTR2), .A2(P3_DataWidth_PTR3), .ZN(_01672__PTR1) );
  OR2_X1 U3909 ( .A1(P3_DataWidth_PTR4), .A2(P3_DataWidth_PTR5), .ZN(_01672__PTR2) );
  OR2_X1 U3910 ( .A1(P3_DataWidth_PTR6), .A2(P3_DataWidth_PTR7), .ZN(_01672__PTR3) );
  OR2_X1 U3911 ( .A1(P3_DataWidth_PTR8), .A2(P3_DataWidth_PTR9), .ZN(_01672__PTR4) );
  OR2_X1 U3912 ( .A1(P3_DataWidth_PTR10), .A2(P3_DataWidth_PTR11), .ZN(_01672__PTR5) );
  OR2_X1 U3913 ( .A1(P3_DataWidth_PTR12), .A2(P3_DataWidth_PTR13), .ZN(_01672__PTR6) );
  OR2_X1 U3914 ( .A1(P3_DataWidth_PTR14), .A2(P3_DataWidth_PTR15), .ZN(_01672__PTR7) );
  OR2_X1 U3915 ( .A1(P3_DataWidth_PTR16), .A2(P3_DataWidth_PTR17), .ZN(_01672__PTR8) );
  OR2_X1 U3916 ( .A1(P3_DataWidth_PTR18), .A2(P3_DataWidth_PTR19), .ZN(_01672__PTR9) );
  OR2_X1 U3917 ( .A1(P3_DataWidth_PTR20), .A2(P3_DataWidth_PTR21), .ZN(_01672__PTR10) );
  OR2_X1 U3918 ( .A1(P3_DataWidth_PTR22), .A2(P3_DataWidth_PTR23), .ZN(_01672__PTR11) );
  OR2_X1 U3919 ( .A1(P3_DataWidth_PTR24), .A2(P3_DataWidth_PTR25), .ZN(_01672__PTR12) );
  OR2_X1 U3920 ( .A1(P3_DataWidth_PTR26), .A2(P3_DataWidth_PTR27), .ZN(_01672__PTR13) );
  OR2_X1 U3921 ( .A1(P3_DataWidth_PTR28), .A2(P3_DataWidth_PTR29), .ZN(_01672__PTR14) );
  OR2_X1 U3922 ( .A1(P3_DataWidth_PTR30), .A2(P3_DataWidth_PTR31), .ZN(_01672__PTR15) );
  OR2_X1 U3923 ( .A1(_01760__PTR0), .A2(_01672__PTR1), .ZN(_01761__PTR0) );
  OR2_X1 U3924 ( .A1(_01672__PTR2), .A2(_01672__PTR3), .ZN(_01673__PTR1) );
  OR2_X1 U3925 ( .A1(_01672__PTR4), .A2(_01672__PTR5), .ZN(_01673__PTR2) );
  OR2_X1 U3926 ( .A1(_01672__PTR6), .A2(_01672__PTR7), .ZN(_01673__PTR3) );
  OR2_X1 U3927 ( .A1(_01672__PTR8), .A2(_01672__PTR9), .ZN(_01673__PTR4) );
  OR2_X1 U3928 ( .A1(_01672__PTR10), .A2(_01672__PTR11), .ZN(_01673__PTR5) );
  OR2_X1 U3929 ( .A1(_01672__PTR12), .A2(_01672__PTR13), .ZN(_01673__PTR6) );
  OR2_X1 U3930 ( .A1(_01672__PTR14), .A2(_01672__PTR15), .ZN(_01673__PTR7) );
  OR2_X1 U3931 ( .A1(_01761__PTR0), .A2(_01673__PTR1), .ZN(_01762__PTR0) );
  OR2_X1 U3932 ( .A1(_01673__PTR2), .A2(_01673__PTR3), .ZN(_01674__PTR1) );
  OR2_X1 U3933 ( .A1(_01673__PTR4), .A2(_01673__PTR5), .ZN(_01674__PTR2) );
  OR2_X1 U3934 ( .A1(_01673__PTR6), .A2(_01673__PTR7), .ZN(_01674__PTR3) );
  OR2_X1 U3935 ( .A1(_01762__PTR0), .A2(_01674__PTR1), .ZN(_01763__PTR0) );
  OR2_X1 U3936 ( .A1(_01674__PTR2), .A2(_01674__PTR3), .ZN(_01675__PTR1) );
  OR2_X1 U3937 ( .A1(_01763__PTR0), .A2(_01675__PTR1), .ZN(_01764_) );
  INV_X1 U3938 ( .A(_01745_), .ZN(_05755_) );
  INV_X1 U3939 ( .A(_01747_), .ZN(_05765_) );
  INV_X1 U3940 ( .A(_01749_), .ZN(_05745_) );
  INV_X1 U3941 ( .A(_01771_), .ZN(_02124__PTR1) );
  INV_X1 U3942 ( .A(_01772_), .ZN(_02124__PTR2) );
  INV_X1 U3943 ( .A(_01754_), .ZN(_02124__PTR3) );
  INV_X1 U3944 ( .A(_01773_), .ZN(_02102__PTR1) );
  INV_X1 U3945 ( .A(_01774_), .ZN(_02098__PTR1) );
  INV_X1 U3946 ( .A(_01775_), .ZN(_02057_) );
  INV_X1 U3947 ( .A(_01776_), .ZN(_02056_) );
  INV_X1 U3948 ( .A(_01777_), .ZN(_02055_) );
  INV_X1 U3949 ( .A(_01778_), .ZN(_02054_) );
  INV_X1 U3950 ( .A(_01779_), .ZN(_01863__PTR0) );
  INV_X1 U3951 ( .A(_01780_), .ZN(_02090__PTR3) );
  INV_X1 U3952 ( .A(_01781_), .ZN(_01863__PTR2) );
  INV_X1 U3953 ( .A(_01782_), .ZN(_02090__PTR4) );
  INV_X1 U3954 ( .A(_01783_), .ZN(_02102__PTR2) );
  INV_X1 U3955 ( .A(_01784_), .ZN(_02098__PTR4) );
  INV_X1 U3956 ( .A(_01785_), .ZN(_02053_) );
  INV_X1 U3957 ( .A(_01786_), .ZN(_02052_) );
  INV_X1 U3958 ( .A(_01787_), .ZN(_01855__PTR2) );
  INV_X1 U3959 ( .A(_01788_), .ZN(_01855__PTR3) );
  INV_X1 U3960 ( .A(_01789_), .ZN(_02051_) );
  INV_X1 U3961 ( .A(_01790_), .ZN(_02050_) );
  INV_X1 U3962 ( .A(_01791_), .ZN(_02024_) );
  INV_X1 U3963 ( .A(_00089_), .ZN(_02023_) );
  INV_X1 U3964 ( .A(_01792_), .ZN(_02413__PTR1) );
  INV_X1 U3965 ( .A(_01793_), .ZN(_02413__PTR2) );
  INV_X1 U3966 ( .A(_01759_), .ZN(_02413__PTR3) );
  INV_X1 U3967 ( .A(_01794_), .ZN(_02391__PTR1) );
  INV_X1 U3968 ( .A(_01795_), .ZN(_02387__PTR1) );
  INV_X1 U3969 ( .A(_01796_), .ZN(_02346_) );
  INV_X1 U3970 ( .A(_01797_), .ZN(_02345_) );
  INV_X1 U3971 ( .A(_01798_), .ZN(_02344_) );
  INV_X1 U3972 ( .A(_01799_), .ZN(_02343_) );
  INV_X1 U3973 ( .A(_01800_), .ZN(_02156__PTR0) );
  INV_X1 U3974 ( .A(_01801_), .ZN(_02379__PTR3) );
  INV_X1 U3975 ( .A(_01802_), .ZN(_02156__PTR2) );
  INV_X1 U3976 ( .A(_01803_), .ZN(_02379__PTR4) );
  INV_X1 U3977 ( .A(_01804_), .ZN(_02391__PTR2) );
  INV_X1 U3978 ( .A(_01805_), .ZN(_02387__PTR4) );
  INV_X1 U3979 ( .A(_01806_), .ZN(_02342_) );
  INV_X1 U3980 ( .A(_01807_), .ZN(_02341_) );
  INV_X1 U3981 ( .A(_01808_), .ZN(_02148__PTR2) );
  INV_X1 U3982 ( .A(_01809_), .ZN(_02148__PTR3) );
  INV_X1 U3983 ( .A(_01810_), .ZN(_02340_) );
  INV_X1 U3984 ( .A(_01811_), .ZN(_02339_) );
  INV_X1 U3985 ( .A(_01812_), .ZN(_02314_) );
  INV_X1 U3986 ( .A(_00045_), .ZN(_02313_) );
  INV_X1 U3987 ( .A(_01813_), .ZN(_02702__PTR1) );
  INV_X1 U3988 ( .A(_01814_), .ZN(_02702__PTR2) );
  INV_X1 U3989 ( .A(_01764_), .ZN(_02702__PTR3) );
  INV_X1 U3990 ( .A(_01815_), .ZN(_02680__PTR1) );
  INV_X1 U3991 ( .A(_01816_), .ZN(_02676__PTR1) );
  INV_X1 U3992 ( .A(_01817_), .ZN(_02635_) );
  INV_X1 U3993 ( .A(_01818_), .ZN(_02634_) );
  INV_X1 U3994 ( .A(_01819_), .ZN(_02633_) );
  INV_X1 U3995 ( .A(_01820_), .ZN(_02632_) );
  INV_X1 U3996 ( .A(_01821_), .ZN(_02445__PTR0) );
  INV_X1 U3997 ( .A(_01822_), .ZN(_02668__PTR3) );
  INV_X1 U3998 ( .A(_01823_), .ZN(_02445__PTR2) );
  INV_X1 U3999 ( .A(_01824_), .ZN(_02668__PTR4) );
  INV_X1 U4000 ( .A(_01825_), .ZN(_02680__PTR2) );
  INV_X1 U4001 ( .A(_01826_), .ZN(_02676__PTR4) );
  INV_X1 U4002 ( .A(_01827_), .ZN(_02631_) );
  INV_X1 U4003 ( .A(_01828_), .ZN(_02630_) );
  INV_X1 U4004 ( .A(_01829_), .ZN(_02437__PTR2) );
  INV_X1 U4005 ( .A(_01830_), .ZN(_02437__PTR3) );
  INV_X1 U4006 ( .A(_01831_), .ZN(_02629_) );
  INV_X1 U4007 ( .A(_01832_), .ZN(_02628_) );
  INV_X1 U4008 ( .A(_01833_), .ZN(_02603_) );
  INV_X1 U4009 ( .A(_00001_), .ZN(_02602_) );
  MUX2_X1 U4010 ( .A(1'b0), .B(_02117__PTR0), .S(_02927_), .Z(_01938__PTR320) );
  MUX2_X1 U4011 ( .A(1'b0), .B(_02117__PTR1), .S(_02927_), .Z(_01938__PTR321) );
  MUX2_X1 U4012 ( .A(1'b0), .B(_02117__PTR2), .S(_02927_), .Z(_01938__PTR322) );
  MUX2_X1 U4013 ( .A(1'b0), .B(_02117__PTR3), .S(_02927_), .Z(_01938__PTR323) );
  MUX2_X1 U4014 ( .A(1'b0), .B(_02117__PTR4), .S(_02927_), .Z(_01938__PTR324) );
  MUX2_X1 U4015 ( .A(1'b0), .B(_02117__PTR5), .S(_02927_), .Z(_01938__PTR325) );
  MUX2_X1 U4016 ( .A(1'b0), .B(_02117__PTR6), .S(_02927_), .Z(_01938__PTR326) );
  MUX2_X1 U4017 ( .A(1'b0), .B(_02117__PTR7), .S(_02927_), .Z(_01938__PTR327) );
  MUX2_X1 U4018 ( .A(1'b0), .B(_02117__PTR8), .S(_02927_), .Z(_01938__PTR328) );
  MUX2_X1 U4019 ( .A(1'b0), .B(_02117__PTR9), .S(_02927_), .Z(_01938__PTR329) );
  MUX2_X1 U4020 ( .A(1'b0), .B(_02117__PTR10), .S(_02927_), .Z(_01938__PTR330) );
  MUX2_X1 U4021 ( .A(1'b0), .B(_02117__PTR11), .S(_02927_), .Z(_01938__PTR331) );
  MUX2_X1 U4022 ( .A(1'b0), .B(_02117__PTR12), .S(_02927_), .Z(_01938__PTR332) );
  MUX2_X1 U4023 ( .A(1'b0), .B(_02117__PTR13), .S(_02927_), .Z(_01938__PTR333) );
  MUX2_X1 U4024 ( .A(1'b0), .B(_02117__PTR14), .S(_02927_), .Z(_01938__PTR334) );
  MUX2_X1 U4025 ( .A(1'b0), .B(_02117__PTR15), .S(_02927_), .Z(_01938__PTR335) );
  MUX2_X1 U4026 ( .A(1'b0), .B(_02117__PTR16), .S(_02927_), .Z(_01938__PTR336) );
  MUX2_X1 U4027 ( .A(1'b0), .B(_02117__PTR17), .S(_02927_), .Z(_01938__PTR337) );
  MUX2_X1 U4028 ( .A(1'b0), .B(_02117__PTR18), .S(_02927_), .Z(_01938__PTR338) );
  MUX2_X1 U4029 ( .A(1'b0), .B(_02117__PTR19), .S(_02927_), .Z(_01938__PTR339) );
  MUX2_X1 U4030 ( .A(1'b0), .B(_02117__PTR20), .S(_02927_), .Z(_01938__PTR340) );
  MUX2_X1 U4031 ( .A(1'b0), .B(_02117__PTR21), .S(_02927_), .Z(_01938__PTR341) );
  MUX2_X1 U4032 ( .A(1'b0), .B(_02117__PTR22), .S(_02927_), .Z(_01938__PTR342) );
  MUX2_X1 U4033 ( .A(1'b0), .B(_02117__PTR23), .S(_02927_), .Z(_01938__PTR343) );
  MUX2_X1 U4034 ( .A(1'b0), .B(_02117__PTR24), .S(_02927_), .Z(_01938__PTR344) );
  MUX2_X1 U4035 ( .A(1'b0), .B(_02117__PTR25), .S(_02927_), .Z(_01938__PTR345) );
  MUX2_X1 U4036 ( .A(1'b0), .B(_02117__PTR26), .S(_02927_), .Z(_01938__PTR346) );
  MUX2_X1 U4037 ( .A(1'b0), .B(_02117__PTR27), .S(_02927_), .Z(_01938__PTR347) );
  MUX2_X1 U4038 ( .A(1'b0), .B(_02117__PTR28), .S(_02927_), .Z(_01938__PTR348) );
  MUX2_X1 U4039 ( .A(1'b0), .B(_02117__PTR29), .S(_02927_), .Z(_01938__PTR349) );
  MUX2_X1 U4040 ( .A(1'b0), .B(_02117__PTR30), .S(_02927_), .Z(_01938__PTR350) );
  MUX2_X1 U4041 ( .A(1'b0), .B(_02117__PTR31), .S(_02927_), .Z(_01938__PTR352) );
  MUX2_X1 U4042 ( .A(1'b0), .B(_02113__PTR0), .S(_02926_), .Z(_01937__PTR80) );
  MUX2_X1 U4043 ( .A(1'b0), .B(_02113__PTR1), .S(_02926_), .Z(_01937__PTR81) );
  MUX2_X1 U4044 ( .A(1'b0), .B(_02113__PTR2), .S(_02926_), .Z(_01937__PTR82) );
  MUX2_X1 U4045 ( .A(1'b0), .B(_02113__PTR3), .S(_02926_), .Z(_01937__PTR83) );
  MUX2_X1 U4046 ( .A(1'b0), .B(_02113__PTR4), .S(_02926_), .Z(_01937__PTR84) );
  MUX2_X1 U4047 ( .A(1'b0), .B(_02113__PTR5), .S(_02926_), .Z(_01937__PTR85) );
  MUX2_X1 U4048 ( .A(1'b0), .B(_02113__PTR6), .S(_02926_), .Z(_01937__PTR86) );
  MUX2_X1 U4049 ( .A(1'b0), .B(_02113__PTR7), .S(_02926_), .Z(_01937__PTR87) );
  MUX2_X1 U4050 ( .A(1'b0), .B(_02113__PTR8), .S(_02926_), .Z(_01937__PTR88) );
  MUX2_X1 U4051 ( .A(1'b0), .B(_02113__PTR9), .S(_02926_), .Z(_01937__PTR89) );
  MUX2_X1 U4052 ( .A(1'b0), .B(_02113__PTR10), .S(_02926_), .Z(_01937__PTR90) );
  MUX2_X1 U4053 ( .A(1'b0), .B(_02113__PTR11), .S(_02926_), .Z(_01937__PTR91) );
  MUX2_X1 U4054 ( .A(1'b0), .B(_02113__PTR12), .S(_02926_), .Z(_01937__PTR92) );
  MUX2_X1 U4055 ( .A(1'b0), .B(_02113__PTR13), .S(_02926_), .Z(_01937__PTR93) );
  MUX2_X1 U4056 ( .A(1'b0), .B(_02113__PTR14), .S(_02926_), .Z(_01937__PTR94) );
  MUX2_X1 U4057 ( .A(1'b0), .B(_02113__PTR15), .S(_02926_), .Z(_01937__PTR95) );
  MUX2_X1 U4058 ( .A(1'b0), .B(_02110__PTR0), .S(_02926_), .Z(_01936__PTR80) );
  MUX2_X1 U4059 ( .A(1'b0), .B(_02110__PTR1), .S(_02926_), .Z(_01936__PTR81) );
  MUX2_X1 U4060 ( .A(1'b0), .B(_02110__PTR2), .S(_02926_), .Z(_01936__PTR82) );
  MUX2_X1 U4061 ( .A(1'b0), .B(_02110__PTR3), .S(_02926_), .Z(_01936__PTR83) );
  MUX2_X1 U4062 ( .A(1'b0), .B(_02110__PTR4), .S(_02926_), .Z(_01936__PTR84) );
  MUX2_X1 U4063 ( .A(1'b0), .B(_02110__PTR5), .S(_02926_), .Z(_01936__PTR85) );
  MUX2_X1 U4064 ( .A(1'b0), .B(_02110__PTR6), .S(_02926_), .Z(_01936__PTR86) );
  MUX2_X1 U4065 ( .A(1'b0), .B(_02110__PTR7), .S(_02926_), .Z(_01936__PTR87) );
  MUX2_X1 U4066 ( .A(1'b0), .B(_02110__PTR8), .S(_02926_), .Z(_01936__PTR88) );
  MUX2_X1 U4067 ( .A(1'b0), .B(_02110__PTR9), .S(_02926_), .Z(_01936__PTR89) );
  MUX2_X1 U4068 ( .A(1'b0), .B(_02110__PTR10), .S(_02926_), .Z(_01936__PTR90) );
  MUX2_X1 U4069 ( .A(1'b0), .B(_02110__PTR11), .S(_02926_), .Z(_01936__PTR91) );
  MUX2_X1 U4070 ( .A(1'b0), .B(_02110__PTR12), .S(_02926_), .Z(_01936__PTR92) );
  MUX2_X1 U4071 ( .A(1'b0), .B(_02110__PTR13), .S(_02926_), .Z(_01936__PTR93) );
  MUX2_X1 U4072 ( .A(1'b0), .B(_02110__PTR14), .S(_02926_), .Z(_01936__PTR94) );
  MUX2_X1 U4073 ( .A(1'b0), .B(_02103__PTR0), .S(_02924_), .Z(_01935__PTR160) );
  MUX2_X1 U4074 ( .A(1'b0), .B(_02103__PTR1), .S(_02924_), .Z(_01935__PTR161) );
  MUX2_X1 U4075 ( .A(1'b0), .B(_02103__PTR2), .S(_02924_), .Z(_01935__PTR162) );
  MUX2_X1 U4076 ( .A(1'b0), .B(_02103__PTR3), .S(_02924_), .Z(_01935__PTR163) );
  MUX2_X1 U4077 ( .A(1'b0), .B(_02103__PTR4), .S(_02924_), .Z(_01935__PTR164) );
  MUX2_X1 U4078 ( .A(1'b0), .B(_02103__PTR5), .S(_02924_), .Z(_01935__PTR165) );
  MUX2_X1 U4079 ( .A(1'b0), .B(_02103__PTR6), .S(_02924_), .Z(_01935__PTR166) );
  MUX2_X1 U4080 ( .A(1'b0), .B(_02103__PTR7), .S(_02924_), .Z(_01935__PTR167) );
  MUX2_X1 U4081 ( .A(1'b0), .B(_02103__PTR8), .S(_02924_), .Z(_01935__PTR168) );
  MUX2_X1 U4082 ( .A(1'b0), .B(_02103__PTR9), .S(_02924_), .Z(_01935__PTR169) );
  MUX2_X1 U4083 ( .A(1'b0), .B(_02103__PTR10), .S(_02924_), .Z(_01935__PTR170) );
  MUX2_X1 U4084 ( .A(1'b0), .B(_02103__PTR11), .S(_02924_), .Z(_01935__PTR171) );
  MUX2_X1 U4085 ( .A(1'b0), .B(_02103__PTR12), .S(_02924_), .Z(_01935__PTR172) );
  MUX2_X1 U4086 ( .A(1'b0), .B(_02103__PTR13), .S(_02924_), .Z(_01935__PTR173) );
  MUX2_X1 U4087 ( .A(1'b0), .B(_02103__PTR14), .S(_02924_), .Z(_01935__PTR174) );
  MUX2_X1 U4088 ( .A(1'b0), .B(_02103__PTR15), .S(_02924_), .Z(_01935__PTR175) );
  MUX2_X1 U4089 ( .A(1'b0), .B(_02103__PTR16), .S(_02924_), .Z(_01935__PTR176) );
  MUX2_X1 U4090 ( .A(1'b0), .B(_02103__PTR17), .S(_02924_), .Z(_01935__PTR177) );
  MUX2_X1 U4091 ( .A(1'b0), .B(_02103__PTR18), .S(_02924_), .Z(_01935__PTR178) );
  MUX2_X1 U4092 ( .A(1'b0), .B(_02103__PTR19), .S(_02924_), .Z(_01935__PTR179) );
  MUX2_X1 U4093 ( .A(1'b0), .B(_02103__PTR20), .S(_02924_), .Z(_01935__PTR180) );
  MUX2_X1 U4094 ( .A(1'b0), .B(_02103__PTR21), .S(_02924_), .Z(_01935__PTR181) );
  MUX2_X1 U4095 ( .A(1'b0), .B(_02103__PTR22), .S(_02924_), .Z(_01935__PTR182) );
  MUX2_X1 U4096 ( .A(1'b0), .B(_02103__PTR23), .S(_02924_), .Z(_01935__PTR183) );
  MUX2_X1 U4097 ( .A(1'b0), .B(_02103__PTR24), .S(_02924_), .Z(_01935__PTR184) );
  MUX2_X1 U4098 ( .A(1'b0), .B(_02103__PTR25), .S(_02924_), .Z(_01935__PTR185) );
  MUX2_X1 U4099 ( .A(1'b0), .B(_02103__PTR26), .S(_02924_), .Z(_01935__PTR186) );
  MUX2_X1 U4100 ( .A(1'b0), .B(_02103__PTR27), .S(_02924_), .Z(_01935__PTR187) );
  MUX2_X1 U4101 ( .A(1'b0), .B(_02103__PTR28), .S(_02924_), .Z(_01935__PTR188) );
  MUX2_X1 U4102 ( .A(1'b0), .B(_02103__PTR29), .S(_02924_), .Z(_01935__PTR189) );
  MUX2_X1 U4103 ( .A(1'b0), .B(_02103__PTR30), .S(_02924_), .Z(_01935__PTR190) );
  MUX2_X1 U4104 ( .A(1'b0), .B(_02103__PTR31), .S(_02924_), .Z(_01935__PTR191) );
  MUX2_X1 U4105 ( .A(1'b0), .B(_02099__PTR0), .S(_02923_), .Z(_01934__PTR160) );
  MUX2_X1 U4106 ( .A(1'b0), .B(_02099__PTR1), .S(_02923_), .Z(_01934__PTR161) );
  MUX2_X1 U4107 ( .A(1'b0), .B(_02099__PTR2), .S(_02923_), .Z(_01934__PTR162) );
  MUX2_X1 U4108 ( .A(1'b0), .B(_02099__PTR3), .S(_02923_), .Z(_01934__PTR163) );
  MUX2_X1 U4109 ( .A(1'b0), .B(_02099__PTR4), .S(_02923_), .Z(_01934__PTR164) );
  MUX2_X1 U4110 ( .A(1'b0), .B(_02099__PTR5), .S(_02923_), .Z(_01934__PTR165) );
  MUX2_X1 U4111 ( .A(1'b0), .B(_02099__PTR6), .S(_02923_), .Z(_01934__PTR166) );
  MUX2_X1 U4112 ( .A(1'b0), .B(_02099__PTR7), .S(_02923_), .Z(_01934__PTR167) );
  MUX2_X1 U4113 ( .A(1'b0), .B(_02099__PTR8), .S(_02923_), .Z(_01934__PTR168) );
  MUX2_X1 U4114 ( .A(1'b0), .B(_02099__PTR9), .S(_02923_), .Z(_01934__PTR169) );
  MUX2_X1 U4115 ( .A(1'b0), .B(_02099__PTR10), .S(_02923_), .Z(_01934__PTR170) );
  MUX2_X1 U4116 ( .A(1'b0), .B(_02099__PTR11), .S(_02923_), .Z(_01934__PTR171) );
  MUX2_X1 U4117 ( .A(1'b0), .B(_02099__PTR12), .S(_02923_), .Z(_01934__PTR172) );
  MUX2_X1 U4118 ( .A(1'b0), .B(_02099__PTR13), .S(_02923_), .Z(_01934__PTR173) );
  MUX2_X1 U4119 ( .A(1'b0), .B(_02099__PTR14), .S(_02923_), .Z(_01934__PTR174) );
  MUX2_X1 U4120 ( .A(1'b0), .B(_02099__PTR15), .S(_02923_), .Z(_01934__PTR175) );
  MUX2_X1 U4121 ( .A(1'b0), .B(_02099__PTR16), .S(_02923_), .Z(_01934__PTR176) );
  MUX2_X1 U4122 ( .A(1'b0), .B(_02099__PTR17), .S(_02923_), .Z(_01934__PTR177) );
  MUX2_X1 U4123 ( .A(1'b0), .B(_02099__PTR18), .S(_02923_), .Z(_01934__PTR178) );
  MUX2_X1 U4124 ( .A(1'b0), .B(_02099__PTR19), .S(_02923_), .Z(_01934__PTR179) );
  MUX2_X1 U4125 ( .A(1'b0), .B(_02099__PTR20), .S(_02923_), .Z(_01934__PTR180) );
  MUX2_X1 U4126 ( .A(1'b0), .B(_02099__PTR21), .S(_02923_), .Z(_01934__PTR181) );
  MUX2_X1 U4127 ( .A(1'b0), .B(_02099__PTR22), .S(_02923_), .Z(_01934__PTR182) );
  MUX2_X1 U4128 ( .A(1'b0), .B(_02099__PTR23), .S(_02923_), .Z(_01934__PTR183) );
  MUX2_X1 U4129 ( .A(1'b0), .B(_02099__PTR24), .S(_02923_), .Z(_01934__PTR184) );
  MUX2_X1 U4130 ( .A(1'b0), .B(_02099__PTR25), .S(_02923_), .Z(_01934__PTR185) );
  MUX2_X1 U4131 ( .A(1'b0), .B(_02099__PTR26), .S(_02923_), .Z(_01934__PTR186) );
  MUX2_X1 U4132 ( .A(1'b0), .B(_02099__PTR27), .S(_02923_), .Z(_01934__PTR187) );
  MUX2_X1 U4133 ( .A(1'b0), .B(_02099__PTR28), .S(_02923_), .Z(_01934__PTR188) );
  MUX2_X1 U4134 ( .A(1'b0), .B(_02099__PTR29), .S(_02923_), .Z(_01934__PTR189) );
  MUX2_X1 U4135 ( .A(1'b0), .B(_02099__PTR30), .S(_02923_), .Z(_01934__PTR190) );
  MUX2_X1 U4136 ( .A(1'b0), .B(_02099__PTR31), .S(_02923_), .Z(_01934__PTR191) );
  MUX2_X1 U4137 ( .A(1'b0), .B(_01860_), .S(_02773_), .Z(_01852__PTR5) );
  MUX2_X1 U4138 ( .A(1'b0), .B(_01856_), .S(_02772_), .Z(_01851__PTR5) );
  MUX2_X1 U4139 ( .A(1'b0), .B(_02091__PTR0), .S(_02921_), .Z(_01932__PTR40) );
  MUX2_X1 U4140 ( .A(1'b0), .B(_02091__PTR1), .S(_02921_), .Z(_01932__PTR41) );
  MUX2_X1 U4141 ( .A(1'b0), .B(_02091__PTR2), .S(_02921_), .Z(_01932__PTR42) );
  MUX2_X1 U4142 ( .A(1'b0), .B(_02091__PTR3), .S(_02921_), .Z(_01932__PTR43) );
  MUX2_X1 U4143 ( .A(1'b0), .B(_02091__PTR4), .S(_02921_), .Z(_01932__PTR44) );
  MUX2_X1 U4144 ( .A(1'b0), .B(_01875_), .S(_02776_), .Z(_01850__PTR5) );
  MUX2_X1 U4145 ( .A(1'b0), .B(_01864_), .S(_02774_), .Z(_01849__PTR5) );
  MUX2_X1 U4146 ( .A(1'b0), .B(_01871_), .S(_02776_), .Z(_01848__PTR5) );
  MUX2_X1 U4147 ( .A(1'b0), .B(_01867_), .S(_02775_), .Z(_01847__PTR5) );
  MUX2_X1 U4148 ( .A(1'b0), .B(_02106__PTR0), .S(_02925_), .Z(_01896__PTR320) );
  MUX2_X1 U4149 ( .A(1'b0), .B(_02106__PTR1), .S(_02925_), .Z(_01896__PTR321) );
  MUX2_X1 U4150 ( .A(1'b0), .B(_02106__PTR2), .S(_02925_), .Z(_01896__PTR322) );
  MUX2_X1 U4151 ( .A(1'b0), .B(_02106__PTR3), .S(_02925_), .Z(_01896__PTR323) );
  MUX2_X1 U4152 ( .A(1'b0), .B(_02106__PTR4), .S(_02925_), .Z(_01896__PTR324) );
  MUX2_X1 U4153 ( .A(1'b0), .B(_02106__PTR5), .S(_02925_), .Z(_01896__PTR325) );
  MUX2_X1 U4154 ( .A(1'b0), .B(_02106__PTR6), .S(_02925_), .Z(_01896__PTR326) );
  MUX2_X1 U4155 ( .A(1'b0), .B(_02106__PTR7), .S(_02925_), .Z(_01896__PTR327) );
  MUX2_X1 U4156 ( .A(1'b0), .B(_02106__PTR8), .S(_02925_), .Z(_01896__PTR328) );
  MUX2_X1 U4157 ( .A(1'b0), .B(_02106__PTR9), .S(_02925_), .Z(_01896__PTR329) );
  MUX2_X1 U4158 ( .A(1'b0), .B(_02106__PTR10), .S(_02925_), .Z(_01896__PTR330) );
  MUX2_X1 U4159 ( .A(1'b0), .B(_02106__PTR11), .S(_02925_), .Z(_01896__PTR331) );
  MUX2_X1 U4160 ( .A(1'b0), .B(_02106__PTR12), .S(_02925_), .Z(_01896__PTR332) );
  MUX2_X1 U4161 ( .A(1'b0), .B(_02106__PTR13), .S(_02925_), .Z(_01896__PTR333) );
  MUX2_X1 U4162 ( .A(1'b0), .B(_02106__PTR14), .S(_02925_), .Z(_01896__PTR334) );
  MUX2_X1 U4163 ( .A(1'b0), .B(_02106__PTR15), .S(_02925_), .Z(_01896__PTR335) );
  MUX2_X1 U4164 ( .A(1'b0), .B(_02106__PTR16), .S(_02925_), .Z(_01896__PTR336) );
  MUX2_X1 U4165 ( .A(1'b0), .B(_02106__PTR17), .S(_02925_), .Z(_01896__PTR337) );
  MUX2_X1 U4166 ( .A(1'b0), .B(_02106__PTR18), .S(_02925_), .Z(_01896__PTR338) );
  MUX2_X1 U4167 ( .A(1'b0), .B(_02106__PTR19), .S(_02925_), .Z(_01896__PTR339) );
  MUX2_X1 U4168 ( .A(1'b0), .B(_02106__PTR20), .S(_02925_), .Z(_01896__PTR340) );
  MUX2_X1 U4169 ( .A(1'b0), .B(_02106__PTR21), .S(_02925_), .Z(_01896__PTR341) );
  MUX2_X1 U4170 ( .A(1'b0), .B(_02106__PTR22), .S(_02925_), .Z(_01896__PTR342) );
  MUX2_X1 U4171 ( .A(1'b0), .B(_02106__PTR23), .S(_02925_), .Z(_01896__PTR343) );
  MUX2_X1 U4172 ( .A(1'b0), .B(_02106__PTR24), .S(_02925_), .Z(_01896__PTR344) );
  MUX2_X1 U4173 ( .A(1'b0), .B(_02106__PTR25), .S(_02925_), .Z(_01896__PTR345) );
  MUX2_X1 U4174 ( .A(1'b0), .B(_02106__PTR26), .S(_02925_), .Z(_01896__PTR346) );
  MUX2_X1 U4175 ( .A(1'b0), .B(_02106__PTR27), .S(_02925_), .Z(_01896__PTR347) );
  MUX2_X1 U4176 ( .A(1'b0), .B(_02106__PTR28), .S(_02925_), .Z(_01896__PTR348) );
  MUX2_X1 U4177 ( .A(1'b0), .B(_02106__PTR29), .S(_02925_), .Z(_01896__PTR349) );
  MUX2_X1 U4178 ( .A(1'b0), .B(_02106__PTR30), .S(_02925_), .Z(_01896__PTR350) );
  MUX2_X1 U4179 ( .A(1'b0), .B(_02106__PTR31), .S(_02925_), .Z(_01896__PTR352) );
  MUX2_X1 U4180 ( .A(1'b0), .B(_02087__PTR0), .S(_02920_), .Z(_01893__PTR160) );
  MUX2_X1 U4181 ( .A(1'b0), .B(_02087__PTR1), .S(_02920_), .Z(_01893__PTR161) );
  MUX2_X1 U4182 ( .A(1'b0), .B(_02087__PTR2), .S(_02920_), .Z(_01893__PTR162) );
  MUX2_X1 U4183 ( .A(1'b0), .B(_02087__PTR3), .S(_02920_), .Z(_01893__PTR163) );
  MUX2_X1 U4184 ( .A(1'b0), .B(_02087__PTR4), .S(_02920_), .Z(_01893__PTR164) );
  MUX2_X1 U4185 ( .A(1'b0), .B(_02087__PTR5), .S(_02920_), .Z(_01893__PTR165) );
  MUX2_X1 U4186 ( .A(1'b0), .B(_02087__PTR6), .S(_02920_), .Z(_01893__PTR166) );
  MUX2_X1 U4187 ( .A(1'b0), .B(_02087__PTR7), .S(_02920_), .Z(_01893__PTR167) );
  MUX2_X1 U4188 ( .A(1'b0), .B(_02087__PTR8), .S(_02920_), .Z(_01893__PTR168) );
  MUX2_X1 U4189 ( .A(1'b0), .B(_02087__PTR9), .S(_02920_), .Z(_01893__PTR169) );
  MUX2_X1 U4190 ( .A(1'b0), .B(_02087__PTR10), .S(_02920_), .Z(_01893__PTR170) );
  MUX2_X1 U4191 ( .A(1'b0), .B(_02087__PTR11), .S(_02920_), .Z(_01893__PTR171) );
  MUX2_X1 U4192 ( .A(1'b0), .B(_02087__PTR12), .S(_02920_), .Z(_01893__PTR172) );
  MUX2_X1 U4193 ( .A(1'b0), .B(_02087__PTR13), .S(_02920_), .Z(_01893__PTR173) );
  MUX2_X1 U4194 ( .A(1'b0), .B(_02087__PTR14), .S(_02920_), .Z(_01893__PTR174) );
  MUX2_X1 U4195 ( .A(1'b0), .B(_02087__PTR15), .S(_02920_), .Z(_01893__PTR175) );
  MUX2_X1 U4196 ( .A(1'b0), .B(_02087__PTR16), .S(_02920_), .Z(_01893__PTR176) );
  MUX2_X1 U4197 ( .A(1'b0), .B(_02087__PTR17), .S(_02920_), .Z(_01893__PTR177) );
  MUX2_X1 U4198 ( .A(1'b0), .B(_02087__PTR18), .S(_02920_), .Z(_01893__PTR178) );
  MUX2_X1 U4199 ( .A(1'b0), .B(_02087__PTR19), .S(_02920_), .Z(_01893__PTR179) );
  MUX2_X1 U4200 ( .A(1'b0), .B(_02087__PTR20), .S(_02920_), .Z(_01893__PTR180) );
  MUX2_X1 U4201 ( .A(1'b0), .B(_02087__PTR21), .S(_02920_), .Z(_01893__PTR181) );
  MUX2_X1 U4202 ( .A(1'b0), .B(_02087__PTR22), .S(_02920_), .Z(_01893__PTR182) );
  MUX2_X1 U4203 ( .A(1'b0), .B(_02087__PTR23), .S(_02920_), .Z(_01893__PTR183) );
  MUX2_X1 U4204 ( .A(1'b0), .B(_02087__PTR24), .S(_02920_), .Z(_01893__PTR184) );
  MUX2_X1 U4205 ( .A(1'b0), .B(_02087__PTR25), .S(_02920_), .Z(_01893__PTR185) );
  MUX2_X1 U4206 ( .A(1'b0), .B(_02087__PTR26), .S(_02920_), .Z(_01893__PTR186) );
  MUX2_X1 U4207 ( .A(1'b0), .B(_02087__PTR27), .S(_02920_), .Z(_01893__PTR187) );
  MUX2_X1 U4208 ( .A(1'b0), .B(_02087__PTR28), .S(_02920_), .Z(_01893__PTR188) );
  MUX2_X1 U4209 ( .A(1'b0), .B(_02087__PTR29), .S(_02920_), .Z(_01893__PTR189) );
  MUX2_X1 U4210 ( .A(1'b0), .B(_02087__PTR30), .S(_02920_), .Z(_01893__PTR190) );
  MUX2_X1 U4211 ( .A(1'b0), .B(_02087__PTR31), .S(_02920_), .Z(_01893__PTR191) );
  MUX2_X1 U4212 ( .A(1'b0), .B(_02095__PTR0), .S(_02922_), .Z(_01892__PTR160) );
  MUX2_X1 U4213 ( .A(1'b0), .B(_02095__PTR1), .S(_02922_), .Z(_01892__PTR161) );
  MUX2_X1 U4214 ( .A(1'b0), .B(_02095__PTR2), .S(_02922_), .Z(_01892__PTR162) );
  MUX2_X1 U4215 ( .A(1'b0), .B(_02095__PTR3), .S(_02922_), .Z(_01892__PTR163) );
  MUX2_X1 U4216 ( .A(1'b0), .B(_02095__PTR4), .S(_02922_), .Z(_01892__PTR164) );
  MUX2_X1 U4217 ( .A(1'b0), .B(_02095__PTR5), .S(_02922_), .Z(_01892__PTR165) );
  MUX2_X1 U4218 ( .A(1'b0), .B(_02095__PTR6), .S(_02922_), .Z(_01892__PTR166) );
  MUX2_X1 U4219 ( .A(1'b0), .B(_02095__PTR7), .S(_02922_), .Z(_01892__PTR167) );
  MUX2_X1 U4220 ( .A(1'b0), .B(_02095__PTR8), .S(_02922_), .Z(_01892__PTR168) );
  MUX2_X1 U4221 ( .A(1'b0), .B(_02095__PTR9), .S(_02922_), .Z(_01892__PTR169) );
  MUX2_X1 U4222 ( .A(1'b0), .B(_02095__PTR10), .S(_02922_), .Z(_01892__PTR170) );
  MUX2_X1 U4223 ( .A(1'b0), .B(_02095__PTR11), .S(_02922_), .Z(_01892__PTR171) );
  MUX2_X1 U4224 ( .A(1'b0), .B(_02095__PTR12), .S(_02922_), .Z(_01892__PTR172) );
  MUX2_X1 U4225 ( .A(1'b0), .B(_02095__PTR13), .S(_02922_), .Z(_01892__PTR173) );
  MUX2_X1 U4226 ( .A(1'b0), .B(_02095__PTR14), .S(_02922_), .Z(_01892__PTR174) );
  MUX2_X1 U4227 ( .A(1'b0), .B(_02095__PTR15), .S(_02922_), .Z(_01892__PTR175) );
  MUX2_X1 U4228 ( .A(1'b0), .B(_02095__PTR16), .S(_02922_), .Z(_01892__PTR176) );
  MUX2_X1 U4229 ( .A(1'b0), .B(_02095__PTR17), .S(_02922_), .Z(_01892__PTR177) );
  MUX2_X1 U4230 ( .A(1'b0), .B(_02095__PTR18), .S(_02922_), .Z(_01892__PTR178) );
  MUX2_X1 U4231 ( .A(1'b0), .B(_02095__PTR19), .S(_02922_), .Z(_01892__PTR179) );
  MUX2_X1 U4232 ( .A(1'b0), .B(_02095__PTR20), .S(_02922_), .Z(_01892__PTR180) );
  MUX2_X1 U4233 ( .A(1'b0), .B(_02095__PTR21), .S(_02922_), .Z(_01892__PTR181) );
  MUX2_X1 U4234 ( .A(1'b0), .B(_02095__PTR22), .S(_02922_), .Z(_01892__PTR182) );
  MUX2_X1 U4235 ( .A(1'b0), .B(_02095__PTR23), .S(_02922_), .Z(_01892__PTR183) );
  MUX2_X1 U4236 ( .A(1'b0), .B(_02095__PTR24), .S(_02922_), .Z(_01892__PTR184) );
  MUX2_X1 U4237 ( .A(1'b0), .B(_02095__PTR25), .S(_02922_), .Z(_01892__PTR185) );
  MUX2_X1 U4238 ( .A(1'b0), .B(_02095__PTR26), .S(_02922_), .Z(_01892__PTR186) );
  MUX2_X1 U4239 ( .A(1'b0), .B(_02095__PTR27), .S(_02922_), .Z(_01892__PTR187) );
  MUX2_X1 U4240 ( .A(1'b0), .B(_02095__PTR28), .S(_02922_), .Z(_01892__PTR188) );
  MUX2_X1 U4241 ( .A(1'b0), .B(_02095__PTR29), .S(_02922_), .Z(_01892__PTR189) );
  MUX2_X1 U4242 ( .A(1'b0), .B(_02095__PTR30), .S(_02922_), .Z(_01892__PTR190) );
  MUX2_X1 U4243 ( .A(1'b0), .B(_02095__PTR31), .S(_02922_), .Z(_01892__PTR191) );
  MUX2_X1 U4244 ( .A(1'b0), .B(_02122__PTR0), .S(_02928_), .Z(_02121__PTR0) );
  MUX2_X1 U4245 ( .A(1'b0), .B(_02122__PTR1), .S(_02928_), .Z(_02121__PTR1) );
  MUX2_X1 U4246 ( .A(1'b0), .B(_02122__PTR2), .S(_02928_), .Z(_02121__PTR2) );
  MUX2_X1 U4247 ( .A(1'b0), .B(_02122__PTR3), .S(_02928_), .Z(_02121__PTR3) );
  MUX2_X1 U4248 ( .A(1'b0), .B(_02415__PTR0), .S(_03174_), .Z(_02414__PTR0) );
  MUX2_X1 U4249 ( .A(1'b0), .B(_02415__PTR1), .S(_03174_), .Z(_02414__PTR1) );
  MUX2_X1 U4250 ( .A(1'b0), .B(_02415__PTR2), .S(_03174_), .Z(_02414__PTR2) );
  MUX2_X1 U4251 ( .A(1'b0), .B(_02415__PTR3), .S(_03174_), .Z(_02414__PTR3) );
  MUX2_X1 U4252 ( .A(1'b0), .B(_02406__PTR0), .S(_03172_), .Z(_02230__PTR320) );
  MUX2_X1 U4253 ( .A(1'b0), .B(_02406__PTR1), .S(_03172_), .Z(_02230__PTR321) );
  MUX2_X1 U4254 ( .A(1'b0), .B(_02406__PTR2), .S(_03172_), .Z(_02230__PTR322) );
  MUX2_X1 U4255 ( .A(1'b0), .B(_02406__PTR3), .S(_03172_), .Z(_02230__PTR323) );
  MUX2_X1 U4256 ( .A(1'b0), .B(_02406__PTR4), .S(_03172_), .Z(_02230__PTR324) );
  MUX2_X1 U4257 ( .A(1'b0), .B(_02406__PTR5), .S(_03172_), .Z(_02230__PTR325) );
  MUX2_X1 U4258 ( .A(1'b0), .B(_02406__PTR6), .S(_03172_), .Z(_02230__PTR326) );
  MUX2_X1 U4259 ( .A(1'b0), .B(_02406__PTR7), .S(_03172_), .Z(_02230__PTR327) );
  MUX2_X1 U4260 ( .A(1'b0), .B(_02406__PTR8), .S(_03172_), .Z(_02230__PTR328) );
  MUX2_X1 U4261 ( .A(1'b0), .B(_02406__PTR9), .S(_03172_), .Z(_02230__PTR329) );
  MUX2_X1 U4262 ( .A(1'b0), .B(_02406__PTR10), .S(_03172_), .Z(_02230__PTR330) );
  MUX2_X1 U4263 ( .A(1'b0), .B(_02406__PTR11), .S(_03172_), .Z(_02230__PTR331) );
  MUX2_X1 U4264 ( .A(1'b0), .B(_02406__PTR12), .S(_03172_), .Z(_02230__PTR332) );
  MUX2_X1 U4265 ( .A(1'b0), .B(_02406__PTR13), .S(_03172_), .Z(_02230__PTR333) );
  MUX2_X1 U4266 ( .A(1'b0), .B(_02406__PTR14), .S(_03172_), .Z(_02230__PTR334) );
  MUX2_X1 U4267 ( .A(1'b0), .B(_02406__PTR15), .S(_03172_), .Z(_02230__PTR335) );
  MUX2_X1 U4268 ( .A(1'b0), .B(_02406__PTR16), .S(_03172_), .Z(_02230__PTR336) );
  MUX2_X1 U4269 ( .A(1'b0), .B(_02406__PTR17), .S(_03172_), .Z(_02230__PTR337) );
  MUX2_X1 U4270 ( .A(1'b0), .B(_02406__PTR18), .S(_03172_), .Z(_02230__PTR338) );
  MUX2_X1 U4271 ( .A(1'b0), .B(_02406__PTR19), .S(_03172_), .Z(_02230__PTR339) );
  MUX2_X1 U4272 ( .A(1'b0), .B(_02406__PTR20), .S(_03172_), .Z(_02230__PTR340) );
  MUX2_X1 U4273 ( .A(1'b0), .B(_02406__PTR21), .S(_03172_), .Z(_02230__PTR341) );
  MUX2_X1 U4274 ( .A(1'b0), .B(_02406__PTR22), .S(_03172_), .Z(_02230__PTR342) );
  MUX2_X1 U4275 ( .A(1'b0), .B(_02406__PTR23), .S(_03172_), .Z(_02230__PTR343) );
  MUX2_X1 U4276 ( .A(1'b0), .B(_02406__PTR24), .S(_03172_), .Z(_02230__PTR344) );
  MUX2_X1 U4277 ( .A(1'b0), .B(_02406__PTR25), .S(_03172_), .Z(_02230__PTR345) );
  MUX2_X1 U4278 ( .A(1'b0), .B(_02406__PTR26), .S(_03172_), .Z(_02230__PTR346) );
  MUX2_X1 U4279 ( .A(1'b0), .B(_02406__PTR27), .S(_03172_), .Z(_02230__PTR347) );
  MUX2_X1 U4280 ( .A(1'b0), .B(_02406__PTR28), .S(_03172_), .Z(_02230__PTR348) );
  MUX2_X1 U4281 ( .A(1'b0), .B(_02406__PTR29), .S(_03172_), .Z(_02230__PTR349) );
  MUX2_X1 U4282 ( .A(1'b0), .B(_02406__PTR30), .S(_03172_), .Z(_02230__PTR350) );
  MUX2_X1 U4283 ( .A(1'b0), .B(_02406__PTR31), .S(_03172_), .Z(_02230__PTR352) );
  MUX2_X1 U4284 ( .A(1'b0), .B(_02402__PTR0), .S(_03171_), .Z(_02229__PTR80) );
  MUX2_X1 U4285 ( .A(1'b0), .B(_02402__PTR1), .S(_03171_), .Z(_02229__PTR81) );
  MUX2_X1 U4286 ( .A(1'b0), .B(_02402__PTR2), .S(_03171_), .Z(_02229__PTR82) );
  MUX2_X1 U4287 ( .A(1'b0), .B(_02402__PTR3), .S(_03171_), .Z(_02229__PTR83) );
  MUX2_X1 U4288 ( .A(1'b0), .B(_02402__PTR4), .S(_03171_), .Z(_02229__PTR84) );
  MUX2_X1 U4289 ( .A(1'b0), .B(_02402__PTR5), .S(_03171_), .Z(_02229__PTR85) );
  MUX2_X1 U4290 ( .A(1'b0), .B(_02402__PTR6), .S(_03171_), .Z(_02229__PTR86) );
  MUX2_X1 U4291 ( .A(1'b0), .B(_02402__PTR7), .S(_03171_), .Z(_02229__PTR87) );
  MUX2_X1 U4292 ( .A(1'b0), .B(_02402__PTR8), .S(_03171_), .Z(_02229__PTR88) );
  MUX2_X1 U4293 ( .A(1'b0), .B(_02402__PTR9), .S(_03171_), .Z(_02229__PTR89) );
  MUX2_X1 U4294 ( .A(1'b0), .B(_02402__PTR10), .S(_03171_), .Z(_02229__PTR90) );
  MUX2_X1 U4295 ( .A(1'b0), .B(_02402__PTR11), .S(_03171_), .Z(_02229__PTR91) );
  MUX2_X1 U4296 ( .A(1'b0), .B(_02402__PTR12), .S(_03171_), .Z(_02229__PTR92) );
  MUX2_X1 U4297 ( .A(1'b0), .B(_02402__PTR13), .S(_03171_), .Z(_02229__PTR93) );
  MUX2_X1 U4298 ( .A(1'b0), .B(_02402__PTR14), .S(_03171_), .Z(_02229__PTR94) );
  MUX2_X1 U4299 ( .A(1'b0), .B(_02402__PTR15), .S(_03171_), .Z(_02229__PTR95) );
  MUX2_X1 U4300 ( .A(1'b0), .B(_02399__PTR0), .S(_03171_), .Z(_02228__PTR80) );
  MUX2_X1 U4301 ( .A(1'b0), .B(_02399__PTR1), .S(_03171_), .Z(_02228__PTR81) );
  MUX2_X1 U4302 ( .A(1'b0), .B(_02399__PTR2), .S(_03171_), .Z(_02228__PTR82) );
  MUX2_X1 U4303 ( .A(1'b0), .B(_02399__PTR3), .S(_03171_), .Z(_02228__PTR83) );
  MUX2_X1 U4304 ( .A(1'b0), .B(_02399__PTR4), .S(_03171_), .Z(_02228__PTR84) );
  MUX2_X1 U4305 ( .A(1'b0), .B(_02399__PTR5), .S(_03171_), .Z(_02228__PTR85) );
  MUX2_X1 U4306 ( .A(1'b0), .B(_02399__PTR6), .S(_03171_), .Z(_02228__PTR86) );
  MUX2_X1 U4307 ( .A(1'b0), .B(_02399__PTR7), .S(_03171_), .Z(_02228__PTR87) );
  MUX2_X1 U4308 ( .A(1'b0), .B(_02399__PTR8), .S(_03171_), .Z(_02228__PTR88) );
  MUX2_X1 U4309 ( .A(1'b0), .B(_02399__PTR9), .S(_03171_), .Z(_02228__PTR89) );
  MUX2_X1 U4310 ( .A(1'b0), .B(_02399__PTR10), .S(_03171_), .Z(_02228__PTR90) );
  MUX2_X1 U4311 ( .A(1'b0), .B(_02399__PTR11), .S(_03171_), .Z(_02228__PTR91) );
  MUX2_X1 U4312 ( .A(1'b0), .B(_02399__PTR12), .S(_03171_), .Z(_02228__PTR92) );
  MUX2_X1 U4313 ( .A(1'b0), .B(_02399__PTR13), .S(_03171_), .Z(_02228__PTR93) );
  MUX2_X1 U4314 ( .A(1'b0), .B(_02399__PTR14), .S(_03171_), .Z(_02228__PTR94) );
  MUX2_X1 U4315 ( .A(1'b0), .B(_02392__PTR0), .S(_03169_), .Z(_02227__PTR160) );
  MUX2_X1 U4316 ( .A(1'b0), .B(_02392__PTR1), .S(_03169_), .Z(_02227__PTR161) );
  MUX2_X1 U4317 ( .A(1'b0), .B(_02392__PTR2), .S(_03169_), .Z(_02227__PTR162) );
  MUX2_X1 U4318 ( .A(1'b0), .B(_02392__PTR3), .S(_03169_), .Z(_02227__PTR163) );
  MUX2_X1 U4319 ( .A(1'b0), .B(_02392__PTR4), .S(_03169_), .Z(_02227__PTR164) );
  MUX2_X1 U4320 ( .A(1'b0), .B(_02392__PTR5), .S(_03169_), .Z(_02227__PTR165) );
  MUX2_X1 U4321 ( .A(1'b0), .B(_02392__PTR6), .S(_03169_), .Z(_02227__PTR166) );
  MUX2_X1 U4322 ( .A(1'b0), .B(_02392__PTR7), .S(_03169_), .Z(_02227__PTR167) );
  MUX2_X1 U4323 ( .A(1'b0), .B(_02392__PTR8), .S(_03169_), .Z(_02227__PTR168) );
  MUX2_X1 U4324 ( .A(1'b0), .B(_02392__PTR9), .S(_03169_), .Z(_02227__PTR169) );
  MUX2_X1 U4325 ( .A(1'b0), .B(_02392__PTR10), .S(_03169_), .Z(_02227__PTR170) );
  MUX2_X1 U4326 ( .A(1'b0), .B(_02392__PTR11), .S(_03169_), .Z(_02227__PTR171) );
  MUX2_X1 U4327 ( .A(1'b0), .B(_02392__PTR12), .S(_03169_), .Z(_02227__PTR172) );
  MUX2_X1 U4328 ( .A(1'b0), .B(_02392__PTR13), .S(_03169_), .Z(_02227__PTR173) );
  MUX2_X1 U4329 ( .A(1'b0), .B(_02392__PTR14), .S(_03169_), .Z(_02227__PTR174) );
  MUX2_X1 U4330 ( .A(1'b0), .B(_02392__PTR15), .S(_03169_), .Z(_02227__PTR175) );
  MUX2_X1 U4331 ( .A(1'b0), .B(_02392__PTR16), .S(_03169_), .Z(_02227__PTR176) );
  MUX2_X1 U4332 ( .A(1'b0), .B(_02392__PTR17), .S(_03169_), .Z(_02227__PTR177) );
  MUX2_X1 U4333 ( .A(1'b0), .B(_02392__PTR18), .S(_03169_), .Z(_02227__PTR178) );
  MUX2_X1 U4334 ( .A(1'b0), .B(_02392__PTR19), .S(_03169_), .Z(_02227__PTR179) );
  MUX2_X1 U4335 ( .A(1'b0), .B(_02392__PTR20), .S(_03169_), .Z(_02227__PTR180) );
  MUX2_X1 U4336 ( .A(1'b0), .B(_02392__PTR21), .S(_03169_), .Z(_02227__PTR181) );
  MUX2_X1 U4337 ( .A(1'b0), .B(_02392__PTR22), .S(_03169_), .Z(_02227__PTR182) );
  MUX2_X1 U4338 ( .A(1'b0), .B(_02392__PTR23), .S(_03169_), .Z(_02227__PTR183) );
  MUX2_X1 U4339 ( .A(1'b0), .B(_02392__PTR24), .S(_03169_), .Z(_02227__PTR184) );
  MUX2_X1 U4340 ( .A(1'b0), .B(_02392__PTR25), .S(_03169_), .Z(_02227__PTR185) );
  MUX2_X1 U4341 ( .A(1'b0), .B(_02392__PTR26), .S(_03169_), .Z(_02227__PTR186) );
  MUX2_X1 U4342 ( .A(1'b0), .B(_02392__PTR27), .S(_03169_), .Z(_02227__PTR187) );
  MUX2_X1 U4343 ( .A(1'b0), .B(_02392__PTR28), .S(_03169_), .Z(_02227__PTR188) );
  MUX2_X1 U4344 ( .A(1'b0), .B(_02392__PTR29), .S(_03169_), .Z(_02227__PTR189) );
  MUX2_X1 U4345 ( .A(1'b0), .B(_02392__PTR30), .S(_03169_), .Z(_02227__PTR190) );
  MUX2_X1 U4346 ( .A(1'b0), .B(_02392__PTR31), .S(_03169_), .Z(_02227__PTR191) );
  MUX2_X1 U4347 ( .A(1'b0), .B(_02388__PTR0), .S(_03168_), .Z(_02226__PTR160) );
  MUX2_X1 U4348 ( .A(1'b0), .B(_02388__PTR1), .S(_03168_), .Z(_02226__PTR161) );
  MUX2_X1 U4349 ( .A(1'b0), .B(_02388__PTR2), .S(_03168_), .Z(_02226__PTR162) );
  MUX2_X1 U4350 ( .A(1'b0), .B(_02388__PTR3), .S(_03168_), .Z(_02226__PTR163) );
  MUX2_X1 U4351 ( .A(1'b0), .B(_02388__PTR4), .S(_03168_), .Z(_02226__PTR164) );
  MUX2_X1 U4352 ( .A(1'b0), .B(_02388__PTR5), .S(_03168_), .Z(_02226__PTR165) );
  MUX2_X1 U4353 ( .A(1'b0), .B(_02388__PTR6), .S(_03168_), .Z(_02226__PTR166) );
  MUX2_X1 U4354 ( .A(1'b0), .B(_02388__PTR7), .S(_03168_), .Z(_02226__PTR167) );
  MUX2_X1 U4355 ( .A(1'b0), .B(_02388__PTR8), .S(_03168_), .Z(_02226__PTR168) );
  MUX2_X1 U4356 ( .A(1'b0), .B(_02388__PTR9), .S(_03168_), .Z(_02226__PTR169) );
  MUX2_X1 U4357 ( .A(1'b0), .B(_02388__PTR10), .S(_03168_), .Z(_02226__PTR170) );
  MUX2_X1 U4358 ( .A(1'b0), .B(_02388__PTR11), .S(_03168_), .Z(_02226__PTR171) );
  MUX2_X1 U4359 ( .A(1'b0), .B(_02388__PTR12), .S(_03168_), .Z(_02226__PTR172) );
  MUX2_X1 U4360 ( .A(1'b0), .B(_02388__PTR13), .S(_03168_), .Z(_02226__PTR173) );
  MUX2_X1 U4361 ( .A(1'b0), .B(_02388__PTR14), .S(_03168_), .Z(_02226__PTR174) );
  MUX2_X1 U4362 ( .A(1'b0), .B(_02388__PTR15), .S(_03168_), .Z(_02226__PTR175) );
  MUX2_X1 U4363 ( .A(1'b0), .B(_02388__PTR16), .S(_03168_), .Z(_02226__PTR176) );
  MUX2_X1 U4364 ( .A(1'b0), .B(_02388__PTR17), .S(_03168_), .Z(_02226__PTR177) );
  MUX2_X1 U4365 ( .A(1'b0), .B(_02388__PTR18), .S(_03168_), .Z(_02226__PTR178) );
  MUX2_X1 U4366 ( .A(1'b0), .B(_02388__PTR19), .S(_03168_), .Z(_02226__PTR179) );
  MUX2_X1 U4367 ( .A(1'b0), .B(_02388__PTR20), .S(_03168_), .Z(_02226__PTR180) );
  MUX2_X1 U4368 ( .A(1'b0), .B(_02388__PTR21), .S(_03168_), .Z(_02226__PTR181) );
  MUX2_X1 U4369 ( .A(1'b0), .B(_02388__PTR22), .S(_03168_), .Z(_02226__PTR182) );
  MUX2_X1 U4370 ( .A(1'b0), .B(_02388__PTR23), .S(_03168_), .Z(_02226__PTR183) );
  MUX2_X1 U4371 ( .A(1'b0), .B(_02388__PTR24), .S(_03168_), .Z(_02226__PTR184) );
  MUX2_X1 U4372 ( .A(1'b0), .B(_02388__PTR25), .S(_03168_), .Z(_02226__PTR185) );
  MUX2_X1 U4373 ( .A(1'b0), .B(_02388__PTR26), .S(_03168_), .Z(_02226__PTR186) );
  MUX2_X1 U4374 ( .A(1'b0), .B(_02388__PTR27), .S(_03168_), .Z(_02226__PTR187) );
  MUX2_X1 U4375 ( .A(1'b0), .B(_02388__PTR28), .S(_03168_), .Z(_02226__PTR188) );
  MUX2_X1 U4376 ( .A(1'b0), .B(_02388__PTR29), .S(_03168_), .Z(_02226__PTR189) );
  MUX2_X1 U4377 ( .A(1'b0), .B(_02388__PTR30), .S(_03168_), .Z(_02226__PTR190) );
  MUX2_X1 U4378 ( .A(1'b0), .B(_02388__PTR31), .S(_03168_), .Z(_02226__PTR191) );
  MUX2_X1 U4379 ( .A(1'b0), .B(_02153_), .S(_03018_), .Z(_02145__PTR5) );
  MUX2_X1 U4380 ( .A(1'b0), .B(_02149_), .S(_03017_), .Z(_02144__PTR5) );
  MUX2_X1 U4381 ( .A(1'b0), .B(_02380__PTR0), .S(_03166_), .Z(_02224__PTR40) );
  MUX2_X1 U4382 ( .A(1'b0), .B(_02380__PTR1), .S(_03166_), .Z(_02224__PTR41) );
  MUX2_X1 U4383 ( .A(1'b0), .B(_02380__PTR2), .S(_03166_), .Z(_02224__PTR42) );
  MUX2_X1 U4384 ( .A(1'b0), .B(_02380__PTR3), .S(_03166_), .Z(_02224__PTR43) );
  MUX2_X1 U4385 ( .A(1'b0), .B(_02380__PTR4), .S(_03166_), .Z(_02224__PTR44) );
  MUX2_X1 U4386 ( .A(1'b0), .B(_02168_), .S(_03021_), .Z(_02143__PTR5) );
  MUX2_X1 U4387 ( .A(1'b0), .B(_02157_), .S(_03019_), .Z(_02142__PTR5) );
  MUX2_X1 U4388 ( .A(1'b0), .B(_02164_), .S(_03021_), .Z(_02141__PTR5) );
  MUX2_X1 U4389 ( .A(1'b0), .B(_02160_), .S(_03020_), .Z(_02140__PTR5) );
  MUX2_X1 U4390 ( .A(1'b0), .B(_02395__PTR0), .S(_03170_), .Z(_02188__PTR320) );
  MUX2_X1 U4391 ( .A(1'b0), .B(_02395__PTR1), .S(_03170_), .Z(_02188__PTR321) );
  MUX2_X1 U4392 ( .A(1'b0), .B(_02395__PTR2), .S(_03170_), .Z(_02188__PTR322) );
  MUX2_X1 U4393 ( .A(1'b0), .B(_02395__PTR3), .S(_03170_), .Z(_02188__PTR323) );
  MUX2_X1 U4394 ( .A(1'b0), .B(_02395__PTR4), .S(_03170_), .Z(_02188__PTR324) );
  MUX2_X1 U4395 ( .A(1'b0), .B(_02395__PTR5), .S(_03170_), .Z(_02188__PTR325) );
  MUX2_X1 U4396 ( .A(1'b0), .B(_02395__PTR6), .S(_03170_), .Z(_02188__PTR326) );
  MUX2_X1 U4397 ( .A(1'b0), .B(_02395__PTR7), .S(_03170_), .Z(_02188__PTR327) );
  MUX2_X1 U4398 ( .A(1'b0), .B(_02395__PTR8), .S(_03170_), .Z(_02188__PTR328) );
  MUX2_X1 U4399 ( .A(1'b0), .B(_02395__PTR9), .S(_03170_), .Z(_02188__PTR329) );
  MUX2_X1 U4400 ( .A(1'b0), .B(_02395__PTR10), .S(_03170_), .Z(_02188__PTR330) );
  MUX2_X1 U4401 ( .A(1'b0), .B(_02395__PTR11), .S(_03170_), .Z(_02188__PTR331) );
  MUX2_X1 U4402 ( .A(1'b0), .B(_02395__PTR12), .S(_03170_), .Z(_02188__PTR332) );
  MUX2_X1 U4403 ( .A(1'b0), .B(_02395__PTR13), .S(_03170_), .Z(_02188__PTR333) );
  MUX2_X1 U4404 ( .A(1'b0), .B(_02395__PTR14), .S(_03170_), .Z(_02188__PTR334) );
  MUX2_X1 U4405 ( .A(1'b0), .B(_02395__PTR15), .S(_03170_), .Z(_02188__PTR335) );
  MUX2_X1 U4406 ( .A(1'b0), .B(_02395__PTR16), .S(_03170_), .Z(_02188__PTR336) );
  MUX2_X1 U4407 ( .A(1'b0), .B(_02395__PTR17), .S(_03170_), .Z(_02188__PTR337) );
  MUX2_X1 U4408 ( .A(1'b0), .B(_02395__PTR18), .S(_03170_), .Z(_02188__PTR338) );
  MUX2_X1 U4409 ( .A(1'b0), .B(_02395__PTR19), .S(_03170_), .Z(_02188__PTR339) );
  MUX2_X1 U4410 ( .A(1'b0), .B(_02395__PTR20), .S(_03170_), .Z(_02188__PTR340) );
  MUX2_X1 U4411 ( .A(1'b0), .B(_02395__PTR21), .S(_03170_), .Z(_02188__PTR341) );
  MUX2_X1 U4412 ( .A(1'b0), .B(_02395__PTR22), .S(_03170_), .Z(_02188__PTR342) );
  MUX2_X1 U4413 ( .A(1'b0), .B(_02395__PTR23), .S(_03170_), .Z(_02188__PTR343) );
  MUX2_X1 U4414 ( .A(1'b0), .B(_02395__PTR24), .S(_03170_), .Z(_02188__PTR344) );
  MUX2_X1 U4415 ( .A(1'b0), .B(_02395__PTR25), .S(_03170_), .Z(_02188__PTR345) );
  MUX2_X1 U4416 ( .A(1'b0), .B(_02395__PTR26), .S(_03170_), .Z(_02188__PTR346) );
  MUX2_X1 U4417 ( .A(1'b0), .B(_02395__PTR27), .S(_03170_), .Z(_02188__PTR347) );
  MUX2_X1 U4418 ( .A(1'b0), .B(_02395__PTR28), .S(_03170_), .Z(_02188__PTR348) );
  MUX2_X1 U4419 ( .A(1'b0), .B(_02395__PTR29), .S(_03170_), .Z(_02188__PTR349) );
  MUX2_X1 U4420 ( .A(1'b0), .B(_02395__PTR30), .S(_03170_), .Z(_02188__PTR350) );
  MUX2_X1 U4421 ( .A(1'b0), .B(_02395__PTR31), .S(_03170_), .Z(_02188__PTR352) );
  MUX2_X1 U4422 ( .A(1'b0), .B(_02376__PTR0), .S(_03165_), .Z(_02185__PTR160) );
  MUX2_X1 U4423 ( .A(1'b0), .B(_02376__PTR1), .S(_03165_), .Z(_02185__PTR161) );
  MUX2_X1 U4424 ( .A(1'b0), .B(_02376__PTR2), .S(_03165_), .Z(_02185__PTR162) );
  MUX2_X1 U4425 ( .A(1'b0), .B(_02376__PTR3), .S(_03165_), .Z(_02185__PTR163) );
  MUX2_X1 U4426 ( .A(1'b0), .B(_02376__PTR4), .S(_03165_), .Z(_02185__PTR164) );
  MUX2_X1 U4427 ( .A(1'b0), .B(_02376__PTR5), .S(_03165_), .Z(_02185__PTR165) );
  MUX2_X1 U4428 ( .A(1'b0), .B(_02376__PTR6), .S(_03165_), .Z(_02185__PTR166) );
  MUX2_X1 U4429 ( .A(1'b0), .B(_02376__PTR7), .S(_03165_), .Z(_02185__PTR167) );
  MUX2_X1 U4430 ( .A(1'b0), .B(_02376__PTR8), .S(_03165_), .Z(_02185__PTR168) );
  MUX2_X1 U4431 ( .A(1'b0), .B(_02376__PTR9), .S(_03165_), .Z(_02185__PTR169) );
  MUX2_X1 U4432 ( .A(1'b0), .B(_02376__PTR10), .S(_03165_), .Z(_02185__PTR170) );
  MUX2_X1 U4433 ( .A(1'b0), .B(_02376__PTR11), .S(_03165_), .Z(_02185__PTR171) );
  MUX2_X1 U4434 ( .A(1'b0), .B(_02376__PTR12), .S(_03165_), .Z(_02185__PTR172) );
  MUX2_X1 U4435 ( .A(1'b0), .B(_02376__PTR13), .S(_03165_), .Z(_02185__PTR173) );
  MUX2_X1 U4436 ( .A(1'b0), .B(_02376__PTR14), .S(_03165_), .Z(_02185__PTR174) );
  MUX2_X1 U4437 ( .A(1'b0), .B(_02376__PTR15), .S(_03165_), .Z(_02185__PTR175) );
  MUX2_X1 U4438 ( .A(1'b0), .B(_02376__PTR16), .S(_03165_), .Z(_02185__PTR176) );
  MUX2_X1 U4439 ( .A(1'b0), .B(_02376__PTR17), .S(_03165_), .Z(_02185__PTR177) );
  MUX2_X1 U4440 ( .A(1'b0), .B(_02376__PTR18), .S(_03165_), .Z(_02185__PTR178) );
  MUX2_X1 U4441 ( .A(1'b0), .B(_02376__PTR19), .S(_03165_), .Z(_02185__PTR179) );
  MUX2_X1 U4442 ( .A(1'b0), .B(_02376__PTR20), .S(_03165_), .Z(_02185__PTR180) );
  MUX2_X1 U4443 ( .A(1'b0), .B(_02376__PTR21), .S(_03165_), .Z(_02185__PTR181) );
  MUX2_X1 U4444 ( .A(1'b0), .B(_02376__PTR22), .S(_03165_), .Z(_02185__PTR182) );
  MUX2_X1 U4445 ( .A(1'b0), .B(_02376__PTR23), .S(_03165_), .Z(_02185__PTR183) );
  MUX2_X1 U4446 ( .A(1'b0), .B(_02376__PTR24), .S(_03165_), .Z(_02185__PTR184) );
  MUX2_X1 U4447 ( .A(1'b0), .B(_02376__PTR25), .S(_03165_), .Z(_02185__PTR185) );
  MUX2_X1 U4448 ( .A(1'b0), .B(_02376__PTR26), .S(_03165_), .Z(_02185__PTR186) );
  MUX2_X1 U4449 ( .A(1'b0), .B(_02376__PTR27), .S(_03165_), .Z(_02185__PTR187) );
  MUX2_X1 U4450 ( .A(1'b0), .B(_02376__PTR28), .S(_03165_), .Z(_02185__PTR188) );
  MUX2_X1 U4451 ( .A(1'b0), .B(_02376__PTR29), .S(_03165_), .Z(_02185__PTR189) );
  MUX2_X1 U4452 ( .A(1'b0), .B(_02376__PTR30), .S(_03165_), .Z(_02185__PTR190) );
  MUX2_X1 U4453 ( .A(1'b0), .B(_02376__PTR31), .S(_03165_), .Z(_02185__PTR191) );
  MUX2_X1 U4454 ( .A(1'b0), .B(_02384__PTR0), .S(_03167_), .Z(_02184__PTR160) );
  MUX2_X1 U4455 ( .A(1'b0), .B(_02384__PTR1), .S(_03167_), .Z(_02184__PTR161) );
  MUX2_X1 U4456 ( .A(1'b0), .B(_02384__PTR2), .S(_03167_), .Z(_02184__PTR162) );
  MUX2_X1 U4457 ( .A(1'b0), .B(_02384__PTR3), .S(_03167_), .Z(_02184__PTR163) );
  MUX2_X1 U4458 ( .A(1'b0), .B(_02384__PTR4), .S(_03167_), .Z(_02184__PTR164) );
  MUX2_X1 U4459 ( .A(1'b0), .B(_02384__PTR5), .S(_03167_), .Z(_02184__PTR165) );
  MUX2_X1 U4460 ( .A(1'b0), .B(_02384__PTR6), .S(_03167_), .Z(_02184__PTR166) );
  MUX2_X1 U4461 ( .A(1'b0), .B(_02384__PTR7), .S(_03167_), .Z(_02184__PTR167) );
  MUX2_X1 U4462 ( .A(1'b0), .B(_02384__PTR8), .S(_03167_), .Z(_02184__PTR168) );
  MUX2_X1 U4463 ( .A(1'b0), .B(_02384__PTR9), .S(_03167_), .Z(_02184__PTR169) );
  MUX2_X1 U4464 ( .A(1'b0), .B(_02384__PTR10), .S(_03167_), .Z(_02184__PTR170) );
  MUX2_X1 U4465 ( .A(1'b0), .B(_02384__PTR11), .S(_03167_), .Z(_02184__PTR171) );
  MUX2_X1 U4466 ( .A(1'b0), .B(_02384__PTR12), .S(_03167_), .Z(_02184__PTR172) );
  MUX2_X1 U4467 ( .A(1'b0), .B(_02384__PTR13), .S(_03167_), .Z(_02184__PTR173) );
  MUX2_X1 U4468 ( .A(1'b0), .B(_02384__PTR14), .S(_03167_), .Z(_02184__PTR174) );
  MUX2_X1 U4469 ( .A(1'b0), .B(_02384__PTR15), .S(_03167_), .Z(_02184__PTR175) );
  MUX2_X1 U4470 ( .A(1'b0), .B(_02384__PTR16), .S(_03167_), .Z(_02184__PTR176) );
  MUX2_X1 U4471 ( .A(1'b0), .B(_02384__PTR17), .S(_03167_), .Z(_02184__PTR177) );
  MUX2_X1 U4472 ( .A(1'b0), .B(_02384__PTR18), .S(_03167_), .Z(_02184__PTR178) );
  MUX2_X1 U4473 ( .A(1'b0), .B(_02384__PTR19), .S(_03167_), .Z(_02184__PTR179) );
  MUX2_X1 U4474 ( .A(1'b0), .B(_02384__PTR20), .S(_03167_), .Z(_02184__PTR180) );
  MUX2_X1 U4475 ( .A(1'b0), .B(_02384__PTR21), .S(_03167_), .Z(_02184__PTR181) );
  MUX2_X1 U4476 ( .A(1'b0), .B(_02384__PTR22), .S(_03167_), .Z(_02184__PTR182) );
  MUX2_X1 U4477 ( .A(1'b0), .B(_02384__PTR23), .S(_03167_), .Z(_02184__PTR183) );
  MUX2_X1 U4478 ( .A(1'b0), .B(_02384__PTR24), .S(_03167_), .Z(_02184__PTR184) );
  MUX2_X1 U4479 ( .A(1'b0), .B(_02384__PTR25), .S(_03167_), .Z(_02184__PTR185) );
  MUX2_X1 U4480 ( .A(1'b0), .B(_02384__PTR26), .S(_03167_), .Z(_02184__PTR186) );
  MUX2_X1 U4481 ( .A(1'b0), .B(_02384__PTR27), .S(_03167_), .Z(_02184__PTR187) );
  MUX2_X1 U4482 ( .A(1'b0), .B(_02384__PTR28), .S(_03167_), .Z(_02184__PTR188) );
  MUX2_X1 U4483 ( .A(1'b0), .B(_02384__PTR29), .S(_03167_), .Z(_02184__PTR189) );
  MUX2_X1 U4484 ( .A(1'b0), .B(_02384__PTR30), .S(_03167_), .Z(_02184__PTR190) );
  MUX2_X1 U4485 ( .A(1'b0), .B(_02384__PTR31), .S(_03167_), .Z(_02184__PTR191) );
  MUX2_X1 U4486 ( .A(1'b0), .B(_02411__PTR0), .S(_03173_), .Z(_02410__PTR0) );
  MUX2_X1 U4487 ( .A(1'b0), .B(_02411__PTR1), .S(_03173_), .Z(_02410__PTR1) );
  MUX2_X1 U4488 ( .A(1'b0), .B(_02411__PTR2), .S(_03173_), .Z(_02410__PTR2) );
  MUX2_X1 U4489 ( .A(1'b0), .B(_02411__PTR3), .S(_03173_), .Z(_02410__PTR3) );
  MUX2_X1 U4490 ( .A(1'b0), .B(_02704__PTR0), .S(_03419_), .Z(_02703__PTR0) );
  MUX2_X1 U4491 ( .A(1'b0), .B(_02704__PTR1), .S(_03419_), .Z(_02703__PTR1) );
  MUX2_X1 U4492 ( .A(1'b0), .B(_02704__PTR2), .S(_03419_), .Z(_02703__PTR2) );
  MUX2_X1 U4493 ( .A(1'b0), .B(_02704__PTR3), .S(_03419_), .Z(_02703__PTR3) );
  MUX2_X1 U4494 ( .A(1'b0), .B(_02695__PTR0), .S(_03417_), .Z(_02519__PTR320) );
  MUX2_X1 U4495 ( .A(1'b0), .B(_02695__PTR1), .S(_03417_), .Z(_02519__PTR321) );
  MUX2_X1 U4496 ( .A(1'b0), .B(_02695__PTR2), .S(_03417_), .Z(_02519__PTR322) );
  MUX2_X1 U4497 ( .A(1'b0), .B(_02695__PTR3), .S(_03417_), .Z(_02519__PTR323) );
  MUX2_X1 U4498 ( .A(1'b0), .B(_02695__PTR4), .S(_03417_), .Z(_02519__PTR324) );
  MUX2_X1 U4499 ( .A(1'b0), .B(_02695__PTR5), .S(_03417_), .Z(_02519__PTR325) );
  MUX2_X1 U4500 ( .A(1'b0), .B(_02695__PTR6), .S(_03417_), .Z(_02519__PTR326) );
  MUX2_X1 U4501 ( .A(1'b0), .B(_02695__PTR7), .S(_03417_), .Z(_02519__PTR327) );
  MUX2_X1 U4502 ( .A(1'b0), .B(_02695__PTR8), .S(_03417_), .Z(_02519__PTR328) );
  MUX2_X1 U4503 ( .A(1'b0), .B(_02695__PTR9), .S(_03417_), .Z(_02519__PTR329) );
  MUX2_X1 U4504 ( .A(1'b0), .B(_02695__PTR10), .S(_03417_), .Z(_02519__PTR330) );
  MUX2_X1 U4505 ( .A(1'b0), .B(_02695__PTR11), .S(_03417_), .Z(_02519__PTR331) );
  MUX2_X1 U4506 ( .A(1'b0), .B(_02695__PTR12), .S(_03417_), .Z(_02519__PTR332) );
  MUX2_X1 U4507 ( .A(1'b0), .B(_02695__PTR13), .S(_03417_), .Z(_02519__PTR333) );
  MUX2_X1 U4508 ( .A(1'b0), .B(_02695__PTR14), .S(_03417_), .Z(_02519__PTR334) );
  MUX2_X1 U4509 ( .A(1'b0), .B(_02695__PTR15), .S(_03417_), .Z(_02519__PTR335) );
  MUX2_X1 U4510 ( .A(1'b0), .B(_02695__PTR16), .S(_03417_), .Z(_02519__PTR336) );
  MUX2_X1 U4511 ( .A(1'b0), .B(_02695__PTR17), .S(_03417_), .Z(_02519__PTR337) );
  MUX2_X1 U4512 ( .A(1'b0), .B(_02695__PTR18), .S(_03417_), .Z(_02519__PTR338) );
  MUX2_X1 U4513 ( .A(1'b0), .B(_02695__PTR19), .S(_03417_), .Z(_02519__PTR339) );
  MUX2_X1 U4514 ( .A(1'b0), .B(_02695__PTR20), .S(_03417_), .Z(_02519__PTR340) );
  MUX2_X1 U4515 ( .A(1'b0), .B(_02695__PTR21), .S(_03417_), .Z(_02519__PTR341) );
  MUX2_X1 U4516 ( .A(1'b0), .B(_02695__PTR22), .S(_03417_), .Z(_02519__PTR342) );
  MUX2_X1 U4517 ( .A(1'b0), .B(_02695__PTR23), .S(_03417_), .Z(_02519__PTR343) );
  MUX2_X1 U4518 ( .A(1'b0), .B(_02695__PTR24), .S(_03417_), .Z(_02519__PTR344) );
  MUX2_X1 U4519 ( .A(1'b0), .B(_02695__PTR25), .S(_03417_), .Z(_02519__PTR345) );
  MUX2_X1 U4520 ( .A(1'b0), .B(_02695__PTR26), .S(_03417_), .Z(_02519__PTR346) );
  MUX2_X1 U4521 ( .A(1'b0), .B(_02695__PTR27), .S(_03417_), .Z(_02519__PTR347) );
  MUX2_X1 U4522 ( .A(1'b0), .B(_02695__PTR28), .S(_03417_), .Z(_02519__PTR348) );
  MUX2_X1 U4523 ( .A(1'b0), .B(_02695__PTR29), .S(_03417_), .Z(_02519__PTR349) );
  MUX2_X1 U4524 ( .A(1'b0), .B(_02695__PTR30), .S(_03417_), .Z(_02519__PTR350) );
  MUX2_X1 U4525 ( .A(1'b0), .B(_02695__PTR31), .S(_03417_), .Z(_02519__PTR352) );
  MUX2_X1 U4526 ( .A(1'b0), .B(_02691__PTR0), .S(_03416_), .Z(_02518__PTR80) );
  MUX2_X1 U4527 ( .A(1'b0), .B(_02691__PTR1), .S(_03416_), .Z(_02518__PTR81) );
  MUX2_X1 U4528 ( .A(1'b0), .B(_02691__PTR2), .S(_03416_), .Z(_02518__PTR82) );
  MUX2_X1 U4529 ( .A(1'b0), .B(_02691__PTR3), .S(_03416_), .Z(_02518__PTR83) );
  MUX2_X1 U4530 ( .A(1'b0), .B(_02691__PTR4), .S(_03416_), .Z(_02518__PTR84) );
  MUX2_X1 U4531 ( .A(1'b0), .B(_02691__PTR5), .S(_03416_), .Z(_02518__PTR85) );
  MUX2_X1 U4532 ( .A(1'b0), .B(_02691__PTR6), .S(_03416_), .Z(_02518__PTR86) );
  MUX2_X1 U4533 ( .A(1'b0), .B(_02691__PTR7), .S(_03416_), .Z(_02518__PTR87) );
  MUX2_X1 U4534 ( .A(1'b0), .B(_02691__PTR8), .S(_03416_), .Z(_02518__PTR88) );
  MUX2_X1 U4535 ( .A(1'b0), .B(_02691__PTR9), .S(_03416_), .Z(_02518__PTR89) );
  MUX2_X1 U4536 ( .A(1'b0), .B(_02691__PTR10), .S(_03416_), .Z(_02518__PTR90) );
  MUX2_X1 U4537 ( .A(1'b0), .B(_02691__PTR11), .S(_03416_), .Z(_02518__PTR91) );
  MUX2_X1 U4538 ( .A(1'b0), .B(_02691__PTR12), .S(_03416_), .Z(_02518__PTR92) );
  MUX2_X1 U4539 ( .A(1'b0), .B(_02691__PTR13), .S(_03416_), .Z(_02518__PTR93) );
  MUX2_X1 U4540 ( .A(1'b0), .B(_02691__PTR14), .S(_03416_), .Z(_02518__PTR94) );
  MUX2_X1 U4541 ( .A(1'b0), .B(_02691__PTR15), .S(_03416_), .Z(_02518__PTR95) );
  MUX2_X1 U4542 ( .A(1'b0), .B(_02688__PTR0), .S(_03416_), .Z(_02517__PTR80) );
  MUX2_X1 U4543 ( .A(1'b0), .B(_02688__PTR1), .S(_03416_), .Z(_02517__PTR81) );
  MUX2_X1 U4544 ( .A(1'b0), .B(_02688__PTR2), .S(_03416_), .Z(_02517__PTR82) );
  MUX2_X1 U4545 ( .A(1'b0), .B(_02688__PTR3), .S(_03416_), .Z(_02517__PTR83) );
  MUX2_X1 U4546 ( .A(1'b0), .B(_02688__PTR4), .S(_03416_), .Z(_02517__PTR84) );
  MUX2_X1 U4547 ( .A(1'b0), .B(_02688__PTR5), .S(_03416_), .Z(_02517__PTR85) );
  MUX2_X1 U4548 ( .A(1'b0), .B(_02688__PTR6), .S(_03416_), .Z(_02517__PTR86) );
  MUX2_X1 U4549 ( .A(1'b0), .B(_02688__PTR7), .S(_03416_), .Z(_02517__PTR87) );
  MUX2_X1 U4550 ( .A(1'b0), .B(_02688__PTR8), .S(_03416_), .Z(_02517__PTR88) );
  MUX2_X1 U4551 ( .A(1'b0), .B(_02688__PTR9), .S(_03416_), .Z(_02517__PTR89) );
  MUX2_X1 U4552 ( .A(1'b0), .B(_02688__PTR10), .S(_03416_), .Z(_02517__PTR90) );
  MUX2_X1 U4553 ( .A(1'b0), .B(_02688__PTR11), .S(_03416_), .Z(_02517__PTR91) );
  MUX2_X1 U4554 ( .A(1'b0), .B(_02688__PTR12), .S(_03416_), .Z(_02517__PTR92) );
  MUX2_X1 U4555 ( .A(1'b0), .B(_02688__PTR13), .S(_03416_), .Z(_02517__PTR93) );
  MUX2_X1 U4556 ( .A(1'b0), .B(_02688__PTR14), .S(_03416_), .Z(_02517__PTR94) );
  MUX2_X1 U4557 ( .A(1'b0), .B(_02681__PTR0), .S(_03414_), .Z(_02516__PTR160) );
  MUX2_X1 U4558 ( .A(1'b0), .B(_02681__PTR1), .S(_03414_), .Z(_02516__PTR161) );
  MUX2_X1 U4559 ( .A(1'b0), .B(_02681__PTR2), .S(_03414_), .Z(_02516__PTR162) );
  MUX2_X1 U4560 ( .A(1'b0), .B(_02681__PTR3), .S(_03414_), .Z(_02516__PTR163) );
  MUX2_X1 U4561 ( .A(1'b0), .B(_02681__PTR4), .S(_03414_), .Z(_02516__PTR164) );
  MUX2_X1 U4562 ( .A(1'b0), .B(_02681__PTR5), .S(_03414_), .Z(_02516__PTR165) );
  MUX2_X1 U4563 ( .A(1'b0), .B(_02681__PTR6), .S(_03414_), .Z(_02516__PTR166) );
  MUX2_X1 U4564 ( .A(1'b0), .B(_02681__PTR7), .S(_03414_), .Z(_02516__PTR167) );
  MUX2_X1 U4565 ( .A(1'b0), .B(_02681__PTR8), .S(_03414_), .Z(_02516__PTR168) );
  MUX2_X1 U4566 ( .A(1'b0), .B(_02681__PTR9), .S(_03414_), .Z(_02516__PTR169) );
  MUX2_X1 U4567 ( .A(1'b0), .B(_02681__PTR10), .S(_03414_), .Z(_02516__PTR170) );
  MUX2_X1 U4568 ( .A(1'b0), .B(_02681__PTR11), .S(_03414_), .Z(_02516__PTR171) );
  MUX2_X1 U4569 ( .A(1'b0), .B(_02681__PTR12), .S(_03414_), .Z(_02516__PTR172) );
  MUX2_X1 U4570 ( .A(1'b0), .B(_02681__PTR13), .S(_03414_), .Z(_02516__PTR173) );
  MUX2_X1 U4571 ( .A(1'b0), .B(_02681__PTR14), .S(_03414_), .Z(_02516__PTR174) );
  MUX2_X1 U4572 ( .A(1'b0), .B(_02681__PTR15), .S(_03414_), .Z(_02516__PTR175) );
  MUX2_X1 U4573 ( .A(1'b0), .B(_02681__PTR16), .S(_03414_), .Z(_02516__PTR176) );
  MUX2_X1 U4574 ( .A(1'b0), .B(_02681__PTR17), .S(_03414_), .Z(_02516__PTR177) );
  MUX2_X1 U4575 ( .A(1'b0), .B(_02681__PTR18), .S(_03414_), .Z(_02516__PTR178) );
  MUX2_X1 U4576 ( .A(1'b0), .B(_02681__PTR19), .S(_03414_), .Z(_02516__PTR179) );
  MUX2_X1 U4577 ( .A(1'b0), .B(_02681__PTR20), .S(_03414_), .Z(_02516__PTR180) );
  MUX2_X1 U4578 ( .A(1'b0), .B(_02681__PTR21), .S(_03414_), .Z(_02516__PTR181) );
  MUX2_X1 U4579 ( .A(1'b0), .B(_02681__PTR22), .S(_03414_), .Z(_02516__PTR182) );
  MUX2_X1 U4580 ( .A(1'b0), .B(_02681__PTR23), .S(_03414_), .Z(_02516__PTR183) );
  MUX2_X1 U4581 ( .A(1'b0), .B(_02681__PTR24), .S(_03414_), .Z(_02516__PTR184) );
  MUX2_X1 U4582 ( .A(1'b0), .B(_02681__PTR25), .S(_03414_), .Z(_02516__PTR185) );
  MUX2_X1 U4583 ( .A(1'b0), .B(_02681__PTR26), .S(_03414_), .Z(_02516__PTR186) );
  MUX2_X1 U4584 ( .A(1'b0), .B(_02681__PTR27), .S(_03414_), .Z(_02516__PTR187) );
  MUX2_X1 U4585 ( .A(1'b0), .B(_02681__PTR28), .S(_03414_), .Z(_02516__PTR188) );
  MUX2_X1 U4586 ( .A(1'b0), .B(_02681__PTR29), .S(_03414_), .Z(_02516__PTR189) );
  MUX2_X1 U4587 ( .A(1'b0), .B(_02681__PTR30), .S(_03414_), .Z(_02516__PTR190) );
  MUX2_X1 U4588 ( .A(1'b0), .B(_02681__PTR31), .S(_03414_), .Z(_02516__PTR191) );
  MUX2_X1 U4589 ( .A(1'b0), .B(_02677__PTR0), .S(_03413_), .Z(_02515__PTR160) );
  MUX2_X1 U4590 ( .A(1'b0), .B(_02677__PTR1), .S(_03413_), .Z(_02515__PTR161) );
  MUX2_X1 U4591 ( .A(1'b0), .B(_02677__PTR2), .S(_03413_), .Z(_02515__PTR162) );
  MUX2_X1 U4592 ( .A(1'b0), .B(_02677__PTR3), .S(_03413_), .Z(_02515__PTR163) );
  MUX2_X1 U4593 ( .A(1'b0), .B(_02677__PTR4), .S(_03413_), .Z(_02515__PTR164) );
  MUX2_X1 U4594 ( .A(1'b0), .B(_02677__PTR5), .S(_03413_), .Z(_02515__PTR165) );
  MUX2_X1 U4595 ( .A(1'b0), .B(_02677__PTR6), .S(_03413_), .Z(_02515__PTR166) );
  MUX2_X1 U4596 ( .A(1'b0), .B(_02677__PTR7), .S(_03413_), .Z(_02515__PTR167) );
  MUX2_X1 U4597 ( .A(1'b0), .B(_02677__PTR8), .S(_03413_), .Z(_02515__PTR168) );
  MUX2_X1 U4598 ( .A(1'b0), .B(_02677__PTR9), .S(_03413_), .Z(_02515__PTR169) );
  MUX2_X1 U4599 ( .A(1'b0), .B(_02677__PTR10), .S(_03413_), .Z(_02515__PTR170) );
  MUX2_X1 U4600 ( .A(1'b0), .B(_02677__PTR11), .S(_03413_), .Z(_02515__PTR171) );
  MUX2_X1 U4601 ( .A(1'b0), .B(_02677__PTR12), .S(_03413_), .Z(_02515__PTR172) );
  MUX2_X1 U4602 ( .A(1'b0), .B(_02677__PTR13), .S(_03413_), .Z(_02515__PTR173) );
  MUX2_X1 U4603 ( .A(1'b0), .B(_02677__PTR14), .S(_03413_), .Z(_02515__PTR174) );
  MUX2_X1 U4604 ( .A(1'b0), .B(_02677__PTR15), .S(_03413_), .Z(_02515__PTR175) );
  MUX2_X1 U4605 ( .A(1'b0), .B(_02677__PTR16), .S(_03413_), .Z(_02515__PTR176) );
  MUX2_X1 U4606 ( .A(1'b0), .B(_02677__PTR17), .S(_03413_), .Z(_02515__PTR177) );
  MUX2_X1 U4607 ( .A(1'b0), .B(_02677__PTR18), .S(_03413_), .Z(_02515__PTR178) );
  MUX2_X1 U4608 ( .A(1'b0), .B(_02677__PTR19), .S(_03413_), .Z(_02515__PTR179) );
  MUX2_X1 U4609 ( .A(1'b0), .B(_02677__PTR20), .S(_03413_), .Z(_02515__PTR180) );
  MUX2_X1 U4610 ( .A(1'b0), .B(_02677__PTR21), .S(_03413_), .Z(_02515__PTR181) );
  MUX2_X1 U4611 ( .A(1'b0), .B(_02677__PTR22), .S(_03413_), .Z(_02515__PTR182) );
  MUX2_X1 U4612 ( .A(1'b0), .B(_02677__PTR23), .S(_03413_), .Z(_02515__PTR183) );
  MUX2_X1 U4613 ( .A(1'b0), .B(_02677__PTR24), .S(_03413_), .Z(_02515__PTR184) );
  MUX2_X1 U4614 ( .A(1'b0), .B(_02677__PTR25), .S(_03413_), .Z(_02515__PTR185) );
  MUX2_X1 U4615 ( .A(1'b0), .B(_02677__PTR26), .S(_03413_), .Z(_02515__PTR186) );
  MUX2_X1 U4616 ( .A(1'b0), .B(_02677__PTR27), .S(_03413_), .Z(_02515__PTR187) );
  MUX2_X1 U4617 ( .A(1'b0), .B(_02677__PTR28), .S(_03413_), .Z(_02515__PTR188) );
  MUX2_X1 U4618 ( .A(1'b0), .B(_02677__PTR29), .S(_03413_), .Z(_02515__PTR189) );
  MUX2_X1 U4619 ( .A(1'b0), .B(_02677__PTR30), .S(_03413_), .Z(_02515__PTR190) );
  MUX2_X1 U4620 ( .A(1'b0), .B(_02677__PTR31), .S(_03413_), .Z(_02515__PTR191) );
  MUX2_X1 U4621 ( .A(1'b0), .B(_02442_), .S(_03263_), .Z(_02434__PTR5) );
  MUX2_X1 U4622 ( .A(1'b0), .B(_02438_), .S(_03262_), .Z(_02433__PTR5) );
  MUX2_X1 U4623 ( .A(1'b0), .B(_02669__PTR0), .S(_03411_), .Z(_02513__PTR40) );
  MUX2_X1 U4624 ( .A(1'b0), .B(_02669__PTR1), .S(_03411_), .Z(_02513__PTR41) );
  MUX2_X1 U4625 ( .A(1'b0), .B(_02669__PTR2), .S(_03411_), .Z(_02513__PTR42) );
  MUX2_X1 U4626 ( .A(1'b0), .B(_02669__PTR3), .S(_03411_), .Z(_02513__PTR43) );
  MUX2_X1 U4627 ( .A(1'b0), .B(_02669__PTR4), .S(_03411_), .Z(_02513__PTR44) );
  MUX2_X1 U4628 ( .A(1'b0), .B(_02457_), .S(_03266_), .Z(_02432__PTR5) );
  MUX2_X1 U4629 ( .A(1'b0), .B(_02446_), .S(_03264_), .Z(_02431__PTR5) );
  MUX2_X1 U4630 ( .A(1'b0), .B(_02453_), .S(_03266_), .Z(_02430__PTR5) );
  MUX2_X1 U4631 ( .A(1'b0), .B(_02449_), .S(_03265_), .Z(_02429__PTR5) );
  MUX2_X1 U4632 ( .A(1'b0), .B(_02684__PTR0), .S(_03415_), .Z(_02477__PTR320) );
  MUX2_X1 U4633 ( .A(1'b0), .B(_02684__PTR1), .S(_03415_), .Z(_02477__PTR321) );
  MUX2_X1 U4634 ( .A(1'b0), .B(_02684__PTR2), .S(_03415_), .Z(_02477__PTR322) );
  MUX2_X1 U4635 ( .A(1'b0), .B(_02684__PTR3), .S(_03415_), .Z(_02477__PTR323) );
  MUX2_X1 U4636 ( .A(1'b0), .B(_02684__PTR4), .S(_03415_), .Z(_02477__PTR324) );
  MUX2_X1 U4637 ( .A(1'b0), .B(_02684__PTR5), .S(_03415_), .Z(_02477__PTR325) );
  MUX2_X1 U4638 ( .A(1'b0), .B(_02684__PTR6), .S(_03415_), .Z(_02477__PTR326) );
  MUX2_X1 U4639 ( .A(1'b0), .B(_02684__PTR7), .S(_03415_), .Z(_02477__PTR327) );
  MUX2_X1 U4640 ( .A(1'b0), .B(_02684__PTR8), .S(_03415_), .Z(_02477__PTR328) );
  MUX2_X1 U4641 ( .A(1'b0), .B(_02684__PTR9), .S(_03415_), .Z(_02477__PTR329) );
  MUX2_X1 U4642 ( .A(1'b0), .B(_02684__PTR10), .S(_03415_), .Z(_02477__PTR330) );
  MUX2_X1 U4643 ( .A(1'b0), .B(_02684__PTR11), .S(_03415_), .Z(_02477__PTR331) );
  MUX2_X1 U4644 ( .A(1'b0), .B(_02684__PTR12), .S(_03415_), .Z(_02477__PTR332) );
  MUX2_X1 U4645 ( .A(1'b0), .B(_02684__PTR13), .S(_03415_), .Z(_02477__PTR333) );
  MUX2_X1 U4646 ( .A(1'b0), .B(_02684__PTR14), .S(_03415_), .Z(_02477__PTR334) );
  MUX2_X1 U4647 ( .A(1'b0), .B(_02684__PTR15), .S(_03415_), .Z(_02477__PTR335) );
  MUX2_X1 U4648 ( .A(1'b0), .B(_02684__PTR16), .S(_03415_), .Z(_02477__PTR336) );
  MUX2_X1 U4649 ( .A(1'b0), .B(_02684__PTR17), .S(_03415_), .Z(_02477__PTR337) );
  MUX2_X1 U4650 ( .A(1'b0), .B(_02684__PTR18), .S(_03415_), .Z(_02477__PTR338) );
  MUX2_X1 U4651 ( .A(1'b0), .B(_02684__PTR19), .S(_03415_), .Z(_02477__PTR339) );
  MUX2_X1 U4652 ( .A(1'b0), .B(_02684__PTR20), .S(_03415_), .Z(_02477__PTR340) );
  MUX2_X1 U4653 ( .A(1'b0), .B(_02684__PTR21), .S(_03415_), .Z(_02477__PTR341) );
  MUX2_X1 U4654 ( .A(1'b0), .B(_02684__PTR22), .S(_03415_), .Z(_02477__PTR342) );
  MUX2_X1 U4655 ( .A(1'b0), .B(_02684__PTR23), .S(_03415_), .Z(_02477__PTR343) );
  MUX2_X1 U4656 ( .A(1'b0), .B(_02684__PTR24), .S(_03415_), .Z(_02477__PTR344) );
  MUX2_X1 U4657 ( .A(1'b0), .B(_02684__PTR25), .S(_03415_), .Z(_02477__PTR345) );
  MUX2_X1 U4658 ( .A(1'b0), .B(_02684__PTR26), .S(_03415_), .Z(_02477__PTR346) );
  MUX2_X1 U4659 ( .A(1'b0), .B(_02684__PTR27), .S(_03415_), .Z(_02477__PTR347) );
  MUX2_X1 U4660 ( .A(1'b0), .B(_02684__PTR28), .S(_03415_), .Z(_02477__PTR348) );
  MUX2_X1 U4661 ( .A(1'b0), .B(_02684__PTR29), .S(_03415_), .Z(_02477__PTR349) );
  MUX2_X1 U4662 ( .A(1'b0), .B(_02684__PTR30), .S(_03415_), .Z(_02477__PTR350) );
  MUX2_X1 U4663 ( .A(1'b0), .B(_02684__PTR31), .S(_03415_), .Z(_02477__PTR352) );
  MUX2_X1 U4664 ( .A(1'b0), .B(_02665__PTR0), .S(_03410_), .Z(_02474__PTR160) );
  MUX2_X1 U4665 ( .A(1'b0), .B(_02665__PTR1), .S(_03410_), .Z(_02474__PTR161) );
  MUX2_X1 U4666 ( .A(1'b0), .B(_02665__PTR2), .S(_03410_), .Z(_02474__PTR162) );
  MUX2_X1 U4667 ( .A(1'b0), .B(_02665__PTR3), .S(_03410_), .Z(_02474__PTR163) );
  MUX2_X1 U4668 ( .A(1'b0), .B(_02665__PTR4), .S(_03410_), .Z(_02474__PTR164) );
  MUX2_X1 U4669 ( .A(1'b0), .B(_02665__PTR5), .S(_03410_), .Z(_02474__PTR165) );
  MUX2_X1 U4670 ( .A(1'b0), .B(_02665__PTR6), .S(_03410_), .Z(_02474__PTR166) );
  MUX2_X1 U4671 ( .A(1'b0), .B(_02665__PTR7), .S(_03410_), .Z(_02474__PTR167) );
  MUX2_X1 U4672 ( .A(1'b0), .B(_02665__PTR8), .S(_03410_), .Z(_02474__PTR168) );
  MUX2_X1 U4673 ( .A(1'b0), .B(_02665__PTR9), .S(_03410_), .Z(_02474__PTR169) );
  MUX2_X1 U4674 ( .A(1'b0), .B(_02665__PTR10), .S(_03410_), .Z(_02474__PTR170) );
  MUX2_X1 U4675 ( .A(1'b0), .B(_02665__PTR11), .S(_03410_), .Z(_02474__PTR171) );
  MUX2_X1 U4676 ( .A(1'b0), .B(_02665__PTR12), .S(_03410_), .Z(_02474__PTR172) );
  MUX2_X1 U4677 ( .A(1'b0), .B(_02665__PTR13), .S(_03410_), .Z(_02474__PTR173) );
  MUX2_X1 U4678 ( .A(1'b0), .B(_02665__PTR14), .S(_03410_), .Z(_02474__PTR174) );
  MUX2_X1 U4679 ( .A(1'b0), .B(_02665__PTR15), .S(_03410_), .Z(_02474__PTR175) );
  MUX2_X1 U4680 ( .A(1'b0), .B(_02665__PTR16), .S(_03410_), .Z(_02474__PTR176) );
  MUX2_X1 U4681 ( .A(1'b0), .B(_02665__PTR17), .S(_03410_), .Z(_02474__PTR177) );
  MUX2_X1 U4682 ( .A(1'b0), .B(_02665__PTR18), .S(_03410_), .Z(_02474__PTR178) );
  MUX2_X1 U4683 ( .A(1'b0), .B(_02665__PTR19), .S(_03410_), .Z(_02474__PTR179) );
  MUX2_X1 U4684 ( .A(1'b0), .B(_02665__PTR20), .S(_03410_), .Z(_02474__PTR180) );
  MUX2_X1 U4685 ( .A(1'b0), .B(_02665__PTR21), .S(_03410_), .Z(_02474__PTR181) );
  MUX2_X1 U4686 ( .A(1'b0), .B(_02665__PTR22), .S(_03410_), .Z(_02474__PTR182) );
  MUX2_X1 U4687 ( .A(1'b0), .B(_02665__PTR23), .S(_03410_), .Z(_02474__PTR183) );
  MUX2_X1 U4688 ( .A(1'b0), .B(_02665__PTR24), .S(_03410_), .Z(_02474__PTR184) );
  MUX2_X1 U4689 ( .A(1'b0), .B(_02665__PTR25), .S(_03410_), .Z(_02474__PTR185) );
  MUX2_X1 U4690 ( .A(1'b0), .B(_02665__PTR26), .S(_03410_), .Z(_02474__PTR186) );
  MUX2_X1 U4691 ( .A(1'b0), .B(_02665__PTR27), .S(_03410_), .Z(_02474__PTR187) );
  MUX2_X1 U4692 ( .A(1'b0), .B(_02665__PTR28), .S(_03410_), .Z(_02474__PTR188) );
  MUX2_X1 U4693 ( .A(1'b0), .B(_02665__PTR29), .S(_03410_), .Z(_02474__PTR189) );
  MUX2_X1 U4694 ( .A(1'b0), .B(_02665__PTR30), .S(_03410_), .Z(_02474__PTR190) );
  MUX2_X1 U4695 ( .A(1'b0), .B(_02665__PTR31), .S(_03410_), .Z(_02474__PTR191) );
  MUX2_X1 U4696 ( .A(1'b0), .B(_02673__PTR0), .S(_03412_), .Z(_02473__PTR160) );
  MUX2_X1 U4697 ( .A(1'b0), .B(_02673__PTR1), .S(_03412_), .Z(_02473__PTR161) );
  MUX2_X1 U4698 ( .A(1'b0), .B(_02673__PTR2), .S(_03412_), .Z(_02473__PTR162) );
  MUX2_X1 U4699 ( .A(1'b0), .B(_02673__PTR3), .S(_03412_), .Z(_02473__PTR163) );
  MUX2_X1 U4700 ( .A(1'b0), .B(_02673__PTR4), .S(_03412_), .Z(_02473__PTR164) );
  MUX2_X1 U4701 ( .A(1'b0), .B(_02673__PTR5), .S(_03412_), .Z(_02473__PTR165) );
  MUX2_X1 U4702 ( .A(1'b0), .B(_02673__PTR6), .S(_03412_), .Z(_02473__PTR166) );
  MUX2_X1 U4703 ( .A(1'b0), .B(_02673__PTR7), .S(_03412_), .Z(_02473__PTR167) );
  MUX2_X1 U4704 ( .A(1'b0), .B(_02673__PTR8), .S(_03412_), .Z(_02473__PTR168) );
  MUX2_X1 U4705 ( .A(1'b0), .B(_02673__PTR9), .S(_03412_), .Z(_02473__PTR169) );
  MUX2_X1 U4706 ( .A(1'b0), .B(_02673__PTR10), .S(_03412_), .Z(_02473__PTR170) );
  MUX2_X1 U4707 ( .A(1'b0), .B(_02673__PTR11), .S(_03412_), .Z(_02473__PTR171) );
  MUX2_X1 U4708 ( .A(1'b0), .B(_02673__PTR12), .S(_03412_), .Z(_02473__PTR172) );
  MUX2_X1 U4709 ( .A(1'b0), .B(_02673__PTR13), .S(_03412_), .Z(_02473__PTR173) );
  MUX2_X1 U4710 ( .A(1'b0), .B(_02673__PTR14), .S(_03412_), .Z(_02473__PTR174) );
  MUX2_X1 U4711 ( .A(1'b0), .B(_02673__PTR15), .S(_03412_), .Z(_02473__PTR175) );
  MUX2_X1 U4712 ( .A(1'b0), .B(_02673__PTR16), .S(_03412_), .Z(_02473__PTR176) );
  MUX2_X1 U4713 ( .A(1'b0), .B(_02673__PTR17), .S(_03412_), .Z(_02473__PTR177) );
  MUX2_X1 U4714 ( .A(1'b0), .B(_02673__PTR18), .S(_03412_), .Z(_02473__PTR178) );
  MUX2_X1 U4715 ( .A(1'b0), .B(_02673__PTR19), .S(_03412_), .Z(_02473__PTR179) );
  MUX2_X1 U4716 ( .A(1'b0), .B(_02673__PTR20), .S(_03412_), .Z(_02473__PTR180) );
  MUX2_X1 U4717 ( .A(1'b0), .B(_02673__PTR21), .S(_03412_), .Z(_02473__PTR181) );
  MUX2_X1 U4718 ( .A(1'b0), .B(_02673__PTR22), .S(_03412_), .Z(_02473__PTR182) );
  MUX2_X1 U4719 ( .A(1'b0), .B(_02673__PTR23), .S(_03412_), .Z(_02473__PTR183) );
  MUX2_X1 U4720 ( .A(1'b0), .B(_02673__PTR24), .S(_03412_), .Z(_02473__PTR184) );
  MUX2_X1 U4721 ( .A(1'b0), .B(_02673__PTR25), .S(_03412_), .Z(_02473__PTR185) );
  MUX2_X1 U4722 ( .A(1'b0), .B(_02673__PTR26), .S(_03412_), .Z(_02473__PTR186) );
  MUX2_X1 U4723 ( .A(1'b0), .B(_02673__PTR27), .S(_03412_), .Z(_02473__PTR187) );
  MUX2_X1 U4724 ( .A(1'b0), .B(_02673__PTR28), .S(_03412_), .Z(_02473__PTR188) );
  MUX2_X1 U4725 ( .A(1'b0), .B(_02673__PTR29), .S(_03412_), .Z(_02473__PTR189) );
  MUX2_X1 U4726 ( .A(1'b0), .B(_02673__PTR30), .S(_03412_), .Z(_02473__PTR190) );
  MUX2_X1 U4727 ( .A(1'b0), .B(_02673__PTR31), .S(_03412_), .Z(_02473__PTR191) );
  MUX2_X1 U4728 ( .A(1'b0), .B(_02700__PTR0), .S(_03418_), .Z(_02699__PTR0) );
  MUX2_X1 U4729 ( .A(1'b0), .B(_02700__PTR1), .S(_03418_), .Z(_02699__PTR1) );
  MUX2_X1 U4730 ( .A(1'b0), .B(_02700__PTR2), .S(_03418_), .Z(_02699__PTR2) );
  MUX2_X1 U4731 ( .A(1'b0), .B(_02700__PTR3), .S(_03418_), .Z(_02699__PTR3) );
  MUX2_X1 U4732 ( .A(1'b0), .B(P2_Datao_PTR0), .S(_05770_), .Z(_05732__PTR0) );
  MUX2_X1 U4733 ( .A(1'b0), .B(P2_Datao_PTR1), .S(_05770_), .Z(_05732__PTR1) );
  MUX2_X1 U4734 ( .A(1'b0), .B(P2_Datao_PTR2), .S(_05770_), .Z(_05732__PTR2) );
  MUX2_X1 U4735 ( .A(1'b0), .B(P2_Datao_PTR3), .S(_05770_), .Z(_05732__PTR3) );
  MUX2_X1 U4736 ( .A(1'b0), .B(P2_Datao_PTR4), .S(_05770_), .Z(_05732__PTR4) );
  MUX2_X1 U4737 ( .A(1'b0), .B(P2_Datao_PTR5), .S(_05770_), .Z(_05732__PTR5) );
  MUX2_X1 U4738 ( .A(1'b0), .B(P2_Datao_PTR6), .S(_05770_), .Z(_05732__PTR6) );
  MUX2_X1 U4739 ( .A(1'b0), .B(P2_Datao_PTR7), .S(_05770_), .Z(_05732__PTR7) );
  MUX2_X1 U4740 ( .A(1'b0), .B(P2_Datao_PTR8), .S(_05770_), .Z(_05732__PTR8) );
  MUX2_X1 U4741 ( .A(1'b0), .B(P2_Datao_PTR9), .S(_05770_), .Z(_05732__PTR9) );
  MUX2_X1 U4742 ( .A(1'b0), .B(P2_Datao_PTR10), .S(_05770_), .Z(_05732__PTR10) );
  MUX2_X1 U4743 ( .A(1'b0), .B(P2_Datao_PTR11), .S(_05770_), .Z(_05732__PTR11) );
  MUX2_X1 U4744 ( .A(1'b0), .B(P2_Datao_PTR12), .S(_05770_), .Z(_05732__PTR12) );
  MUX2_X1 U4745 ( .A(1'b0), .B(P2_Datao_PTR13), .S(_05770_), .Z(_05732__PTR13) );
  MUX2_X1 U4746 ( .A(1'b0), .B(P2_Datao_PTR14), .S(_05770_), .Z(_05732__PTR14) );
  MUX2_X1 U4747 ( .A(1'b0), .B(P2_Datao_PTR15), .S(_05770_), .Z(_05732__PTR15) );
  MUX2_X1 U4748 ( .A(1'b0), .B(P2_Datao_PTR16), .S(_05770_), .Z(_05732__PTR16) );
  MUX2_X1 U4749 ( .A(1'b0), .B(P2_Datao_PTR17), .S(_05770_), .Z(_05732__PTR17) );
  MUX2_X1 U4750 ( .A(1'b0), .B(P2_Datao_PTR18), .S(_05770_), .Z(_05732__PTR18) );
  MUX2_X1 U4751 ( .A(1'b0), .B(P2_Datao_PTR19), .S(_05770_), .Z(_05732__PTR19) );
  MUX2_X1 U4752 ( .A(1'b0), .B(P2_Datao_PTR20), .S(_05770_), .Z(_05732__PTR20) );
  MUX2_X1 U4753 ( .A(1'b0), .B(P2_Datao_PTR21), .S(_05770_), .Z(_05732__PTR21) );
  MUX2_X1 U4754 ( .A(1'b0), .B(P2_Datao_PTR22), .S(_05770_), .Z(_05732__PTR22) );
  MUX2_X1 U4755 ( .A(1'b0), .B(P2_Datao_PTR23), .S(_05770_), .Z(_05732__PTR23) );
  MUX2_X1 U4756 ( .A(1'b0), .B(P2_Datao_PTR24), .S(_05770_), .Z(_05732__PTR24) );
  MUX2_X1 U4757 ( .A(1'b0), .B(P2_Datao_PTR25), .S(_05770_), .Z(_05732__PTR25) );
  MUX2_X1 U4758 ( .A(1'b0), .B(P2_Datao_PTR26), .S(_05770_), .Z(_05732__PTR26) );
  MUX2_X1 U4759 ( .A(1'b0), .B(P2_Datao_PTR27), .S(_05770_), .Z(_05732__PTR27) );
  MUX2_X1 U4760 ( .A(1'b0), .B(P2_Datao_PTR28), .S(_05770_), .Z(_05732__PTR28) );
  MUX2_X1 U4761 ( .A(1'b0), .B(P2_Datao_PTR29), .S(_05770_), .Z(_05732__PTR29) );
  MUX2_X1 U4762 ( .A(1'b0), .B(P2_Datao_PTR30), .S(_05770_), .Z(_05732__PTR30) );
  MUX2_X1 U4763 ( .A(1'b0), .B(P2_Datao_PTR31), .S(_05770_), .Z(_05732__PTR31) );
  MUX2_X1 U4764 ( .A(_05732__PTR0), .B(P1_Datao_PTR0), .S(_05760_), .Z(_05733__PTR0) );
  MUX2_X1 U4765 ( .A(_05732__PTR1), .B(P1_Datao_PTR1), .S(_05760_), .Z(_05733__PTR1) );
  MUX2_X1 U4766 ( .A(_05732__PTR2), .B(P1_Datao_PTR2), .S(_05760_), .Z(_05733__PTR2) );
  MUX2_X1 U4767 ( .A(_05732__PTR3), .B(P1_Datao_PTR3), .S(_05760_), .Z(_05733__PTR3) );
  MUX2_X1 U4768 ( .A(_05732__PTR4), .B(P1_Datao_PTR4), .S(_05760_), .Z(_05733__PTR4) );
  MUX2_X1 U4769 ( .A(_05732__PTR5), .B(P1_Datao_PTR5), .S(_05760_), .Z(_05733__PTR5) );
  MUX2_X1 U4770 ( .A(_05732__PTR6), .B(P1_Datao_PTR6), .S(_05760_), .Z(_05733__PTR6) );
  MUX2_X1 U4771 ( .A(_05732__PTR7), .B(P1_Datao_PTR7), .S(_05760_), .Z(_05733__PTR7) );
  MUX2_X1 U4772 ( .A(_05732__PTR8), .B(P1_Datao_PTR8), .S(_05760_), .Z(_05733__PTR8) );
  MUX2_X1 U4773 ( .A(_05732__PTR9), .B(P1_Datao_PTR9), .S(_05760_), .Z(_05733__PTR9) );
  MUX2_X1 U4774 ( .A(_05732__PTR10), .B(P1_Datao_PTR10), .S(_05760_), .Z(_05733__PTR10) );
  MUX2_X1 U4775 ( .A(_05732__PTR11), .B(P1_Datao_PTR11), .S(_05760_), .Z(_05733__PTR11) );
  MUX2_X1 U4776 ( .A(_05732__PTR12), .B(P1_Datao_PTR12), .S(_05760_), .Z(_05733__PTR12) );
  MUX2_X1 U4777 ( .A(_05732__PTR13), .B(P1_Datao_PTR13), .S(_05760_), .Z(_05733__PTR13) );
  MUX2_X1 U4778 ( .A(_05732__PTR14), .B(P1_Datao_PTR14), .S(_05760_), .Z(_05733__PTR14) );
  MUX2_X1 U4779 ( .A(_05732__PTR15), .B(P1_Datao_PTR15), .S(_05760_), .Z(_05733__PTR15) );
  MUX2_X1 U4780 ( .A(_05732__PTR16), .B(P1_Datao_PTR16), .S(_05760_), .Z(_05733__PTR16) );
  MUX2_X1 U4781 ( .A(_05732__PTR17), .B(P1_Datao_PTR17), .S(_05760_), .Z(_05733__PTR17) );
  MUX2_X1 U4782 ( .A(_05732__PTR18), .B(P1_Datao_PTR18), .S(_05760_), .Z(_05733__PTR18) );
  MUX2_X1 U4783 ( .A(_05732__PTR19), .B(P1_Datao_PTR19), .S(_05760_), .Z(_05733__PTR19) );
  MUX2_X1 U4784 ( .A(_05732__PTR20), .B(P1_Datao_PTR20), .S(_05760_), .Z(_05733__PTR20) );
  MUX2_X1 U4785 ( .A(_05732__PTR21), .B(P1_Datao_PTR21), .S(_05760_), .Z(_05733__PTR21) );
  MUX2_X1 U4786 ( .A(_05732__PTR22), .B(P1_Datao_PTR22), .S(_05760_), .Z(_05733__PTR22) );
  MUX2_X1 U4787 ( .A(_05732__PTR23), .B(P1_Datao_PTR23), .S(_05760_), .Z(_05733__PTR23) );
  MUX2_X1 U4788 ( .A(_05732__PTR24), .B(P1_Datao_PTR24), .S(_05760_), .Z(_05733__PTR24) );
  MUX2_X1 U4789 ( .A(_05732__PTR25), .B(P1_Datao_PTR25), .S(_05760_), .Z(_05733__PTR25) );
  MUX2_X1 U4790 ( .A(_05732__PTR26), .B(P1_Datao_PTR26), .S(_05760_), .Z(_05733__PTR26) );
  MUX2_X1 U4791 ( .A(_05732__PTR27), .B(P1_Datao_PTR27), .S(_05760_), .Z(_05733__PTR27) );
  MUX2_X1 U4792 ( .A(_05732__PTR28), .B(P1_Datao_PTR28), .S(_05760_), .Z(_05733__PTR28) );
  MUX2_X1 U4793 ( .A(_05732__PTR29), .B(P1_Datao_PTR29), .S(_05760_), .Z(_05733__PTR29) );
  MUX2_X1 U4794 ( .A(_05732__PTR30), .B(P1_Datao_PTR30), .S(_05760_), .Z(_05733__PTR30) );
  MUX2_X1 U4795 ( .A(_05732__PTR31), .B(P1_Datao_PTR31), .S(_05760_), .Z(_05733__PTR31) );
  INV_X1 U4796 ( .A(_05760_), .ZN(_05734_) );
  INV_X1 U4797 ( .A(_05770_), .ZN(_05735_) );
  MUX2_X1 U4798 ( .A(_05735_), .B(1'b1), .S(_05760_), .Z(_05736_) );
  INV_X1 U4799 ( .A(_05741_), .ZN(_05750_) );
  INV_X1 U4800 ( .A(_05749_), .ZN(_05751_) );
  MUX2_X1 U4801 ( .A(_05751_), .B(1'b1), .S(_05741_), .Z(_05752_) );
  MUX2_X1 U4802 ( .A(buf1_PTR0), .B(datai_PTR0), .S(_05718__PTR29), .Z(di1_PTR0) );
  MUX2_X1 U4803 ( .A(buf1_PTR1), .B(datai_PTR1), .S(_05718__PTR29), .Z(di1_PTR1) );
  MUX2_X1 U4804 ( .A(buf1_PTR2), .B(datai_PTR2), .S(_05718__PTR29), .Z(di1_PTR2) );
  MUX2_X1 U4805 ( .A(buf1_PTR3), .B(datai_PTR3), .S(_05718__PTR29), .Z(di1_PTR3) );
  MUX2_X1 U4806 ( .A(buf1_PTR4), .B(datai_PTR4), .S(_05718__PTR29), .Z(di1_PTR4) );
  MUX2_X1 U4807 ( .A(buf1_PTR5), .B(datai_PTR5), .S(_05718__PTR29), .Z(di1_PTR5) );
  MUX2_X1 U4808 ( .A(buf1_PTR6), .B(datai_PTR6), .S(_05718__PTR29), .Z(di1_PTR6) );
  MUX2_X1 U4809 ( .A(buf1_PTR7), .B(datai_PTR7), .S(_05718__PTR29), .Z(di1_PTR7) );
  MUX2_X1 U4810 ( .A(buf1_PTR8), .B(datai_PTR8), .S(_05718__PTR29), .Z(di1_PTR8) );
  MUX2_X1 U4811 ( .A(buf1_PTR9), .B(datai_PTR9), .S(_05718__PTR29), .Z(di1_PTR9) );
  MUX2_X1 U4812 ( .A(buf1_PTR10), .B(datai_PTR10), .S(_05718__PTR29), .Z(di1_PTR10) );
  MUX2_X1 U4813 ( .A(buf1_PTR11), .B(datai_PTR11), .S(_05718__PTR29), .Z(di1_PTR11) );
  MUX2_X1 U4814 ( .A(buf1_PTR12), .B(datai_PTR12), .S(_05718__PTR29), .Z(di1_PTR12) );
  MUX2_X1 U4815 ( .A(buf1_PTR13), .B(datai_PTR13), .S(_05718__PTR29), .Z(di1_PTR13) );
  MUX2_X1 U4816 ( .A(buf1_PTR14), .B(datai_PTR14), .S(_05718__PTR29), .Z(di1_PTR14) );
  MUX2_X1 U4817 ( .A(buf1_PTR15), .B(datai_PTR15), .S(_05718__PTR29), .Z(di1_PTR15) );
  MUX2_X1 U4818 ( .A(buf1_PTR16), .B(datai_PTR16), .S(_05718__PTR29), .Z(di1_PTR16) );
  MUX2_X1 U4819 ( .A(buf1_PTR17), .B(datai_PTR17), .S(_05718__PTR29), .Z(di1_PTR17) );
  MUX2_X1 U4820 ( .A(buf1_PTR18), .B(datai_PTR18), .S(_05718__PTR29), .Z(di1_PTR18) );
  MUX2_X1 U4821 ( .A(buf1_PTR19), .B(datai_PTR19), .S(_05718__PTR29), .Z(di1_PTR19) );
  MUX2_X1 U4822 ( .A(buf1_PTR20), .B(datai_PTR20), .S(_05718__PTR29), .Z(di1_PTR20) );
  MUX2_X1 U4823 ( .A(buf1_PTR21), .B(datai_PTR21), .S(_05718__PTR29), .Z(di1_PTR21) );
  MUX2_X1 U4824 ( .A(buf1_PTR22), .B(datai_PTR22), .S(_05718__PTR29), .Z(di1_PTR22) );
  MUX2_X1 U4825 ( .A(buf1_PTR23), .B(datai_PTR23), .S(_05718__PTR29), .Z(di1_PTR23) );
  MUX2_X1 U4826 ( .A(buf1_PTR24), .B(datai_PTR24), .S(_05718__PTR29), .Z(di1_PTR24) );
  MUX2_X1 U4827 ( .A(buf1_PTR25), .B(datai_PTR25), .S(_05718__PTR29), .Z(di1_PTR25) );
  MUX2_X1 U4828 ( .A(buf1_PTR26), .B(datai_PTR26), .S(_05718__PTR29), .Z(di1_PTR26) );
  MUX2_X1 U4829 ( .A(buf1_PTR27), .B(datai_PTR27), .S(_05718__PTR29), .Z(di1_PTR27) );
  MUX2_X1 U4830 ( .A(buf1_PTR28), .B(datai_PTR28), .S(_05718__PTR29), .Z(di1_PTR28) );
  MUX2_X1 U4831 ( .A(buf1_PTR29), .B(datai_PTR29), .S(_05718__PTR29), .Z(di1_PTR29) );
  MUX2_X1 U4832 ( .A(buf1_PTR30), .B(datai_PTR30), .S(_05718__PTR29), .Z(di1_PTR30) );
  MUX2_X1 U4833 ( .A(buf1_PTR31), .B(datai_PTR31), .S(_05718__PTR29), .Z(P1_Datai_PTR31) );
  MUX2_X1 U4834 ( .A(buf1_PTR0), .B(buf2_PTR0), .S(_05713__PTR29), .Z(di2_PTR0) );
  MUX2_X1 U4835 ( .A(buf1_PTR1), .B(buf2_PTR1), .S(_05713__PTR29), .Z(di2_PTR1) );
  MUX2_X1 U4836 ( .A(buf1_PTR2), .B(buf2_PTR2), .S(_05713__PTR29), .Z(di2_PTR2) );
  MUX2_X1 U4837 ( .A(buf1_PTR3), .B(buf2_PTR3), .S(_05713__PTR29), .Z(di2_PTR3) );
  MUX2_X1 U4838 ( .A(buf1_PTR4), .B(buf2_PTR4), .S(_05713__PTR29), .Z(di2_PTR4) );
  MUX2_X1 U4839 ( .A(buf1_PTR5), .B(buf2_PTR5), .S(_05713__PTR29), .Z(di2_PTR5) );
  MUX2_X1 U4840 ( .A(buf1_PTR6), .B(buf2_PTR6), .S(_05713__PTR29), .Z(di2_PTR6) );
  MUX2_X1 U4841 ( .A(buf1_PTR7), .B(buf2_PTR7), .S(_05713__PTR29), .Z(di2_PTR7) );
  MUX2_X1 U4842 ( .A(buf1_PTR8), .B(buf2_PTR8), .S(_05713__PTR29), .Z(di2_PTR8) );
  MUX2_X1 U4843 ( .A(buf1_PTR9), .B(buf2_PTR9), .S(_05713__PTR29), .Z(di2_PTR9) );
  MUX2_X1 U4844 ( .A(buf1_PTR10), .B(buf2_PTR10), .S(_05713__PTR29), .Z(di2_PTR10) );
  MUX2_X1 U4845 ( .A(buf1_PTR11), .B(buf2_PTR11), .S(_05713__PTR29), .Z(di2_PTR11) );
  MUX2_X1 U4846 ( .A(buf1_PTR12), .B(buf2_PTR12), .S(_05713__PTR29), .Z(di2_PTR12) );
  MUX2_X1 U4847 ( .A(buf1_PTR13), .B(buf2_PTR13), .S(_05713__PTR29), .Z(di2_PTR13) );
  MUX2_X1 U4848 ( .A(buf1_PTR14), .B(buf2_PTR14), .S(_05713__PTR29), .Z(di2_PTR14) );
  MUX2_X1 U4849 ( .A(buf1_PTR15), .B(buf2_PTR15), .S(_05713__PTR29), .Z(di2_PTR15) );
  MUX2_X1 U4850 ( .A(buf1_PTR16), .B(buf2_PTR16), .S(_05713__PTR29), .Z(di2_PTR16) );
  MUX2_X1 U4851 ( .A(buf1_PTR17), .B(buf2_PTR17), .S(_05713__PTR29), .Z(di2_PTR17) );
  MUX2_X1 U4852 ( .A(buf1_PTR18), .B(buf2_PTR18), .S(_05713__PTR29), .Z(di2_PTR18) );
  MUX2_X1 U4853 ( .A(buf1_PTR19), .B(buf2_PTR19), .S(_05713__PTR29), .Z(di2_PTR19) );
  MUX2_X1 U4854 ( .A(buf1_PTR20), .B(buf2_PTR20), .S(_05713__PTR29), .Z(di2_PTR20) );
  MUX2_X1 U4855 ( .A(buf1_PTR21), .B(buf2_PTR21), .S(_05713__PTR29), .Z(di2_PTR21) );
  MUX2_X1 U4856 ( .A(buf1_PTR22), .B(buf2_PTR22), .S(_05713__PTR29), .Z(di2_PTR22) );
  MUX2_X1 U4857 ( .A(buf1_PTR23), .B(buf2_PTR23), .S(_05713__PTR29), .Z(di2_PTR23) );
  MUX2_X1 U4858 ( .A(buf1_PTR24), .B(buf2_PTR24), .S(_05713__PTR29), .Z(di2_PTR24) );
  MUX2_X1 U4859 ( .A(buf1_PTR25), .B(buf2_PTR25), .S(_05713__PTR29), .Z(di2_PTR25) );
  MUX2_X1 U4860 ( .A(buf1_PTR26), .B(buf2_PTR26), .S(_05713__PTR29), .Z(di2_PTR26) );
  MUX2_X1 U4861 ( .A(buf1_PTR27), .B(buf2_PTR27), .S(_05713__PTR29), .Z(di2_PTR27) );
  MUX2_X1 U4862 ( .A(buf1_PTR28), .B(buf2_PTR28), .S(_05713__PTR29), .Z(di2_PTR28) );
  MUX2_X1 U4863 ( .A(buf1_PTR29), .B(buf2_PTR29), .S(_05713__PTR29), .Z(di2_PTR29) );
  MUX2_X1 U4864 ( .A(buf1_PTR30), .B(buf2_PTR30), .S(_05713__PTR29), .Z(di2_PTR30) );
  MUX2_X1 U4865 ( .A(buf1_PTR31), .B(buf2_PTR31), .S(_05713__PTR29), .Z(P2_Datai_PTR31) );
  MUX2_X1 U4866 ( .A(P2_Address_PTR0), .B(P3_Address_PTR0), .S(_05762_), .Z(address2_PTR0) );
  MUX2_X1 U4867 ( .A(P2_Address_PTR1), .B(P3_Address_PTR1), .S(_05762_), .Z(address2_PTR1) );
  MUX2_X1 U4868 ( .A(P2_Address_PTR2), .B(P3_Address_PTR2), .S(_05762_), .Z(address2_PTR2) );
  MUX2_X1 U4869 ( .A(P2_Address_PTR3), .B(P3_Address_PTR3), .S(_05762_), .Z(address2_PTR3) );
  MUX2_X1 U4870 ( .A(P2_Address_PTR4), .B(P3_Address_PTR4), .S(_05762_), .Z(address2_PTR4) );
  MUX2_X1 U4871 ( .A(P2_Address_PTR5), .B(P3_Address_PTR5), .S(_05762_), .Z(address2_PTR5) );
  MUX2_X1 U4872 ( .A(P2_Address_PTR6), .B(P3_Address_PTR6), .S(_05762_), .Z(address2_PTR6) );
  MUX2_X1 U4873 ( .A(P2_Address_PTR7), .B(P3_Address_PTR7), .S(_05762_), .Z(address2_PTR7) );
  MUX2_X1 U4874 ( .A(P2_Address_PTR8), .B(P3_Address_PTR8), .S(_05762_), .Z(address2_PTR8) );
  MUX2_X1 U4875 ( .A(P2_Address_PTR9), .B(P3_Address_PTR9), .S(_05762_), .Z(address2_PTR9) );
  MUX2_X1 U4876 ( .A(P2_Address_PTR10), .B(P3_Address_PTR10), .S(_05762_), .Z(address2_PTR10) );
  MUX2_X1 U4877 ( .A(P2_Address_PTR11), .B(P3_Address_PTR11), .S(_05762_), .Z(address2_PTR11) );
  MUX2_X1 U4878 ( .A(P2_Address_PTR12), .B(P3_Address_PTR12), .S(_05762_), .Z(address2_PTR12) );
  MUX2_X1 U4879 ( .A(P2_Address_PTR13), .B(P3_Address_PTR13), .S(_05762_), .Z(address2_PTR13) );
  MUX2_X1 U4880 ( .A(P2_Address_PTR14), .B(P3_Address_PTR14), .S(_05762_), .Z(address2_PTR14) );
  MUX2_X1 U4881 ( .A(P2_Address_PTR15), .B(P3_Address_PTR15), .S(_05762_), .Z(address2_PTR15) );
  MUX2_X1 U4882 ( .A(P2_Address_PTR16), .B(P3_Address_PTR16), .S(_05762_), .Z(address2_PTR16) );
  MUX2_X1 U4883 ( .A(P2_Address_PTR17), .B(P3_Address_PTR17), .S(_05762_), .Z(address2_PTR17) );
  MUX2_X1 U4884 ( .A(P2_Address_PTR18), .B(P3_Address_PTR18), .S(_05762_), .Z(address2_PTR18) );
  MUX2_X1 U4885 ( .A(P2_Address_PTR19), .B(P3_Address_PTR19), .S(_05762_), .Z(address2_PTR19) );
  MUX2_X1 U4886 ( .A(P2_Address_PTR20), .B(P3_Address_PTR20), .S(_05762_), .Z(address2_PTR20) );
  MUX2_X1 U4887 ( .A(P2_Address_PTR21), .B(P3_Address_PTR21), .S(_05762_), .Z(address2_PTR21) );
  MUX2_X1 U4888 ( .A(P2_Address_PTR22), .B(P3_Address_PTR22), .S(_05762_), .Z(address2_PTR22) );
  MUX2_X1 U4889 ( .A(P2_Address_PTR23), .B(P3_Address_PTR23), .S(_05762_), .Z(address2_PTR23) );
  MUX2_X1 U4890 ( .A(P2_Address_PTR24), .B(P3_Address_PTR24), .S(_05762_), .Z(address2_PTR24) );
  MUX2_X1 U4891 ( .A(P2_Address_PTR25), .B(P3_Address_PTR25), .S(_05762_), .Z(address2_PTR25) );
  MUX2_X1 U4892 ( .A(P2_Address_PTR26), .B(P3_Address_PTR26), .S(_05762_), .Z(address2_PTR26) );
  MUX2_X1 U4893 ( .A(P2_Address_PTR27), .B(P3_Address_PTR27), .S(_05762_), .Z(address2_PTR27) );
  MUX2_X1 U4894 ( .A(P2_Address_PTR28), .B(P3_Address_PTR28), .S(_05762_), .Z(address2_PTR28) );
  MUX2_X1 U4895 ( .A(P2_Address_PTR29), .B(P3_Address_PTR29), .S(_05762_), .Z(address2_PTR29) );
  MUX2_X1 U4896 ( .A(1'b0), .B(_01836__PTR0), .S(_01770__PTR2), .Z(_01930__PTR64) );
  MUX2_X1 U4897 ( .A(1'b0), .B(_01836__PTR1), .S(_01770__PTR2), .Z(_01930__PTR65) );
  MUX2_X1 U4898 ( .A(1'b0), .B(_01836__PTR2), .S(_01770__PTR2), .Z(_01930__PTR66) );
  MUX2_X1 U4899 ( .A(1'b0), .B(_01836__PTR3), .S(_01770__PTR2), .Z(_01930__PTR67) );
  MUX2_X1 U4900 ( .A(1'b0), .B(1'b0), .S(_01770__PTR2), .Z(_01930__PTR68) );
  MUX2_X1 U4901 ( .A(1'b0), .B(_01884__PTR3), .S(_01770__PTR2), .Z(_01932__PTR64) );
  MUX2_X1 U4902 ( .A(1'b0), .B(_01884__PTR4), .S(_01770__PTR2), .Z(_01932__PTR65) );
  MUX2_X1 U4903 ( .A(1'b0), .B(_01884__PTR5), .S(_01770__PTR2), .Z(_01932__PTR66) );
  MUX2_X1 U4904 ( .A(1'b0), .B(_01884__PTR6), .S(_01770__PTR2), .Z(_01932__PTR67) );
  MUX2_X1 U4905 ( .A(1'b0), .B(_02082__PTR0), .S(_01770__PTR2), .Z(_01928__PTR64) );
  MUX2_X1 U4906 ( .A(1'b0), .B(_02082__PTR1), .S(_01770__PTR2), .Z(_01928__PTR65) );
  MUX2_X1 U4907 ( .A(1'b0), .B(_02082__PTR2), .S(_01770__PTR2), .Z(_01928__PTR66) );
  MUX2_X1 U4908 ( .A(1'b0), .B(_02082__PTR3), .S(_01770__PTR2), .Z(_01928__PTR67) );
  MUX2_X1 U4909 ( .A(1'b0), .B(_02082__PTR4), .S(_01770__PTR2), .Z(_01928__PTR68) );
  MUX2_X1 U4910 ( .A(1'b0), .B(_02082__PTR5), .S(_01770__PTR2), .Z(_01928__PTR69) );
  MUX2_X1 U4911 ( .A(1'b0), .B(_02082__PTR6), .S(_01770__PTR2), .Z(_01928__PTR70) );
  MUX2_X1 U4912 ( .A(1'b0), .B(_02082__PTR7), .S(_01770__PTR2), .Z(_01928__PTR71) );
  MUX2_X1 U4913 ( .A(1'b0), .B(_02081__PTR0), .S(_01770__PTR2), .Z(_01926__PTR64) );
  MUX2_X1 U4914 ( .A(1'b0), .B(_02081__PTR1), .S(_01770__PTR2), .Z(_01926__PTR65) );
  MUX2_X1 U4915 ( .A(1'b0), .B(_02081__PTR2), .S(_01770__PTR2), .Z(_01926__PTR66) );
  MUX2_X1 U4916 ( .A(1'b0), .B(_02081__PTR3), .S(_01770__PTR2), .Z(_01926__PTR67) );
  MUX2_X1 U4917 ( .A(1'b0), .B(_02081__PTR4), .S(_01770__PTR2), .Z(_01926__PTR68) );
  MUX2_X1 U4918 ( .A(1'b0), .B(_02081__PTR5), .S(_01770__PTR2), .Z(_01926__PTR69) );
  MUX2_X1 U4919 ( .A(1'b0), .B(_02081__PTR6), .S(_01770__PTR2), .Z(_01926__PTR70) );
  MUX2_X1 U4920 ( .A(1'b0), .B(_02081__PTR7), .S(_01770__PTR2), .Z(_01926__PTR71) );
  MUX2_X1 U4921 ( .A(1'b0), .B(_02080__PTR0), .S(_01770__PTR2), .Z(_01924__PTR64) );
  MUX2_X1 U4922 ( .A(1'b0), .B(_02080__PTR1), .S(_01770__PTR2), .Z(_01924__PTR65) );
  MUX2_X1 U4923 ( .A(1'b0), .B(_02080__PTR2), .S(_01770__PTR2), .Z(_01924__PTR66) );
  MUX2_X1 U4924 ( .A(1'b0), .B(_02080__PTR3), .S(_01770__PTR2), .Z(_01924__PTR67) );
  MUX2_X1 U4925 ( .A(1'b0), .B(_02080__PTR4), .S(_01770__PTR2), .Z(_01924__PTR68) );
  MUX2_X1 U4926 ( .A(1'b0), .B(_02080__PTR5), .S(_01770__PTR2), .Z(_01924__PTR69) );
  MUX2_X1 U4927 ( .A(1'b0), .B(_02080__PTR6), .S(_01770__PTR2), .Z(_01924__PTR70) );
  MUX2_X1 U4928 ( .A(1'b0), .B(_02080__PTR7), .S(_01770__PTR2), .Z(_01924__PTR71) );
  MUX2_X1 U4929 ( .A(1'b0), .B(_02079__PTR0), .S(_01770__PTR2), .Z(_01922__PTR64) );
  MUX2_X1 U4930 ( .A(1'b0), .B(_02079__PTR1), .S(_01770__PTR2), .Z(_01922__PTR65) );
  MUX2_X1 U4931 ( .A(1'b0), .B(_02079__PTR2), .S(_01770__PTR2), .Z(_01922__PTR66) );
  MUX2_X1 U4932 ( .A(1'b0), .B(_02079__PTR3), .S(_01770__PTR2), .Z(_01922__PTR67) );
  MUX2_X1 U4933 ( .A(1'b0), .B(_02079__PTR4), .S(_01770__PTR2), .Z(_01922__PTR68) );
  MUX2_X1 U4934 ( .A(1'b0), .B(_02079__PTR5), .S(_01770__PTR2), .Z(_01922__PTR69) );
  MUX2_X1 U4935 ( .A(1'b0), .B(_02079__PTR6), .S(_01770__PTR2), .Z(_01922__PTR70) );
  MUX2_X1 U4936 ( .A(1'b0), .B(_02079__PTR7), .S(_01770__PTR2), .Z(_01922__PTR71) );
  MUX2_X1 U4937 ( .A(1'b0), .B(_02078__PTR0), .S(_01770__PTR2), .Z(_01920__PTR64) );
  MUX2_X1 U4938 ( .A(1'b0), .B(_02078__PTR1), .S(_01770__PTR2), .Z(_01920__PTR65) );
  MUX2_X1 U4939 ( .A(1'b0), .B(_02078__PTR2), .S(_01770__PTR2), .Z(_01920__PTR66) );
  MUX2_X1 U4940 ( .A(1'b0), .B(_02078__PTR3), .S(_01770__PTR2), .Z(_01920__PTR67) );
  MUX2_X1 U4941 ( .A(1'b0), .B(_02078__PTR4), .S(_01770__PTR2), .Z(_01920__PTR68) );
  MUX2_X1 U4942 ( .A(1'b0), .B(_02078__PTR5), .S(_01770__PTR2), .Z(_01920__PTR69) );
  MUX2_X1 U4943 ( .A(1'b0), .B(_02078__PTR6), .S(_01770__PTR2), .Z(_01920__PTR70) );
  MUX2_X1 U4944 ( .A(1'b0), .B(_02078__PTR7), .S(_01770__PTR2), .Z(_01920__PTR71) );
  MUX2_X1 U4945 ( .A(1'b0), .B(_02077__PTR0), .S(_01770__PTR2), .Z(_01918__PTR64) );
  MUX2_X1 U4946 ( .A(1'b0), .B(_02077__PTR1), .S(_01770__PTR2), .Z(_01918__PTR65) );
  MUX2_X1 U4947 ( .A(1'b0), .B(_02077__PTR2), .S(_01770__PTR2), .Z(_01918__PTR66) );
  MUX2_X1 U4948 ( .A(1'b0), .B(_02077__PTR3), .S(_01770__PTR2), .Z(_01918__PTR67) );
  MUX2_X1 U4949 ( .A(1'b0), .B(_02077__PTR4), .S(_01770__PTR2), .Z(_01918__PTR68) );
  MUX2_X1 U4950 ( .A(1'b0), .B(_02077__PTR5), .S(_01770__PTR2), .Z(_01918__PTR69) );
  MUX2_X1 U4951 ( .A(1'b0), .B(_02077__PTR6), .S(_01770__PTR2), .Z(_01918__PTR70) );
  MUX2_X1 U4952 ( .A(1'b0), .B(_02077__PTR7), .S(_01770__PTR2), .Z(_01918__PTR71) );
  MUX2_X1 U4953 ( .A(1'b0), .B(_02076__PTR0), .S(_01770__PTR2), .Z(_01916__PTR64) );
  MUX2_X1 U4954 ( .A(1'b0), .B(_02076__PTR1), .S(_01770__PTR2), .Z(_01916__PTR65) );
  MUX2_X1 U4955 ( .A(1'b0), .B(_02076__PTR2), .S(_01770__PTR2), .Z(_01916__PTR66) );
  MUX2_X1 U4956 ( .A(1'b0), .B(_02076__PTR3), .S(_01770__PTR2), .Z(_01916__PTR67) );
  MUX2_X1 U4957 ( .A(1'b0), .B(_02076__PTR4), .S(_01770__PTR2), .Z(_01916__PTR68) );
  MUX2_X1 U4958 ( .A(1'b0), .B(_02076__PTR5), .S(_01770__PTR2), .Z(_01916__PTR69) );
  MUX2_X1 U4959 ( .A(1'b0), .B(_02076__PTR6), .S(_01770__PTR2), .Z(_01916__PTR70) );
  MUX2_X1 U4960 ( .A(1'b0), .B(_02076__PTR7), .S(_01770__PTR2), .Z(_01916__PTR71) );
  MUX2_X1 U4961 ( .A(1'b0), .B(_02075__PTR0), .S(_01770__PTR2), .Z(_01914__PTR64) );
  MUX2_X1 U4962 ( .A(1'b0), .B(_02075__PTR1), .S(_01770__PTR2), .Z(_01914__PTR65) );
  MUX2_X1 U4963 ( .A(1'b0), .B(_02075__PTR2), .S(_01770__PTR2), .Z(_01914__PTR66) );
  MUX2_X1 U4964 ( .A(1'b0), .B(_02075__PTR3), .S(_01770__PTR2), .Z(_01914__PTR67) );
  MUX2_X1 U4965 ( .A(1'b0), .B(_02075__PTR4), .S(_01770__PTR2), .Z(_01914__PTR68) );
  MUX2_X1 U4966 ( .A(1'b0), .B(_02075__PTR5), .S(_01770__PTR2), .Z(_01914__PTR69) );
  MUX2_X1 U4967 ( .A(1'b0), .B(_02075__PTR6), .S(_01770__PTR2), .Z(_01914__PTR70) );
  MUX2_X1 U4968 ( .A(1'b0), .B(_02075__PTR7), .S(_01770__PTR2), .Z(_01914__PTR71) );
  MUX2_X1 U4969 ( .A(1'b0), .B(_02074__PTR0), .S(_01770__PTR2), .Z(_01912__PTR64) );
  MUX2_X1 U4970 ( .A(1'b0), .B(_02074__PTR1), .S(_01770__PTR2), .Z(_01912__PTR65) );
  MUX2_X1 U4971 ( .A(1'b0), .B(_02074__PTR2), .S(_01770__PTR2), .Z(_01912__PTR66) );
  MUX2_X1 U4972 ( .A(1'b0), .B(_02074__PTR3), .S(_01770__PTR2), .Z(_01912__PTR67) );
  MUX2_X1 U4973 ( .A(1'b0), .B(_02074__PTR4), .S(_01770__PTR2), .Z(_01912__PTR68) );
  MUX2_X1 U4974 ( .A(1'b0), .B(_02074__PTR5), .S(_01770__PTR2), .Z(_01912__PTR69) );
  MUX2_X1 U4975 ( .A(1'b0), .B(_02074__PTR6), .S(_01770__PTR2), .Z(_01912__PTR70) );
  MUX2_X1 U4976 ( .A(1'b0), .B(_02074__PTR7), .S(_01770__PTR2), .Z(_01912__PTR71) );
  MUX2_X1 U4977 ( .A(1'b0), .B(_02073__PTR0), .S(_01770__PTR2), .Z(_01910__PTR64) );
  MUX2_X1 U4978 ( .A(1'b0), .B(_02073__PTR1), .S(_01770__PTR2), .Z(_01910__PTR65) );
  MUX2_X1 U4979 ( .A(1'b0), .B(_02073__PTR2), .S(_01770__PTR2), .Z(_01910__PTR66) );
  MUX2_X1 U4980 ( .A(1'b0), .B(_02073__PTR3), .S(_01770__PTR2), .Z(_01910__PTR67) );
  MUX2_X1 U4981 ( .A(1'b0), .B(_02073__PTR4), .S(_01770__PTR2), .Z(_01910__PTR68) );
  MUX2_X1 U4982 ( .A(1'b0), .B(_02073__PTR5), .S(_01770__PTR2), .Z(_01910__PTR69) );
  MUX2_X1 U4983 ( .A(1'b0), .B(_02073__PTR6), .S(_01770__PTR2), .Z(_01910__PTR70) );
  MUX2_X1 U4984 ( .A(1'b0), .B(_02073__PTR7), .S(_01770__PTR2), .Z(_01910__PTR71) );
  MUX2_X1 U4985 ( .A(1'b0), .B(_02072__PTR0), .S(_01770__PTR2), .Z(_01908__PTR64) );
  MUX2_X1 U4986 ( .A(1'b0), .B(_02072__PTR1), .S(_01770__PTR2), .Z(_01908__PTR65) );
  MUX2_X1 U4987 ( .A(1'b0), .B(_02072__PTR2), .S(_01770__PTR2), .Z(_01908__PTR66) );
  MUX2_X1 U4988 ( .A(1'b0), .B(_02072__PTR3), .S(_01770__PTR2), .Z(_01908__PTR67) );
  MUX2_X1 U4989 ( .A(1'b0), .B(_02072__PTR4), .S(_01770__PTR2), .Z(_01908__PTR68) );
  MUX2_X1 U4990 ( .A(1'b0), .B(_02072__PTR5), .S(_01770__PTR2), .Z(_01908__PTR69) );
  MUX2_X1 U4991 ( .A(1'b0), .B(_02072__PTR6), .S(_01770__PTR2), .Z(_01908__PTR70) );
  MUX2_X1 U4992 ( .A(1'b0), .B(_02072__PTR7), .S(_01770__PTR2), .Z(_01908__PTR71) );
  MUX2_X1 U4993 ( .A(1'b0), .B(_02071__PTR0), .S(_01770__PTR2), .Z(_01906__PTR64) );
  MUX2_X1 U4994 ( .A(1'b0), .B(_02071__PTR1), .S(_01770__PTR2), .Z(_01906__PTR65) );
  MUX2_X1 U4995 ( .A(1'b0), .B(_02071__PTR2), .S(_01770__PTR2), .Z(_01906__PTR66) );
  MUX2_X1 U4996 ( .A(1'b0), .B(_02071__PTR3), .S(_01770__PTR2), .Z(_01906__PTR67) );
  MUX2_X1 U4997 ( .A(1'b0), .B(_02071__PTR4), .S(_01770__PTR2), .Z(_01906__PTR68) );
  MUX2_X1 U4998 ( .A(1'b0), .B(_02071__PTR5), .S(_01770__PTR2), .Z(_01906__PTR69) );
  MUX2_X1 U4999 ( .A(1'b0), .B(_02071__PTR6), .S(_01770__PTR2), .Z(_01906__PTR70) );
  MUX2_X1 U5000 ( .A(1'b0), .B(_02071__PTR7), .S(_01770__PTR2), .Z(_01906__PTR71) );
  MUX2_X1 U5001 ( .A(1'b0), .B(_02070__PTR0), .S(_01770__PTR2), .Z(_01904__PTR64) );
  MUX2_X1 U5002 ( .A(1'b0), .B(_02070__PTR1), .S(_01770__PTR2), .Z(_01904__PTR65) );
  MUX2_X1 U5003 ( .A(1'b0), .B(_02070__PTR2), .S(_01770__PTR2), .Z(_01904__PTR66) );
  MUX2_X1 U5004 ( .A(1'b0), .B(_02070__PTR3), .S(_01770__PTR2), .Z(_01904__PTR67) );
  MUX2_X1 U5005 ( .A(1'b0), .B(_02070__PTR4), .S(_01770__PTR2), .Z(_01904__PTR68) );
  MUX2_X1 U5006 ( .A(1'b0), .B(_02070__PTR5), .S(_01770__PTR2), .Z(_01904__PTR69) );
  MUX2_X1 U5007 ( .A(1'b0), .B(_02070__PTR6), .S(_01770__PTR2), .Z(_01904__PTR70) );
  MUX2_X1 U5008 ( .A(1'b0), .B(_02070__PTR7), .S(_01770__PTR2), .Z(_01904__PTR71) );
  MUX2_X1 U5009 ( .A(1'b0), .B(_02069__PTR0), .S(_01770__PTR2), .Z(_01902__PTR64) );
  MUX2_X1 U5010 ( .A(1'b0), .B(_02069__PTR1), .S(_01770__PTR2), .Z(_01902__PTR65) );
  MUX2_X1 U5011 ( .A(1'b0), .B(_02069__PTR2), .S(_01770__PTR2), .Z(_01902__PTR66) );
  MUX2_X1 U5012 ( .A(1'b0), .B(_02069__PTR3), .S(_01770__PTR2), .Z(_01902__PTR67) );
  MUX2_X1 U5013 ( .A(1'b0), .B(_02069__PTR4), .S(_01770__PTR2), .Z(_01902__PTR68) );
  MUX2_X1 U5014 ( .A(1'b0), .B(_02069__PTR5), .S(_01770__PTR2), .Z(_01902__PTR69) );
  MUX2_X1 U5015 ( .A(1'b0), .B(_02069__PTR6), .S(_01770__PTR2), .Z(_01902__PTR70) );
  MUX2_X1 U5016 ( .A(1'b0), .B(_02069__PTR7), .S(_01770__PTR2), .Z(_01902__PTR71) );
  MUX2_X1 U5017 ( .A(1'b0), .B(_02068__PTR0), .S(_01770__PTR2), .Z(_01900__PTR64) );
  MUX2_X1 U5018 ( .A(1'b0), .B(_02068__PTR1), .S(_01770__PTR2), .Z(_01900__PTR65) );
  MUX2_X1 U5019 ( .A(1'b0), .B(_02068__PTR2), .S(_01770__PTR2), .Z(_01900__PTR66) );
  MUX2_X1 U5020 ( .A(1'b0), .B(_02068__PTR3), .S(_01770__PTR2), .Z(_01900__PTR67) );
  MUX2_X1 U5021 ( .A(1'b0), .B(_02068__PTR4), .S(_01770__PTR2), .Z(_01900__PTR68) );
  MUX2_X1 U5022 ( .A(1'b0), .B(_02068__PTR5), .S(_01770__PTR2), .Z(_01900__PTR69) );
  MUX2_X1 U5023 ( .A(1'b0), .B(_02068__PTR6), .S(_01770__PTR2), .Z(_01900__PTR70) );
  MUX2_X1 U5024 ( .A(1'b0), .B(_02068__PTR7), .S(_01770__PTR2), .Z(_01900__PTR71) );
  MUX2_X1 U5025 ( .A(1'b0), .B(_02067__PTR0), .S(_01770__PTR2), .Z(_01898__PTR64) );
  MUX2_X1 U5026 ( .A(1'b0), .B(_02067__PTR1), .S(_01770__PTR2), .Z(_01898__PTR65) );
  MUX2_X1 U5027 ( .A(1'b0), .B(_02067__PTR2), .S(_01770__PTR2), .Z(_01898__PTR66) );
  MUX2_X1 U5028 ( .A(1'b0), .B(_02067__PTR3), .S(_01770__PTR2), .Z(_01898__PTR67) );
  MUX2_X1 U5029 ( .A(1'b0), .B(_02067__PTR4), .S(_01770__PTR2), .Z(_01898__PTR68) );
  MUX2_X1 U5030 ( .A(1'b0), .B(_02067__PTR5), .S(_01770__PTR2), .Z(_01898__PTR69) );
  MUX2_X1 U5031 ( .A(1'b0), .B(_02067__PTR6), .S(_01770__PTR2), .Z(_01898__PTR70) );
  MUX2_X1 U5032 ( .A(1'b0), .B(_02067__PTR7), .S(_01770__PTR2), .Z(_01898__PTR71) );
  MUX2_X1 U5033 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR0), .Z(_02082__PTR0) );
  MUX2_X1 U5034 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR0), .Z(_02082__PTR1) );
  MUX2_X1 U5035 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR0), .Z(_02082__PTR2) );
  MUX2_X1 U5036 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR0), .Z(_02082__PTR3) );
  MUX2_X1 U5037 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR0), .Z(_02082__PTR4) );
  MUX2_X1 U5038 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR0), .Z(_02082__PTR5) );
  MUX2_X1 U5039 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR0), .Z(_02082__PTR6) );
  MUX2_X1 U5040 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR0), .Z(_02082__PTR7) );
  MUX2_X1 U5041 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR1), .Z(_02081__PTR0) );
  MUX2_X1 U5042 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR1), .Z(_02081__PTR1) );
  MUX2_X1 U5043 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR1), .Z(_02081__PTR2) );
  MUX2_X1 U5044 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR1), .Z(_02081__PTR3) );
  MUX2_X1 U5045 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR1), .Z(_02081__PTR4) );
  MUX2_X1 U5046 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR1), .Z(_02081__PTR5) );
  MUX2_X1 U5047 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR1), .Z(_02081__PTR6) );
  MUX2_X1 U5048 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR1), .Z(_02081__PTR7) );
  MUX2_X1 U5049 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR2), .Z(_02080__PTR0) );
  MUX2_X1 U5050 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR2), .Z(_02080__PTR1) );
  MUX2_X1 U5051 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR2), .Z(_02080__PTR2) );
  MUX2_X1 U5052 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR2), .Z(_02080__PTR3) );
  MUX2_X1 U5053 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR2), .Z(_02080__PTR4) );
  MUX2_X1 U5054 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR2), .Z(_02080__PTR5) );
  MUX2_X1 U5055 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR2), .Z(_02080__PTR6) );
  MUX2_X1 U5056 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR2), .Z(_02080__PTR7) );
  MUX2_X1 U5057 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR3), .Z(_02079__PTR0) );
  MUX2_X1 U5058 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR3), .Z(_02079__PTR1) );
  MUX2_X1 U5059 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR3), .Z(_02079__PTR2) );
  MUX2_X1 U5060 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR3), .Z(_02079__PTR3) );
  MUX2_X1 U5061 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR3), .Z(_02079__PTR4) );
  MUX2_X1 U5062 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR3), .Z(_02079__PTR5) );
  MUX2_X1 U5063 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR3), .Z(_02079__PTR6) );
  MUX2_X1 U5064 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR3), .Z(_02079__PTR7) );
  MUX2_X1 U5065 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR4), .Z(_02078__PTR0) );
  MUX2_X1 U5066 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR4), .Z(_02078__PTR1) );
  MUX2_X1 U5067 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR4), .Z(_02078__PTR2) );
  MUX2_X1 U5068 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR4), .Z(_02078__PTR3) );
  MUX2_X1 U5069 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR4), .Z(_02078__PTR4) );
  MUX2_X1 U5070 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR4), .Z(_02078__PTR5) );
  MUX2_X1 U5071 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR4), .Z(_02078__PTR6) );
  MUX2_X1 U5072 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR4), .Z(_02078__PTR7) );
  MUX2_X1 U5073 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR5), .Z(_02077__PTR0) );
  MUX2_X1 U5074 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR5), .Z(_02077__PTR1) );
  MUX2_X1 U5075 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR5), .Z(_02077__PTR2) );
  MUX2_X1 U5076 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR5), .Z(_02077__PTR3) );
  MUX2_X1 U5077 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR5), .Z(_02077__PTR4) );
  MUX2_X1 U5078 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR5), .Z(_02077__PTR5) );
  MUX2_X1 U5079 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR5), .Z(_02077__PTR6) );
  MUX2_X1 U5080 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR5), .Z(_02077__PTR7) );
  MUX2_X1 U5081 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR6), .Z(_02076__PTR0) );
  MUX2_X1 U5082 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR6), .Z(_02076__PTR1) );
  MUX2_X1 U5083 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR6), .Z(_02076__PTR2) );
  MUX2_X1 U5084 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR6), .Z(_02076__PTR3) );
  MUX2_X1 U5085 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR6), .Z(_02076__PTR4) );
  MUX2_X1 U5086 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR6), .Z(_02076__PTR5) );
  MUX2_X1 U5087 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR6), .Z(_02076__PTR6) );
  MUX2_X1 U5088 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR6), .Z(_02076__PTR7) );
  MUX2_X1 U5089 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR7), .Z(_02075__PTR0) );
  MUX2_X1 U5090 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR7), .Z(_02075__PTR1) );
  MUX2_X1 U5091 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR7), .Z(_02075__PTR2) );
  MUX2_X1 U5092 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR7), .Z(_02075__PTR3) );
  MUX2_X1 U5093 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR7), .Z(_02075__PTR4) );
  MUX2_X1 U5094 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR7), .Z(_02075__PTR5) );
  MUX2_X1 U5095 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR7), .Z(_02075__PTR6) );
  MUX2_X1 U5096 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR7), .Z(_02075__PTR7) );
  MUX2_X1 U5097 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR8), .Z(_02074__PTR0) );
  MUX2_X1 U5098 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR8), .Z(_02074__PTR1) );
  MUX2_X1 U5099 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR8), .Z(_02074__PTR2) );
  MUX2_X1 U5100 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR8), .Z(_02074__PTR3) );
  MUX2_X1 U5101 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR8), .Z(_02074__PTR4) );
  MUX2_X1 U5102 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR8), .Z(_02074__PTR5) );
  MUX2_X1 U5103 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR8), .Z(_02074__PTR6) );
  MUX2_X1 U5104 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR8), .Z(_02074__PTR7) );
  MUX2_X1 U5105 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR9), .Z(_02073__PTR0) );
  MUX2_X1 U5106 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR9), .Z(_02073__PTR1) );
  MUX2_X1 U5107 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR9), .Z(_02073__PTR2) );
  MUX2_X1 U5108 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR9), .Z(_02073__PTR3) );
  MUX2_X1 U5109 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR9), .Z(_02073__PTR4) );
  MUX2_X1 U5110 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR9), .Z(_02073__PTR5) );
  MUX2_X1 U5111 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR9), .Z(_02073__PTR6) );
  MUX2_X1 U5112 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR9), .Z(_02073__PTR7) );
  MUX2_X1 U5113 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR10), .Z(_02072__PTR0) );
  MUX2_X1 U5114 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR10), .Z(_02072__PTR1) );
  MUX2_X1 U5115 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR10), .Z(_02072__PTR2) );
  MUX2_X1 U5116 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR10), .Z(_02072__PTR3) );
  MUX2_X1 U5117 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR10), .Z(_02072__PTR4) );
  MUX2_X1 U5118 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR10), .Z(_02072__PTR5) );
  MUX2_X1 U5119 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR10), .Z(_02072__PTR6) );
  MUX2_X1 U5120 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR10), .Z(_02072__PTR7) );
  MUX2_X1 U5121 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR11), .Z(_02071__PTR0) );
  MUX2_X1 U5122 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR11), .Z(_02071__PTR1) );
  MUX2_X1 U5123 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR11), .Z(_02071__PTR2) );
  MUX2_X1 U5124 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR11), .Z(_02071__PTR3) );
  MUX2_X1 U5125 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR11), .Z(_02071__PTR4) );
  MUX2_X1 U5126 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR11), .Z(_02071__PTR5) );
  MUX2_X1 U5127 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR11), .Z(_02071__PTR6) );
  MUX2_X1 U5128 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR11), .Z(_02071__PTR7) );
  MUX2_X1 U5129 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR12), .Z(_02070__PTR0) );
  MUX2_X1 U5130 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR12), .Z(_02070__PTR1) );
  MUX2_X1 U5131 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR12), .Z(_02070__PTR2) );
  MUX2_X1 U5132 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR12), .Z(_02070__PTR3) );
  MUX2_X1 U5133 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR12), .Z(_02070__PTR4) );
  MUX2_X1 U5134 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR12), .Z(_02070__PTR5) );
  MUX2_X1 U5135 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR12), .Z(_02070__PTR6) );
  MUX2_X1 U5136 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR12), .Z(_02070__PTR7) );
  MUX2_X1 U5137 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR13), .Z(_02069__PTR0) );
  MUX2_X1 U5138 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR13), .Z(_02069__PTR1) );
  MUX2_X1 U5139 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR13), .Z(_02069__PTR2) );
  MUX2_X1 U5140 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR13), .Z(_02069__PTR3) );
  MUX2_X1 U5141 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR13), .Z(_02069__PTR4) );
  MUX2_X1 U5142 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR13), .Z(_02069__PTR5) );
  MUX2_X1 U5143 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR13), .Z(_02069__PTR6) );
  MUX2_X1 U5144 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR13), .Z(_02069__PTR7) );
  MUX2_X1 U5145 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR14), .Z(_02068__PTR0) );
  MUX2_X1 U5146 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR14), .Z(_02068__PTR1) );
  MUX2_X1 U5147 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR14), .Z(_02068__PTR2) );
  MUX2_X1 U5148 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR14), .Z(_02068__PTR3) );
  MUX2_X1 U5149 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR14), .Z(_02068__PTR4) );
  MUX2_X1 U5150 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR14), .Z(_02068__PTR5) );
  MUX2_X1 U5151 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR14), .Z(_02068__PTR6) );
  MUX2_X1 U5152 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR14), .Z(_02068__PTR7) );
  MUX2_X1 U5153 ( .A(1'b0), .B(_01883__PTR0), .S(_01835__PTR15), .Z(_02067__PTR0) );
  MUX2_X1 U5154 ( .A(1'b0), .B(_01883__PTR1), .S(_01835__PTR15), .Z(_02067__PTR1) );
  MUX2_X1 U5155 ( .A(1'b0), .B(_01883__PTR2), .S(_01835__PTR15), .Z(_02067__PTR2) );
  MUX2_X1 U5156 ( .A(1'b0), .B(_01883__PTR3), .S(_01835__PTR15), .Z(_02067__PTR3) );
  MUX2_X1 U5157 ( .A(1'b0), .B(_01883__PTR4), .S(_01835__PTR15), .Z(_02067__PTR4) );
  MUX2_X1 U5158 ( .A(1'b0), .B(_01883__PTR5), .S(_01835__PTR15), .Z(_02067__PTR5) );
  MUX2_X1 U5159 ( .A(1'b0), .B(_01883__PTR6), .S(_01835__PTR15), .Z(_02067__PTR6) );
  MUX2_X1 U5160 ( .A(1'b0), .B(_01883__PTR7), .S(_01835__PTR15), .Z(_02067__PTR7) );
  MUX2_X1 U5161 ( .A(1'b0), .B(_02066__PTR0), .S(_01894__PTR28), .Z(_01930__PTR56) );
  MUX2_X1 U5162 ( .A(1'b0), .B(_02066__PTR4), .S(_01894__PTR28), .Z(_01930__PTR60) );
  MUX2_X1 U5163 ( .A(1'b0), .B(1'b1), .S(P1_P1_Flush), .Z(_02066__PTR0) );
  MUX2_X1 U5164 ( .A(1'b0), .B(1'b0), .S(P1_P1_Flush), .Z(_02066__PTR4) );
  MUX2_X1 U5165 ( .A(P1_P1_InstQueueRd_Addr_PTR0), .B(_02065__PTR0), .S(P1_P1_Flush), .Z(_01932__PTR56) );
  MUX2_X1 U5166 ( .A(P1_P1_InstQueueRd_Addr_PTR1), .B(_02065__PTR1), .S(P1_P1_Flush), .Z(_01932__PTR57) );
  MUX2_X1 U5167 ( .A(P1_P1_InstQueueRd_Addr_PTR2), .B(_02065__PTR2), .S(P1_P1_Flush), .Z(_01932__PTR58) );
  MUX2_X1 U5168 ( .A(P1_P1_InstQueueRd_Addr_PTR3), .B(1'b0), .S(P1_P1_Flush), .Z(_01932__PTR59) );
  MUX2_X1 U5169 ( .A(P1_P1_InstQueueRd_Addr_PTR4), .B(1'b0), .S(P1_P1_Flush), .Z(_01932__PTR60) );
  MUX2_X1 U5170 ( .A(1'b1), .B(_02084__PTR0), .S(P1_P1_InstAddrPointer_PTR0), .Z(_02065__PTR0) );
  MUX2_X1 U5171 ( .A(1'b0), .B(_02831__PTR1), .S(P1_P1_InstAddrPointer_PTR0), .Z(_02065__PTR1) );
  MUX2_X1 U5172 ( .A(1'b0), .B(_02830__PTR1), .S(P1_P1_InstAddrPointer_PTR0), .Z(_02065__PTR2) );
  MUX2_X1 U5173 ( .A(_02949__PTR1), .B(P1_P1_InstAddrPointer_PTR1), .S(_02744__PTR31), .Z(_02829__PTR1) );
  MUX2_X1 U5174 ( .A(1'b1), .B(1'b0), .S(P1_READY_n), .Z(_01894__PTR26) );
  MUX2_X1 U5175 ( .A(1'b0), .B(1'b0), .S(P1_READY_n), .Z(_01849__PTR6) );
  MUX2_X1 U5176 ( .A(_02121__PTR0), .B(1'b1), .S(_02064_), .Z(_01894__PTR20) );
  MUX2_X1 U5177 ( .A(_02121__PTR1), .B(1'b1), .S(_02064_), .Z(_01894__PTR21) );
  MUX2_X1 U5178 ( .A(_02121__PTR2), .B(1'b1), .S(_02064_), .Z(_01894__PTR22) );
  MUX2_X1 U5179 ( .A(_02121__PTR3), .B(1'b0), .S(_02064_), .Z(_01894__PTR23) );
  MUX2_X1 U5180 ( .A(P1_Datao_PTR16), .B(_02046__PTR16), .S(_02006_), .Z(_02114__PTR48) );
  MUX2_X1 U5181 ( .A(P1_Datao_PTR17), .B(_02046__PTR17), .S(_02006_), .Z(_02114__PTR49) );
  MUX2_X1 U5182 ( .A(P1_Datao_PTR18), .B(_02046__PTR18), .S(_02006_), .Z(_02114__PTR50) );
  MUX2_X1 U5183 ( .A(P1_Datao_PTR19), .B(_02046__PTR19), .S(_02006_), .Z(_02114__PTR51) );
  MUX2_X1 U5184 ( .A(P1_Datao_PTR20), .B(_02046__PTR20), .S(_02006_), .Z(_02114__PTR52) );
  MUX2_X1 U5185 ( .A(P1_Datao_PTR21), .B(_02046__PTR21), .S(_02006_), .Z(_02114__PTR53) );
  MUX2_X1 U5186 ( .A(P1_Datao_PTR22), .B(_02046__PTR22), .S(_02006_), .Z(_02114__PTR54) );
  MUX2_X1 U5187 ( .A(P1_Datao_PTR23), .B(_02046__PTR23), .S(_02006_), .Z(_02114__PTR55) );
  MUX2_X1 U5188 ( .A(P1_Datao_PTR24), .B(_02046__PTR24), .S(_02006_), .Z(_02114__PTR56) );
  MUX2_X1 U5189 ( .A(P1_Datao_PTR25), .B(_02046__PTR25), .S(_02006_), .Z(_02114__PTR57) );
  MUX2_X1 U5190 ( .A(P1_Datao_PTR26), .B(_02046__PTR26), .S(_02006_), .Z(_02114__PTR58) );
  MUX2_X1 U5191 ( .A(P1_Datao_PTR27), .B(_02046__PTR27), .S(_02006_), .Z(_02114__PTR59) );
  MUX2_X1 U5192 ( .A(P1_Datao_PTR28), .B(_02046__PTR28), .S(_02006_), .Z(_02114__PTR60) );
  MUX2_X1 U5193 ( .A(P1_Datao_PTR29), .B(_02046__PTR29), .S(_02006_), .Z(_02114__PTR61) );
  MUX2_X1 U5194 ( .A(P1_Datao_PTR30), .B(_02046__PTR30), .S(_02006_), .Z(_02114__PTR62) );
  MUX2_X1 U5195 ( .A(P1_Datao_PTR31), .B(_02031__PTR31), .S(_02006_), .Z(_02114__PTR95) );
  MUX2_X1 U5196 ( .A(P1_Datao_PTR0), .B(_02031__PTR0), .S(_02006_), .Z(_02114__PTR64) );
  MUX2_X1 U5197 ( .A(P1_Datao_PTR1), .B(_02031__PTR1), .S(_02006_), .Z(_02114__PTR65) );
  MUX2_X1 U5198 ( .A(P1_Datao_PTR2), .B(_02031__PTR2), .S(_02006_), .Z(_02114__PTR66) );
  MUX2_X1 U5199 ( .A(P1_Datao_PTR3), .B(_02031__PTR3), .S(_02006_), .Z(_02114__PTR67) );
  MUX2_X1 U5200 ( .A(P1_Datao_PTR4), .B(_02031__PTR4), .S(_02006_), .Z(_02114__PTR68) );
  MUX2_X1 U5201 ( .A(P1_Datao_PTR5), .B(_02031__PTR5), .S(_02006_), .Z(_02114__PTR69) );
  MUX2_X1 U5202 ( .A(P1_Datao_PTR6), .B(_02031__PTR6), .S(_02006_), .Z(_02114__PTR70) );
  MUX2_X1 U5203 ( .A(P1_Datao_PTR7), .B(_02031__PTR7), .S(_02006_), .Z(_02114__PTR71) );
  MUX2_X1 U5204 ( .A(P1_Datao_PTR8), .B(_02031__PTR8), .S(_02006_), .Z(_02114__PTR72) );
  MUX2_X1 U5205 ( .A(P1_Datao_PTR9), .B(_02031__PTR9), .S(_02006_), .Z(_02114__PTR73) );
  MUX2_X1 U5206 ( .A(P1_Datao_PTR10), .B(_02031__PTR10), .S(_02006_), .Z(_02114__PTR74) );
  MUX2_X1 U5207 ( .A(P1_Datao_PTR11), .B(_02031__PTR11), .S(_02006_), .Z(_02114__PTR75) );
  MUX2_X1 U5208 ( .A(P1_Datao_PTR12), .B(_02031__PTR12), .S(_02006_), .Z(_02114__PTR76) );
  MUX2_X1 U5209 ( .A(P1_Datao_PTR13), .B(_02031__PTR13), .S(_02006_), .Z(_02114__PTR77) );
  MUX2_X1 U5210 ( .A(P1_Datao_PTR14), .B(_02031__PTR14), .S(_02006_), .Z(_02114__PTR78) );
  MUX2_X1 U5211 ( .A(P1_Datao_PTR15), .B(_02031__PTR15), .S(_02006_), .Z(_02114__PTR79) );
  MUX2_X1 U5212 ( .A(P1_Datao_PTR16), .B(_02031__PTR16), .S(_02006_), .Z(_02114__PTR80) );
  MUX2_X1 U5213 ( .A(P1_Datao_PTR17), .B(_02031__PTR17), .S(_02006_), .Z(_02114__PTR81) );
  MUX2_X1 U5214 ( .A(P1_Datao_PTR18), .B(_02031__PTR18), .S(_02006_), .Z(_02114__PTR82) );
  MUX2_X1 U5215 ( .A(P1_Datao_PTR19), .B(_02031__PTR19), .S(_02006_), .Z(_02114__PTR83) );
  MUX2_X1 U5216 ( .A(P1_Datao_PTR20), .B(_02031__PTR20), .S(_02006_), .Z(_02114__PTR84) );
  MUX2_X1 U5217 ( .A(P1_Datao_PTR21), .B(_02031__PTR21), .S(_02006_), .Z(_02114__PTR85) );
  MUX2_X1 U5218 ( .A(P1_Datao_PTR22), .B(_02031__PTR22), .S(_02006_), .Z(_02114__PTR86) );
  MUX2_X1 U5219 ( .A(P1_Datao_PTR23), .B(_02031__PTR23), .S(_02006_), .Z(_02114__PTR87) );
  MUX2_X1 U5220 ( .A(P1_Datao_PTR24), .B(_02031__PTR24), .S(_02006_), .Z(_02114__PTR88) );
  MUX2_X1 U5221 ( .A(P1_Datao_PTR25), .B(_02031__PTR25), .S(_02006_), .Z(_02114__PTR89) );
  MUX2_X1 U5222 ( .A(P1_Datao_PTR26), .B(_02031__PTR26), .S(_02006_), .Z(_02114__PTR90) );
  MUX2_X1 U5223 ( .A(P1_Datao_PTR27), .B(_02031__PTR27), .S(_02006_), .Z(_02114__PTR91) );
  MUX2_X1 U5224 ( .A(P1_Datao_PTR28), .B(_02031__PTR28), .S(_02006_), .Z(_02114__PTR92) );
  MUX2_X1 U5225 ( .A(P1_Datao_PTR29), .B(_02031__PTR29), .S(_02006_), .Z(_02114__PTR93) );
  MUX2_X1 U5226 ( .A(P1_Datao_PTR30), .B(_02031__PTR30), .S(_02006_), .Z(_02114__PTR94) );
  MUX2_X1 U5227 ( .A(P1_RequestPending), .B(_02047_), .S(_02006_), .Z(_01861__PTR0) );
  MUX2_X1 U5228 ( .A(1'b1), .B(P1_READY_n), .S(_02025_), .Z(_02047_) );
  MUX2_X1 U5229 ( .A(P1_MemoryFetch), .B(1'b0), .S(_02006_), .Z(_01868__PTR0) );
  MUX2_X1 U5230 ( .A(1'b0), .B(_02036_), .S(_02006_), .Z(_01853__PTR0) );
  MUX2_X1 U5231 ( .A(1'b1), .B(_02035_), .S(_02006_), .Z(_01857__PTR0) );
  MUX2_X1 U5232 ( .A(P1_P1_State2_PTR0), .B(_02034__PTR0), .S(_02006_), .Z(_02118__PTR4) );
  MUX2_X1 U5233 ( .A(P1_P1_State2_PTR1), .B(_02034__PTR1), .S(_02006_), .Z(_02118__PTR5) );
  MUX2_X1 U5234 ( .A(P1_P1_State2_PTR2), .B(_02034__PTR2), .S(_02006_), .Z(_02118__PTR6) );
  MUX2_X1 U5235 ( .A(P1_P1_State2_PTR3), .B(_02034__PTR3), .S(_02006_), .Z(_02118__PTR7) );
  MUX2_X1 U5236 ( .A(P1_Datao_PTR16), .B(1'b0), .S(_02025_), .Z(_02046__PTR16) );
  MUX2_X1 U5237 ( .A(P1_Datao_PTR17), .B(1'b0), .S(_02025_), .Z(_02046__PTR17) );
  MUX2_X1 U5238 ( .A(P1_Datao_PTR18), .B(1'b0), .S(_02025_), .Z(_02046__PTR18) );
  MUX2_X1 U5239 ( .A(P1_Datao_PTR19), .B(1'b0), .S(_02025_), .Z(_02046__PTR19) );
  MUX2_X1 U5240 ( .A(P1_Datao_PTR20), .B(1'b0), .S(_02025_), .Z(_02046__PTR20) );
  MUX2_X1 U5241 ( .A(P1_Datao_PTR21), .B(1'b0), .S(_02025_), .Z(_02046__PTR21) );
  MUX2_X1 U5242 ( .A(P1_Datao_PTR22), .B(1'b0), .S(_02025_), .Z(_02046__PTR22) );
  MUX2_X1 U5243 ( .A(P1_Datao_PTR23), .B(1'b0), .S(_02025_), .Z(_02046__PTR23) );
  MUX2_X1 U5244 ( .A(P1_Datao_PTR24), .B(1'b0), .S(_02025_), .Z(_02046__PTR24) );
  MUX2_X1 U5245 ( .A(P1_Datao_PTR25), .B(1'b0), .S(_02025_), .Z(_02046__PTR25) );
  MUX2_X1 U5246 ( .A(P1_Datao_PTR26), .B(1'b0), .S(_02025_), .Z(_02046__PTR26) );
  MUX2_X1 U5247 ( .A(P1_Datao_PTR27), .B(1'b0), .S(_02025_), .Z(_02046__PTR27) );
  MUX2_X1 U5248 ( .A(P1_Datao_PTR28), .B(1'b0), .S(_02025_), .Z(_02046__PTR28) );
  MUX2_X1 U5249 ( .A(P1_Datao_PTR29), .B(1'b0), .S(_02025_), .Z(_02046__PTR29) );
  MUX2_X1 U5250 ( .A(P1_Datao_PTR30), .B(1'b0), .S(_02025_), .Z(_02046__PTR30) );
  MUX2_X1 U5251 ( .A(P1_Datao_PTR31), .B(1'b0), .S(_02025_), .Z(_02031__PTR31) );
  MUX2_X1 U5252 ( .A(P1_Datao_PTR0), .B(P1_EAX_PTR0), .S(_02025_), .Z(_02031__PTR0) );
  MUX2_X1 U5253 ( .A(P1_Datao_PTR1), .B(P1_EAX_PTR1), .S(_02025_), .Z(_02031__PTR1) );
  MUX2_X1 U5254 ( .A(P1_Datao_PTR2), .B(P1_EAX_PTR2), .S(_02025_), .Z(_02031__PTR2) );
  MUX2_X1 U5255 ( .A(P1_Datao_PTR3), .B(P1_EAX_PTR3), .S(_02025_), .Z(_02031__PTR3) );
  MUX2_X1 U5256 ( .A(P1_Datao_PTR4), .B(P1_EAX_PTR4), .S(_02025_), .Z(_02031__PTR4) );
  MUX2_X1 U5257 ( .A(P1_Datao_PTR5), .B(P1_EAX_PTR5), .S(_02025_), .Z(_02031__PTR5) );
  MUX2_X1 U5258 ( .A(P1_Datao_PTR6), .B(P1_EAX_PTR6), .S(_02025_), .Z(_02031__PTR6) );
  MUX2_X1 U5259 ( .A(P1_Datao_PTR7), .B(P1_EAX_PTR7), .S(_02025_), .Z(_02031__PTR7) );
  MUX2_X1 U5260 ( .A(P1_Datao_PTR8), .B(P1_EAX_PTR8), .S(_02025_), .Z(_02031__PTR8) );
  MUX2_X1 U5261 ( .A(P1_Datao_PTR9), .B(P1_EAX_PTR9), .S(_02025_), .Z(_02031__PTR9) );
  MUX2_X1 U5262 ( .A(P1_Datao_PTR10), .B(P1_EAX_PTR10), .S(_02025_), .Z(_02031__PTR10) );
  MUX2_X1 U5263 ( .A(P1_Datao_PTR11), .B(P1_EAX_PTR11), .S(_02025_), .Z(_02031__PTR11) );
  MUX2_X1 U5264 ( .A(P1_Datao_PTR12), .B(P1_EAX_PTR12), .S(_02025_), .Z(_02031__PTR12) );
  MUX2_X1 U5265 ( .A(P1_Datao_PTR13), .B(P1_EAX_PTR13), .S(_02025_), .Z(_02031__PTR13) );
  MUX2_X1 U5266 ( .A(P1_Datao_PTR14), .B(P1_EAX_PTR14), .S(_02025_), .Z(_02031__PTR14) );
  MUX2_X1 U5267 ( .A(P1_Datao_PTR15), .B(P1_EAX_PTR15), .S(_02025_), .Z(_02031__PTR15) );
  MUX2_X1 U5268 ( .A(P1_Datao_PTR16), .B(_02825__PTR0), .S(_02025_), .Z(_02031__PTR16) );
  MUX2_X1 U5269 ( .A(P1_Datao_PTR17), .B(_02826__PTR1), .S(_02025_), .Z(_02031__PTR17) );
  MUX2_X1 U5270 ( .A(P1_Datao_PTR18), .B(_02826__PTR2), .S(_02025_), .Z(_02031__PTR18) );
  MUX2_X1 U5271 ( .A(P1_Datao_PTR19), .B(_02826__PTR3), .S(_02025_), .Z(_02031__PTR19) );
  MUX2_X1 U5272 ( .A(P1_Datao_PTR20), .B(_02826__PTR4), .S(_02025_), .Z(_02031__PTR20) );
  MUX2_X1 U5273 ( .A(P1_Datao_PTR21), .B(_02826__PTR5), .S(_02025_), .Z(_02031__PTR21) );
  MUX2_X1 U5274 ( .A(P1_Datao_PTR22), .B(_02826__PTR6), .S(_02025_), .Z(_02031__PTR22) );
  MUX2_X1 U5275 ( .A(P1_Datao_PTR23), .B(_02826__PTR7), .S(_02025_), .Z(_02031__PTR23) );
  MUX2_X1 U5276 ( .A(P1_Datao_PTR24), .B(_02826__PTR8), .S(_02025_), .Z(_02031__PTR24) );
  MUX2_X1 U5277 ( .A(P1_Datao_PTR25), .B(_02826__PTR9), .S(_02025_), .Z(_02031__PTR25) );
  MUX2_X1 U5278 ( .A(P1_Datao_PTR26), .B(_02826__PTR10), .S(_02025_), .Z(_02031__PTR26) );
  MUX2_X1 U5279 ( .A(P1_Datao_PTR27), .B(_02826__PTR11), .S(_02025_), .Z(_02031__PTR27) );
  MUX2_X1 U5280 ( .A(P1_Datao_PTR28), .B(_02826__PTR12), .S(_02025_), .Z(_02031__PTR28) );
  MUX2_X1 U5281 ( .A(P1_Datao_PTR29), .B(_02826__PTR13), .S(_02025_), .Z(_02031__PTR29) );
  MUX2_X1 U5282 ( .A(P1_Datao_PTR30), .B(_02826__PTR14), .S(_02025_), .Z(_02031__PTR30) );
  MUX2_X1 U5283 ( .A(P1_ReadRequest), .B(1'b0), .S(_02006_), .Z(_01865__PTR0) );
  MUX2_X1 U5284 ( .A(P1_RequestPending), .B(_02032_), .S(_02006_), .Z(_01861__PTR2) );
  MUX2_X1 U5285 ( .A(P1_P1_InstQueueRd_Addr_PTR1), .B(_02020__PTR1), .S(_02025_), .Z(_02038__PTR1) );
  MUX2_X1 U5286 ( .A(P1_P1_InstQueueRd_Addr_PTR2), .B(_02020__PTR2), .S(_02025_), .Z(_02038__PTR2) );
  MUX2_X1 U5287 ( .A(P1_P1_InstQueueRd_Addr_PTR3), .B(_02020__PTR3), .S(_02025_), .Z(_02038__PTR3) );
  MUX2_X1 U5288 ( .A(P1_P1_InstQueueRd_Addr_PTR4), .B(_02020__PTR4), .S(_02025_), .Z(_02038__PTR4) );
  MUX2_X1 U5289 ( .A(P1_P1_InstAddrPointer_PTR1), .B(_02019__PTR1), .S(_02025_), .Z(_02037__PTR1) );
  MUX2_X1 U5290 ( .A(P1_P1_InstAddrPointer_PTR2), .B(_02019__PTR2), .S(_02025_), .Z(_02037__PTR2) );
  MUX2_X1 U5291 ( .A(P1_P1_InstAddrPointer_PTR3), .B(_02019__PTR3), .S(_02025_), .Z(_02037__PTR3) );
  MUX2_X1 U5292 ( .A(P1_P1_InstAddrPointer_PTR4), .B(_02019__PTR4), .S(_02025_), .Z(_02037__PTR4) );
  MUX2_X1 U5293 ( .A(P1_P1_InstAddrPointer_PTR5), .B(_02019__PTR5), .S(_02025_), .Z(_02037__PTR5) );
  MUX2_X1 U5294 ( .A(P1_P1_InstAddrPointer_PTR6), .B(_02019__PTR6), .S(_02025_), .Z(_02037__PTR6) );
  MUX2_X1 U5295 ( .A(P1_P1_InstAddrPointer_PTR7), .B(_02019__PTR7), .S(_02025_), .Z(_02037__PTR7) );
  MUX2_X1 U5296 ( .A(P1_P1_InstAddrPointer_PTR8), .B(_02019__PTR8), .S(_02025_), .Z(_02037__PTR8) );
  MUX2_X1 U5297 ( .A(P1_P1_InstAddrPointer_PTR9), .B(_02019__PTR9), .S(_02025_), .Z(_02037__PTR9) );
  MUX2_X1 U5298 ( .A(P1_P1_InstAddrPointer_PTR10), .B(_02019__PTR10), .S(_02025_), .Z(_02037__PTR10) );
  MUX2_X1 U5299 ( .A(P1_P1_InstAddrPointer_PTR11), .B(_02019__PTR11), .S(_02025_), .Z(_02037__PTR11) );
  MUX2_X1 U5300 ( .A(P1_P1_InstAddrPointer_PTR12), .B(_02019__PTR12), .S(_02025_), .Z(_02037__PTR12) );
  MUX2_X1 U5301 ( .A(P1_P1_InstAddrPointer_PTR13), .B(_02019__PTR13), .S(_02025_), .Z(_02037__PTR13) );
  MUX2_X1 U5302 ( .A(P1_P1_InstAddrPointer_PTR14), .B(_02019__PTR14), .S(_02025_), .Z(_02037__PTR14) );
  MUX2_X1 U5303 ( .A(P1_P1_InstAddrPointer_PTR15), .B(_02019__PTR15), .S(_02025_), .Z(_02037__PTR15) );
  MUX2_X1 U5304 ( .A(P1_P1_InstAddrPointer_PTR16), .B(_02019__PTR16), .S(_02025_), .Z(_02037__PTR16) );
  MUX2_X1 U5305 ( .A(P1_P1_InstAddrPointer_PTR17), .B(_02019__PTR17), .S(_02025_), .Z(_02037__PTR17) );
  MUX2_X1 U5306 ( .A(P1_P1_InstAddrPointer_PTR18), .B(_02019__PTR18), .S(_02025_), .Z(_02037__PTR18) );
  MUX2_X1 U5307 ( .A(P1_P1_InstAddrPointer_PTR19), .B(_02019__PTR19), .S(_02025_), .Z(_02037__PTR19) );
  MUX2_X1 U5308 ( .A(P1_P1_InstAddrPointer_PTR20), .B(_02019__PTR20), .S(_02025_), .Z(_02037__PTR20) );
  MUX2_X1 U5309 ( .A(P1_P1_InstAddrPointer_PTR21), .B(_02019__PTR21), .S(_02025_), .Z(_02037__PTR21) );
  MUX2_X1 U5310 ( .A(P1_P1_InstAddrPointer_PTR22), .B(_02019__PTR22), .S(_02025_), .Z(_02037__PTR22) );
  MUX2_X1 U5311 ( .A(P1_P1_InstAddrPointer_PTR23), .B(_02019__PTR23), .S(_02025_), .Z(_02037__PTR23) );
  MUX2_X1 U5312 ( .A(P1_P1_InstAddrPointer_PTR24), .B(_02019__PTR24), .S(_02025_), .Z(_02037__PTR24) );
  MUX2_X1 U5313 ( .A(P1_P1_InstAddrPointer_PTR25), .B(_02019__PTR25), .S(_02025_), .Z(_02037__PTR25) );
  MUX2_X1 U5314 ( .A(P1_P1_InstAddrPointer_PTR26), .B(_02019__PTR26), .S(_02025_), .Z(_02037__PTR26) );
  MUX2_X1 U5315 ( .A(P1_P1_InstAddrPointer_PTR27), .B(_02019__PTR27), .S(_02025_), .Z(_02037__PTR27) );
  MUX2_X1 U5316 ( .A(P1_P1_InstAddrPointer_PTR28), .B(_02019__PTR28), .S(_02025_), .Z(_02037__PTR28) );
  MUX2_X1 U5317 ( .A(P1_P1_InstAddrPointer_PTR29), .B(_02019__PTR29), .S(_02025_), .Z(_02037__PTR29) );
  MUX2_X1 U5318 ( .A(P1_P1_InstAddrPointer_PTR30), .B(_02019__PTR30), .S(_02025_), .Z(_02037__PTR30) );
  MUX2_X1 U5319 ( .A(P1_P1_InstAddrPointer_PTR31), .B(_02019__PTR31), .S(_02025_), .Z(_02037__PTR31) );
  MUX2_X1 U5320 ( .A(P1_P1_Flush), .B(_02018_), .S(_02025_), .Z(_02036_) );
  MUX2_X1 U5321 ( .A(P1_P1_More), .B(_02017_), .S(_02025_), .Z(_02035_) );
  MUX2_X1 U5322 ( .A(P1_P1_State2_PTR0), .B(_02030__PTR0), .S(_02025_), .Z(_02034__PTR0) );
  MUX2_X1 U5323 ( .A(P1_P1_State2_PTR1), .B(_02030__PTR1), .S(_02025_), .Z(_02034__PTR1) );
  MUX2_X1 U5324 ( .A(P1_P1_State2_PTR2), .B(_02030__PTR2), .S(_02025_), .Z(_02034__PTR2) );
  MUX2_X1 U5325 ( .A(P1_P1_State2_PTR3), .B(_02030__PTR3), .S(_02025_), .Z(_02034__PTR3) );
  MUX2_X1 U5326 ( .A(P1_EBX_PTR0), .B(_02015__PTR0), .S(_02025_), .Z(_02033__PTR0) );
  MUX2_X1 U5327 ( .A(P1_EBX_PTR1), .B(_02029__PTR1), .S(_02025_), .Z(_02033__PTR1) );
  MUX2_X1 U5328 ( .A(P1_EBX_PTR2), .B(_02029__PTR2), .S(_02025_), .Z(_02033__PTR2) );
  MUX2_X1 U5329 ( .A(P1_EBX_PTR3), .B(_02029__PTR3), .S(_02025_), .Z(_02033__PTR3) );
  MUX2_X1 U5330 ( .A(P1_EBX_PTR4), .B(_02029__PTR4), .S(_02025_), .Z(_02033__PTR4) );
  MUX2_X1 U5331 ( .A(P1_EBX_PTR5), .B(_02029__PTR5), .S(_02025_), .Z(_02033__PTR5) );
  MUX2_X1 U5332 ( .A(P1_EBX_PTR6), .B(_02029__PTR6), .S(_02025_), .Z(_02033__PTR6) );
  MUX2_X1 U5333 ( .A(P1_EBX_PTR7), .B(_02029__PTR7), .S(_02025_), .Z(_02033__PTR7) );
  MUX2_X1 U5334 ( .A(P1_EBX_PTR8), .B(_02029__PTR8), .S(_02025_), .Z(_02033__PTR8) );
  MUX2_X1 U5335 ( .A(P1_EBX_PTR9), .B(_02029__PTR9), .S(_02025_), .Z(_02033__PTR9) );
  MUX2_X1 U5336 ( .A(P1_EBX_PTR10), .B(_02029__PTR10), .S(_02025_), .Z(_02033__PTR10) );
  MUX2_X1 U5337 ( .A(P1_EBX_PTR11), .B(_02029__PTR11), .S(_02025_), .Z(_02033__PTR11) );
  MUX2_X1 U5338 ( .A(P1_EBX_PTR12), .B(_02029__PTR12), .S(_02025_), .Z(_02033__PTR12) );
  MUX2_X1 U5339 ( .A(P1_EBX_PTR13), .B(_02029__PTR13), .S(_02025_), .Z(_02033__PTR13) );
  MUX2_X1 U5340 ( .A(P1_EBX_PTR14), .B(_02029__PTR14), .S(_02025_), .Z(_02033__PTR14) );
  MUX2_X1 U5341 ( .A(P1_EBX_PTR15), .B(_02029__PTR15), .S(_02025_), .Z(_02033__PTR15) );
  MUX2_X1 U5342 ( .A(P1_EBX_PTR16), .B(_02029__PTR16), .S(_02025_), .Z(_02033__PTR16) );
  MUX2_X1 U5343 ( .A(P1_EBX_PTR17), .B(_02029__PTR17), .S(_02025_), .Z(_02033__PTR17) );
  MUX2_X1 U5344 ( .A(P1_EBX_PTR18), .B(_02029__PTR18), .S(_02025_), .Z(_02033__PTR18) );
  MUX2_X1 U5345 ( .A(P1_EBX_PTR19), .B(_02029__PTR19), .S(_02025_), .Z(_02033__PTR19) );
  MUX2_X1 U5346 ( .A(P1_EBX_PTR20), .B(_02029__PTR20), .S(_02025_), .Z(_02033__PTR20) );
  MUX2_X1 U5347 ( .A(P1_EBX_PTR21), .B(_02029__PTR21), .S(_02025_), .Z(_02033__PTR21) );
  MUX2_X1 U5348 ( .A(P1_EBX_PTR22), .B(_02029__PTR22), .S(_02025_), .Z(_02033__PTR22) );
  MUX2_X1 U5349 ( .A(P1_EBX_PTR23), .B(_02029__PTR23), .S(_02025_), .Z(_02033__PTR23) );
  MUX2_X1 U5350 ( .A(P1_EBX_PTR24), .B(_02029__PTR24), .S(_02025_), .Z(_02033__PTR24) );
  MUX2_X1 U5351 ( .A(P1_EBX_PTR25), .B(_02029__PTR25), .S(_02025_), .Z(_02033__PTR25) );
  MUX2_X1 U5352 ( .A(P1_EBX_PTR26), .B(_02029__PTR26), .S(_02025_), .Z(_02033__PTR26) );
  MUX2_X1 U5353 ( .A(P1_EBX_PTR27), .B(_02029__PTR27), .S(_02025_), .Z(_02033__PTR27) );
  MUX2_X1 U5354 ( .A(P1_EBX_PTR28), .B(_02029__PTR28), .S(_02025_), .Z(_02033__PTR28) );
  MUX2_X1 U5355 ( .A(P1_EBX_PTR29), .B(_02029__PTR29), .S(_02025_), .Z(_02033__PTR29) );
  MUX2_X1 U5356 ( .A(P1_EBX_PTR30), .B(_02029__PTR30), .S(_02025_), .Z(_02033__PTR30) );
  MUX2_X1 U5357 ( .A(P1_EBX_PTR31), .B(_02029__PTR31), .S(_02025_), .Z(_02033__PTR31) );
  MUX2_X1 U5358 ( .A(1'b1), .B(_02028_), .S(_02025_), .Z(_02032_) );
  MUX2_X1 U5359 ( .A(_02027__PTR0), .B(P1_P1_State2_PTR0), .S(P1_READY_n), .Z(_02030__PTR0) );
  MUX2_X1 U5360 ( .A(_02027__PTR1), .B(P1_P1_State2_PTR1), .S(P1_READY_n), .Z(_02030__PTR1) );
  MUX2_X1 U5361 ( .A(_02027__PTR2), .B(P1_P1_State2_PTR2), .S(P1_READY_n), .Z(_02030__PTR2) );
  MUX2_X1 U5362 ( .A(_02027__PTR3), .B(P1_P1_State2_PTR3), .S(P1_READY_n), .Z(_02030__PTR3) );
  MUX2_X1 U5363 ( .A(_02026__PTR1), .B(P1_EBX_PTR1), .S(P1_READY_n), .Z(_02029__PTR1) );
  MUX2_X1 U5364 ( .A(_02026__PTR2), .B(P1_EBX_PTR2), .S(P1_READY_n), .Z(_02029__PTR2) );
  MUX2_X1 U5365 ( .A(_02026__PTR3), .B(P1_EBX_PTR3), .S(P1_READY_n), .Z(_02029__PTR3) );
  MUX2_X1 U5366 ( .A(_02026__PTR4), .B(P1_EBX_PTR4), .S(P1_READY_n), .Z(_02029__PTR4) );
  MUX2_X1 U5367 ( .A(_02026__PTR5), .B(P1_EBX_PTR5), .S(P1_READY_n), .Z(_02029__PTR5) );
  MUX2_X1 U5368 ( .A(_02026__PTR6), .B(P1_EBX_PTR6), .S(P1_READY_n), .Z(_02029__PTR6) );
  MUX2_X1 U5369 ( .A(_02026__PTR7), .B(P1_EBX_PTR7), .S(P1_READY_n), .Z(_02029__PTR7) );
  MUX2_X1 U5370 ( .A(_02026__PTR8), .B(P1_EBX_PTR8), .S(P1_READY_n), .Z(_02029__PTR8) );
  MUX2_X1 U5371 ( .A(_02026__PTR9), .B(P1_EBX_PTR9), .S(P1_READY_n), .Z(_02029__PTR9) );
  MUX2_X1 U5372 ( .A(_02026__PTR10), .B(P1_EBX_PTR10), .S(P1_READY_n), .Z(_02029__PTR10) );
  MUX2_X1 U5373 ( .A(_02026__PTR11), .B(P1_EBX_PTR11), .S(P1_READY_n), .Z(_02029__PTR11) );
  MUX2_X1 U5374 ( .A(_02026__PTR12), .B(P1_EBX_PTR12), .S(P1_READY_n), .Z(_02029__PTR12) );
  MUX2_X1 U5375 ( .A(_02026__PTR13), .B(P1_EBX_PTR13), .S(P1_READY_n), .Z(_02029__PTR13) );
  MUX2_X1 U5376 ( .A(_02026__PTR14), .B(P1_EBX_PTR14), .S(P1_READY_n), .Z(_02029__PTR14) );
  MUX2_X1 U5377 ( .A(_02026__PTR15), .B(P1_EBX_PTR15), .S(P1_READY_n), .Z(_02029__PTR15) );
  MUX2_X1 U5378 ( .A(_02026__PTR16), .B(P1_EBX_PTR16), .S(P1_READY_n), .Z(_02029__PTR16) );
  MUX2_X1 U5379 ( .A(_02026__PTR17), .B(P1_EBX_PTR17), .S(P1_READY_n), .Z(_02029__PTR17) );
  MUX2_X1 U5380 ( .A(_02026__PTR18), .B(P1_EBX_PTR18), .S(P1_READY_n), .Z(_02029__PTR18) );
  MUX2_X1 U5381 ( .A(_02026__PTR19), .B(P1_EBX_PTR19), .S(P1_READY_n), .Z(_02029__PTR19) );
  MUX2_X1 U5382 ( .A(_02026__PTR20), .B(P1_EBX_PTR20), .S(P1_READY_n), .Z(_02029__PTR20) );
  MUX2_X1 U5383 ( .A(_02026__PTR21), .B(P1_EBX_PTR21), .S(P1_READY_n), .Z(_02029__PTR21) );
  MUX2_X1 U5384 ( .A(_02026__PTR22), .B(P1_EBX_PTR22), .S(P1_READY_n), .Z(_02029__PTR22) );
  MUX2_X1 U5385 ( .A(_02026__PTR23), .B(P1_EBX_PTR23), .S(P1_READY_n), .Z(_02029__PTR23) );
  MUX2_X1 U5386 ( .A(_02026__PTR24), .B(P1_EBX_PTR24), .S(P1_READY_n), .Z(_02029__PTR24) );
  MUX2_X1 U5387 ( .A(_02026__PTR25), .B(P1_EBX_PTR25), .S(P1_READY_n), .Z(_02029__PTR25) );
  MUX2_X1 U5388 ( .A(_02026__PTR26), .B(P1_EBX_PTR26), .S(P1_READY_n), .Z(_02029__PTR26) );
  MUX2_X1 U5389 ( .A(_02026__PTR27), .B(P1_EBX_PTR27), .S(P1_READY_n), .Z(_02029__PTR27) );
  MUX2_X1 U5390 ( .A(_02026__PTR28), .B(P1_EBX_PTR28), .S(P1_READY_n), .Z(_02029__PTR28) );
  MUX2_X1 U5391 ( .A(_02026__PTR29), .B(P1_EBX_PTR29), .S(P1_READY_n), .Z(_02029__PTR29) );
  MUX2_X1 U5392 ( .A(_02026__PTR30), .B(P1_EBX_PTR30), .S(P1_READY_n), .Z(_02029__PTR30) );
  MUX2_X1 U5393 ( .A(_02026__PTR31), .B(P1_EBX_PTR31), .S(P1_READY_n), .Z(_02029__PTR31) );
  MUX2_X1 U5394 ( .A(_01894__PTR9), .B(1'b1), .S(P1_READY_n), .Z(_02028_) );
  MUX2_X1 U5395 ( .A(1'b0), .B(P1_P1_State2_PTR0), .S(P1_StateBS16), .Z(_02027__PTR0) );
  MUX2_X1 U5396 ( .A(1'b1), .B(P1_P1_State2_PTR1), .S(P1_StateBS16), .Z(_02027__PTR1) );
  MUX2_X1 U5397 ( .A(1'b1), .B(P1_P1_State2_PTR2), .S(P1_StateBS16), .Z(_02027__PTR2) );
  MUX2_X1 U5398 ( .A(1'b0), .B(P1_P1_State2_PTR3), .S(P1_StateBS16), .Z(_02027__PTR3) );
  MUX2_X1 U5399 ( .A(_01882__PTR7), .B(P1_EBX_PTR1), .S(P1_StateBS16), .Z(_02026__PTR1) );
  MUX2_X1 U5400 ( .A(_02822__PTR1), .B(P1_EBX_PTR2), .S(P1_StateBS16), .Z(_02026__PTR2) );
  MUX2_X1 U5401 ( .A(_02822__PTR2), .B(P1_EBX_PTR3), .S(P1_StateBS16), .Z(_02026__PTR3) );
  MUX2_X1 U5402 ( .A(_02822__PTR3), .B(P1_EBX_PTR4), .S(P1_StateBS16), .Z(_02026__PTR4) );
  MUX2_X1 U5403 ( .A(_02822__PTR4), .B(P1_EBX_PTR5), .S(P1_StateBS16), .Z(_02026__PTR5) );
  MUX2_X1 U5404 ( .A(_02822__PTR5), .B(P1_EBX_PTR6), .S(P1_StateBS16), .Z(_02026__PTR6) );
  MUX2_X1 U5405 ( .A(_02822__PTR6), .B(P1_EBX_PTR7), .S(P1_StateBS16), .Z(_02026__PTR7) );
  MUX2_X1 U5406 ( .A(_02822__PTR7), .B(P1_EBX_PTR8), .S(P1_StateBS16), .Z(_02026__PTR8) );
  MUX2_X1 U5407 ( .A(_02822__PTR8), .B(P1_EBX_PTR9), .S(P1_StateBS16), .Z(_02026__PTR9) );
  MUX2_X1 U5408 ( .A(_02822__PTR9), .B(P1_EBX_PTR10), .S(P1_StateBS16), .Z(_02026__PTR10) );
  MUX2_X1 U5409 ( .A(_02822__PTR10), .B(P1_EBX_PTR11), .S(P1_StateBS16), .Z(_02026__PTR11) );
  MUX2_X1 U5410 ( .A(_02822__PTR11), .B(P1_EBX_PTR12), .S(P1_StateBS16), .Z(_02026__PTR12) );
  MUX2_X1 U5411 ( .A(_02822__PTR12), .B(P1_EBX_PTR13), .S(P1_StateBS16), .Z(_02026__PTR13) );
  MUX2_X1 U5412 ( .A(_02822__PTR13), .B(P1_EBX_PTR14), .S(P1_StateBS16), .Z(_02026__PTR14) );
  MUX2_X1 U5413 ( .A(_02822__PTR14), .B(P1_EBX_PTR15), .S(P1_StateBS16), .Z(_02026__PTR15) );
  MUX2_X1 U5414 ( .A(_02822__PTR15), .B(P1_EBX_PTR16), .S(P1_StateBS16), .Z(_02026__PTR16) );
  MUX2_X1 U5415 ( .A(_02822__PTR16), .B(P1_EBX_PTR17), .S(P1_StateBS16), .Z(_02026__PTR17) );
  MUX2_X1 U5416 ( .A(_02822__PTR17), .B(P1_EBX_PTR18), .S(P1_StateBS16), .Z(_02026__PTR18) );
  MUX2_X1 U5417 ( .A(_02822__PTR18), .B(P1_EBX_PTR19), .S(P1_StateBS16), .Z(_02026__PTR19) );
  MUX2_X1 U5418 ( .A(_02822__PTR19), .B(P1_EBX_PTR20), .S(P1_StateBS16), .Z(_02026__PTR20) );
  MUX2_X1 U5419 ( .A(_02822__PTR20), .B(P1_EBX_PTR21), .S(P1_StateBS16), .Z(_02026__PTR21) );
  MUX2_X1 U5420 ( .A(_02822__PTR21), .B(P1_EBX_PTR22), .S(P1_StateBS16), .Z(_02026__PTR22) );
  MUX2_X1 U5421 ( .A(_02822__PTR22), .B(P1_EBX_PTR23), .S(P1_StateBS16), .Z(_02026__PTR23) );
  MUX2_X1 U5422 ( .A(_02822__PTR23), .B(P1_EBX_PTR24), .S(P1_StateBS16), .Z(_02026__PTR24) );
  MUX2_X1 U5423 ( .A(_02822__PTR24), .B(P1_EBX_PTR25), .S(P1_StateBS16), .Z(_02026__PTR25) );
  MUX2_X1 U5424 ( .A(_02822__PTR25), .B(P1_EBX_PTR26), .S(P1_StateBS16), .Z(_02026__PTR26) );
  MUX2_X1 U5425 ( .A(_02822__PTR26), .B(P1_EBX_PTR27), .S(P1_StateBS16), .Z(_02026__PTR27) );
  MUX2_X1 U5426 ( .A(_02822__PTR27), .B(P1_EBX_PTR28), .S(P1_StateBS16), .Z(_02026__PTR28) );
  MUX2_X1 U5427 ( .A(_02822__PTR28), .B(P1_EBX_PTR29), .S(P1_StateBS16), .Z(_02026__PTR29) );
  MUX2_X1 U5428 ( .A(_02822__PTR29), .B(P1_EBX_PTR30), .S(P1_StateBS16), .Z(_02026__PTR30) );
  MUX2_X1 U5429 ( .A(_02822__PTR30), .B(P1_EBX_PTR31), .S(P1_StateBS16), .Z(_02026__PTR31) );
  MUX2_X1 U5430 ( .A(_02818__PTR3), .B(P1_P1_InstQueueRd_Addr_PTR4), .S(P1_READY_n), .Z(_02045__PTR4) );
  MUX2_X1 U5431 ( .A(_01890__PTR4), .B(P1_P1_InstQueueRd_Addr_PTR1), .S(P1_READY_n), .Z(_02020__PTR1) );
  MUX2_X1 U5432 ( .A(_01890__PTR5), .B(P1_P1_InstQueueRd_Addr_PTR2), .S(P1_READY_n), .Z(_02020__PTR2) );
  MUX2_X1 U5433 ( .A(_01890__PTR6), .B(P1_P1_InstQueueRd_Addr_PTR3), .S(P1_READY_n), .Z(_02020__PTR3) );
  MUX2_X1 U5434 ( .A(1'b0), .B(P1_P1_InstQueueRd_Addr_PTR4), .S(P1_READY_n), .Z(_02020__PTR4) );
  MUX2_X1 U5435 ( .A(P1_P1_lWord_PTR0), .B(P1_EAX_PTR0), .S(_02006_), .Z(_02111__PTR16) );
  MUX2_X1 U5436 ( .A(P1_P1_lWord_PTR1), .B(P1_EAX_PTR1), .S(_02006_), .Z(_02111__PTR17) );
  MUX2_X1 U5437 ( .A(P1_P1_lWord_PTR2), .B(P1_EAX_PTR2), .S(_02006_), .Z(_02111__PTR18) );
  MUX2_X1 U5438 ( .A(P1_P1_lWord_PTR3), .B(P1_EAX_PTR3), .S(_02006_), .Z(_02111__PTR19) );
  MUX2_X1 U5439 ( .A(P1_P1_lWord_PTR4), .B(P1_EAX_PTR4), .S(_02006_), .Z(_02111__PTR20) );
  MUX2_X1 U5440 ( .A(P1_P1_lWord_PTR5), .B(P1_EAX_PTR5), .S(_02006_), .Z(_02111__PTR21) );
  MUX2_X1 U5441 ( .A(P1_P1_lWord_PTR6), .B(P1_EAX_PTR6), .S(_02006_), .Z(_02111__PTR22) );
  MUX2_X1 U5442 ( .A(P1_P1_lWord_PTR7), .B(P1_EAX_PTR7), .S(_02006_), .Z(_02111__PTR23) );
  MUX2_X1 U5443 ( .A(P1_P1_lWord_PTR8), .B(P1_EAX_PTR8), .S(_02006_), .Z(_02111__PTR24) );
  MUX2_X1 U5444 ( .A(P1_P1_lWord_PTR9), .B(P1_EAX_PTR9), .S(_02006_), .Z(_02111__PTR25) );
  MUX2_X1 U5445 ( .A(P1_P1_lWord_PTR10), .B(P1_EAX_PTR10), .S(_02006_), .Z(_02111__PTR26) );
  MUX2_X1 U5446 ( .A(P1_P1_lWord_PTR11), .B(P1_EAX_PTR11), .S(_02006_), .Z(_02111__PTR27) );
  MUX2_X1 U5447 ( .A(P1_P1_lWord_PTR12), .B(P1_EAX_PTR12), .S(_02006_), .Z(_02111__PTR28) );
  MUX2_X1 U5448 ( .A(P1_P1_lWord_PTR13), .B(P1_EAX_PTR13), .S(_02006_), .Z(_02111__PTR29) );
  MUX2_X1 U5449 ( .A(P1_P1_lWord_PTR14), .B(P1_EAX_PTR14), .S(_02006_), .Z(_02111__PTR30) );
  MUX2_X1 U5450 ( .A(P1_P1_lWord_PTR15), .B(P1_EAX_PTR15), .S(_02006_), .Z(_02111__PTR31) );
  MUX2_X1 U5451 ( .A(P1_P1_lWord_PTR0), .B(_02014__PTR0), .S(_02006_), .Z(_02111__PTR32) );
  MUX2_X1 U5452 ( .A(P1_P1_lWord_PTR1), .B(_02014__PTR1), .S(_02006_), .Z(_02111__PTR33) );
  MUX2_X1 U5453 ( .A(P1_P1_lWord_PTR2), .B(_02014__PTR2), .S(_02006_), .Z(_02111__PTR34) );
  MUX2_X1 U5454 ( .A(P1_P1_lWord_PTR3), .B(_02014__PTR3), .S(_02006_), .Z(_02111__PTR35) );
  MUX2_X1 U5455 ( .A(P1_P1_lWord_PTR4), .B(_02014__PTR4), .S(_02006_), .Z(_02111__PTR36) );
  MUX2_X1 U5456 ( .A(P1_P1_lWord_PTR5), .B(_02014__PTR5), .S(_02006_), .Z(_02111__PTR37) );
  MUX2_X1 U5457 ( .A(P1_P1_lWord_PTR6), .B(_02014__PTR6), .S(_02006_), .Z(_02111__PTR38) );
  MUX2_X1 U5458 ( .A(P1_P1_lWord_PTR7), .B(_02014__PTR7), .S(_02006_), .Z(_02111__PTR39) );
  MUX2_X1 U5459 ( .A(P1_P1_lWord_PTR8), .B(_02014__PTR8), .S(_02006_), .Z(_02111__PTR40) );
  MUX2_X1 U5460 ( .A(P1_P1_lWord_PTR9), .B(_02014__PTR9), .S(_02006_), .Z(_02111__PTR41) );
  MUX2_X1 U5461 ( .A(P1_P1_lWord_PTR10), .B(_02014__PTR10), .S(_02006_), .Z(_02111__PTR42) );
  MUX2_X1 U5462 ( .A(P1_P1_lWord_PTR11), .B(_02014__PTR11), .S(_02006_), .Z(_02111__PTR43) );
  MUX2_X1 U5463 ( .A(P1_P1_lWord_PTR12), .B(_02014__PTR12), .S(_02006_), .Z(_02111__PTR44) );
  MUX2_X1 U5464 ( .A(P1_P1_lWord_PTR13), .B(_02014__PTR13), .S(_02006_), .Z(_02111__PTR45) );
  MUX2_X1 U5465 ( .A(P1_P1_lWord_PTR14), .B(_02014__PTR14), .S(_02006_), .Z(_02111__PTR46) );
  MUX2_X1 U5466 ( .A(P1_P1_lWord_PTR15), .B(_02014__PTR15), .S(_02006_), .Z(_02111__PTR47) );
  MUX2_X1 U5467 ( .A(1'b0), .B(_02018_), .S(_02006_), .Z(_01853__PTR1) );
  MUX2_X1 U5468 ( .A(1'b1), .B(_02017_), .S(_02006_), .Z(_01857__PTR1) );
  MUX2_X1 U5469 ( .A(di1_PTR16), .B(P1_EAX_PTR16), .S(P1_READY_n), .Z(_02044__PTR16) );
  MUX2_X1 U5470 ( .A(di1_PTR17), .B(P1_EAX_PTR17), .S(P1_READY_n), .Z(_02044__PTR17) );
  MUX2_X1 U5471 ( .A(di1_PTR18), .B(P1_EAX_PTR18), .S(P1_READY_n), .Z(_02044__PTR18) );
  MUX2_X1 U5472 ( .A(di1_PTR19), .B(P1_EAX_PTR19), .S(P1_READY_n), .Z(_02044__PTR19) );
  MUX2_X1 U5473 ( .A(di1_PTR20), .B(P1_EAX_PTR20), .S(P1_READY_n), .Z(_02044__PTR20) );
  MUX2_X1 U5474 ( .A(di1_PTR21), .B(P1_EAX_PTR21), .S(P1_READY_n), .Z(_02044__PTR21) );
  MUX2_X1 U5475 ( .A(di1_PTR22), .B(P1_EAX_PTR22), .S(P1_READY_n), .Z(_02044__PTR22) );
  MUX2_X1 U5476 ( .A(di1_PTR23), .B(P1_EAX_PTR23), .S(P1_READY_n), .Z(_02044__PTR23) );
  MUX2_X1 U5477 ( .A(di1_PTR24), .B(P1_EAX_PTR24), .S(P1_READY_n), .Z(_02044__PTR24) );
  MUX2_X1 U5478 ( .A(di1_PTR25), .B(P1_EAX_PTR25), .S(P1_READY_n), .Z(_02044__PTR25) );
  MUX2_X1 U5479 ( .A(di1_PTR26), .B(P1_EAX_PTR26), .S(P1_READY_n), .Z(_02044__PTR26) );
  MUX2_X1 U5480 ( .A(di1_PTR27), .B(P1_EAX_PTR27), .S(P1_READY_n), .Z(_02044__PTR27) );
  MUX2_X1 U5481 ( .A(di1_PTR28), .B(P1_EAX_PTR28), .S(P1_READY_n), .Z(_02044__PTR28) );
  MUX2_X1 U5482 ( .A(di1_PTR29), .B(P1_EAX_PTR29), .S(P1_READY_n), .Z(_02044__PTR29) );
  MUX2_X1 U5483 ( .A(di1_PTR30), .B(P1_EAX_PTR30), .S(P1_READY_n), .Z(_02044__PTR30) );
  MUX2_X1 U5484 ( .A(P1_Datai_PTR31), .B(P1_EAX_PTR31), .S(P1_READY_n), .Z(_02044__PTR31) );
  MUX2_X1 U5485 ( .A(di1_PTR0), .B(P1_EAX_PTR0), .S(P1_READY_n), .Z(_02016__PTR0) );
  MUX2_X1 U5486 ( .A(di1_PTR1), .B(P1_EAX_PTR1), .S(P1_READY_n), .Z(_02016__PTR1) );
  MUX2_X1 U5487 ( .A(di1_PTR2), .B(P1_EAX_PTR2), .S(P1_READY_n), .Z(_02016__PTR2) );
  MUX2_X1 U5488 ( .A(di1_PTR3), .B(P1_EAX_PTR3), .S(P1_READY_n), .Z(_02016__PTR3) );
  MUX2_X1 U5489 ( .A(di1_PTR4), .B(P1_EAX_PTR4), .S(P1_READY_n), .Z(_02016__PTR4) );
  MUX2_X1 U5490 ( .A(di1_PTR5), .B(P1_EAX_PTR5), .S(P1_READY_n), .Z(_02016__PTR5) );
  MUX2_X1 U5491 ( .A(di1_PTR6), .B(P1_EAX_PTR6), .S(P1_READY_n), .Z(_02016__PTR6) );
  MUX2_X1 U5492 ( .A(di1_PTR7), .B(P1_EAX_PTR7), .S(P1_READY_n), .Z(_02016__PTR7) );
  MUX2_X1 U5493 ( .A(di1_PTR8), .B(P1_EAX_PTR8), .S(P1_READY_n), .Z(_02016__PTR8) );
  MUX2_X1 U5494 ( .A(di1_PTR9), .B(P1_EAX_PTR9), .S(P1_READY_n), .Z(_02016__PTR9) );
  MUX2_X1 U5495 ( .A(di1_PTR10), .B(P1_EAX_PTR10), .S(P1_READY_n), .Z(_02016__PTR10) );
  MUX2_X1 U5496 ( .A(di1_PTR11), .B(P1_EAX_PTR11), .S(P1_READY_n), .Z(_02016__PTR11) );
  MUX2_X1 U5497 ( .A(di1_PTR12), .B(P1_EAX_PTR12), .S(P1_READY_n), .Z(_02016__PTR12) );
  MUX2_X1 U5498 ( .A(di1_PTR13), .B(P1_EAX_PTR13), .S(P1_READY_n), .Z(_02016__PTR13) );
  MUX2_X1 U5499 ( .A(di1_PTR14), .B(P1_EAX_PTR14), .S(P1_READY_n), .Z(_02016__PTR14) );
  MUX2_X1 U5500 ( .A(di1_PTR15), .B(P1_EAX_PTR15), .S(P1_READY_n), .Z(_02016__PTR15) );
  MUX2_X1 U5501 ( .A(di1_PTR0), .B(P1_EAX_PTR16), .S(P1_READY_n), .Z(_02016__PTR16) );
  MUX2_X1 U5502 ( .A(di1_PTR1), .B(P1_EAX_PTR17), .S(P1_READY_n), .Z(_02016__PTR17) );
  MUX2_X1 U5503 ( .A(di1_PTR2), .B(P1_EAX_PTR18), .S(P1_READY_n), .Z(_02016__PTR18) );
  MUX2_X1 U5504 ( .A(di1_PTR3), .B(P1_EAX_PTR19), .S(P1_READY_n), .Z(_02016__PTR19) );
  MUX2_X1 U5505 ( .A(di1_PTR4), .B(P1_EAX_PTR20), .S(P1_READY_n), .Z(_02016__PTR20) );
  MUX2_X1 U5506 ( .A(di1_PTR5), .B(P1_EAX_PTR21), .S(P1_READY_n), .Z(_02016__PTR21) );
  MUX2_X1 U5507 ( .A(di1_PTR6), .B(P1_EAX_PTR22), .S(P1_READY_n), .Z(_02016__PTR22) );
  MUX2_X1 U5508 ( .A(di1_PTR7), .B(P1_EAX_PTR23), .S(P1_READY_n), .Z(_02016__PTR23) );
  MUX2_X1 U5509 ( .A(di1_PTR8), .B(P1_EAX_PTR24), .S(P1_READY_n), .Z(_02016__PTR24) );
  MUX2_X1 U5510 ( .A(di1_PTR9), .B(P1_EAX_PTR25), .S(P1_READY_n), .Z(_02016__PTR25) );
  MUX2_X1 U5511 ( .A(di1_PTR10), .B(P1_EAX_PTR26), .S(P1_READY_n), .Z(_02016__PTR26) );
  MUX2_X1 U5512 ( .A(di1_PTR11), .B(P1_EAX_PTR27), .S(P1_READY_n), .Z(_02016__PTR27) );
  MUX2_X1 U5513 ( .A(di1_PTR12), .B(P1_EAX_PTR28), .S(P1_READY_n), .Z(_02016__PTR28) );
  MUX2_X1 U5514 ( .A(di1_PTR13), .B(P1_EAX_PTR29), .S(P1_READY_n), .Z(_02016__PTR29) );
  MUX2_X1 U5515 ( .A(di1_PTR14), .B(P1_EAX_PTR30), .S(P1_READY_n), .Z(_02016__PTR30) );
  MUX2_X1 U5516 ( .A(1'b0), .B(P1_EAX_PTR31), .S(P1_READY_n), .Z(_02016__PTR31) );
  MUX2_X1 U5517 ( .A(P1_P1_uWord_PTR0), .B(_02825__PTR0), .S(_02006_), .Z(_02107__PTR15) );
  MUX2_X1 U5518 ( .A(P1_P1_uWord_PTR1), .B(_02826__PTR1), .S(_02006_), .Z(_02107__PTR16) );
  MUX2_X1 U5519 ( .A(P1_P1_uWord_PTR2), .B(_02826__PTR2), .S(_02006_), .Z(_02107__PTR17) );
  MUX2_X1 U5520 ( .A(P1_P1_uWord_PTR3), .B(_02826__PTR3), .S(_02006_), .Z(_02107__PTR18) );
  MUX2_X1 U5521 ( .A(P1_P1_uWord_PTR4), .B(_02826__PTR4), .S(_02006_), .Z(_02107__PTR19) );
  MUX2_X1 U5522 ( .A(P1_P1_uWord_PTR5), .B(_02826__PTR5), .S(_02006_), .Z(_02107__PTR20) );
  MUX2_X1 U5523 ( .A(P1_P1_uWord_PTR6), .B(_02826__PTR6), .S(_02006_), .Z(_02107__PTR21) );
  MUX2_X1 U5524 ( .A(P1_P1_uWord_PTR7), .B(_02826__PTR7), .S(_02006_), .Z(_02107__PTR22) );
  MUX2_X1 U5525 ( .A(P1_P1_uWord_PTR8), .B(_02826__PTR8), .S(_02006_), .Z(_02107__PTR23) );
  MUX2_X1 U5526 ( .A(P1_P1_uWord_PTR9), .B(_02826__PTR9), .S(_02006_), .Z(_02107__PTR24) );
  MUX2_X1 U5527 ( .A(P1_P1_uWord_PTR10), .B(_02826__PTR10), .S(_02006_), .Z(_02107__PTR25) );
  MUX2_X1 U5528 ( .A(P1_P1_uWord_PTR11), .B(_02826__PTR11), .S(_02006_), .Z(_02107__PTR26) );
  MUX2_X1 U5529 ( .A(P1_P1_uWord_PTR12), .B(_02826__PTR12), .S(_02006_), .Z(_02107__PTR27) );
  MUX2_X1 U5530 ( .A(P1_P1_uWord_PTR13), .B(_02826__PTR13), .S(_02006_), .Z(_02107__PTR28) );
  MUX2_X1 U5531 ( .A(P1_P1_uWord_PTR14), .B(_02826__PTR14), .S(_02006_), .Z(_02107__PTR29) );
  MUX2_X1 U5532 ( .A(P1_P1_uWord_PTR0), .B(_02013__PTR0), .S(_02006_), .Z(_02107__PTR30) );
  MUX2_X1 U5533 ( .A(P1_P1_uWord_PTR1), .B(_02013__PTR1), .S(_02006_), .Z(_02107__PTR31) );
  MUX2_X1 U5534 ( .A(P1_P1_uWord_PTR2), .B(_02013__PTR2), .S(_02006_), .Z(_02107__PTR32) );
  MUX2_X1 U5535 ( .A(P1_P1_uWord_PTR3), .B(_02013__PTR3), .S(_02006_), .Z(_02107__PTR33) );
  MUX2_X1 U5536 ( .A(P1_P1_uWord_PTR4), .B(_02013__PTR4), .S(_02006_), .Z(_02107__PTR34) );
  MUX2_X1 U5537 ( .A(P1_P1_uWord_PTR5), .B(_02013__PTR5), .S(_02006_), .Z(_02107__PTR35) );
  MUX2_X1 U5538 ( .A(P1_P1_uWord_PTR6), .B(_02013__PTR6), .S(_02006_), .Z(_02107__PTR36) );
  MUX2_X1 U5539 ( .A(P1_P1_uWord_PTR7), .B(_02013__PTR7), .S(_02006_), .Z(_02107__PTR37) );
  MUX2_X1 U5540 ( .A(P1_P1_uWord_PTR8), .B(_02013__PTR8), .S(_02006_), .Z(_02107__PTR38) );
  MUX2_X1 U5541 ( .A(P1_P1_uWord_PTR9), .B(_02013__PTR9), .S(_02006_), .Z(_02107__PTR39) );
  MUX2_X1 U5542 ( .A(P1_P1_uWord_PTR10), .B(_02013__PTR10), .S(_02006_), .Z(_02107__PTR40) );
  MUX2_X1 U5543 ( .A(P1_P1_uWord_PTR11), .B(_02013__PTR11), .S(_02006_), .Z(_02107__PTR41) );
  MUX2_X1 U5544 ( .A(P1_P1_uWord_PTR12), .B(_02013__PTR12), .S(_02006_), .Z(_02107__PTR42) );
  MUX2_X1 U5545 ( .A(P1_P1_uWord_PTR13), .B(_02013__PTR13), .S(_02006_), .Z(_02107__PTR43) );
  MUX2_X1 U5546 ( .A(P1_P1_uWord_PTR14), .B(_02013__PTR14), .S(_02006_), .Z(_02107__PTR44) );
  MUX2_X1 U5547 ( .A(P1_CodeFetch), .B(1'b0), .S(_02006_), .Z(_01872__PTR0) );
  MUX2_X1 U5548 ( .A(P1_MemoryFetch), .B(1'b1), .S(_02006_), .Z(_01868__PTR1) );
  MUX2_X1 U5549 ( .A(P1_ReadRequest), .B(1'b1), .S(_02006_), .Z(_01865__PTR1) );
  MUX2_X1 U5550 ( .A(P1_RequestPending), .B(P1_READY_n), .S(_02006_), .Z(_01861__PTR1) );
  MUX2_X1 U5551 ( .A(P1_P1_InstQueueRd_Addr_PTR4), .B(_02045__PTR4), .S(_02006_), .Z(_02088__PTR19) );
  MUX2_X1 U5552 ( .A(P1_P1_InstQueueRd_Addr_PTR1), .B(_02038__PTR1), .S(_02006_), .Z(_02088__PTR11) );
  MUX2_X1 U5553 ( .A(P1_P1_InstQueueRd_Addr_PTR2), .B(_02038__PTR2), .S(_02006_), .Z(_02088__PTR12) );
  MUX2_X1 U5554 ( .A(P1_P1_InstQueueRd_Addr_PTR3), .B(_02038__PTR3), .S(_02006_), .Z(_02088__PTR13) );
  MUX2_X1 U5555 ( .A(P1_P1_InstQueueRd_Addr_PTR4), .B(_02038__PTR4), .S(_02006_), .Z(_02088__PTR14) );
  MUX2_X1 U5556 ( .A(P1_P1_InstQueueRd_Addr_PTR1), .B(_02020__PTR1), .S(_02006_), .Z(_02088__PTR21) );
  MUX2_X1 U5557 ( .A(P1_P1_InstQueueRd_Addr_PTR2), .B(_02020__PTR2), .S(_02006_), .Z(_02088__PTR22) );
  MUX2_X1 U5558 ( .A(P1_P1_InstQueueRd_Addr_PTR3), .B(_02020__PTR3), .S(_02006_), .Z(_02088__PTR23) );
  MUX2_X1 U5559 ( .A(P1_P1_InstQueueRd_Addr_PTR4), .B(_02020__PTR4), .S(_02006_), .Z(_02088__PTR24) );
  MUX2_X1 U5560 ( .A(_02084__PTR33), .B(P1_P1_InstAddrPointer_PTR1), .S(P1_READY_n), .Z(_02019__PTR1) );
  MUX2_X1 U5561 ( .A(_02084__PTR34), .B(P1_P1_InstAddrPointer_PTR2), .S(P1_READY_n), .Z(_02019__PTR2) );
  MUX2_X1 U5562 ( .A(_02084__PTR35), .B(P1_P1_InstAddrPointer_PTR3), .S(P1_READY_n), .Z(_02019__PTR3) );
  MUX2_X1 U5563 ( .A(_02084__PTR36), .B(P1_P1_InstAddrPointer_PTR4), .S(P1_READY_n), .Z(_02019__PTR4) );
  MUX2_X1 U5564 ( .A(_02084__PTR37), .B(P1_P1_InstAddrPointer_PTR5), .S(P1_READY_n), .Z(_02019__PTR5) );
  MUX2_X1 U5565 ( .A(_02084__PTR38), .B(P1_P1_InstAddrPointer_PTR6), .S(P1_READY_n), .Z(_02019__PTR6) );
  MUX2_X1 U5566 ( .A(_02084__PTR39), .B(P1_P1_InstAddrPointer_PTR7), .S(P1_READY_n), .Z(_02019__PTR7) );
  MUX2_X1 U5567 ( .A(_02084__PTR40), .B(P1_P1_InstAddrPointer_PTR8), .S(P1_READY_n), .Z(_02019__PTR8) );
  MUX2_X1 U5568 ( .A(_02084__PTR41), .B(P1_P1_InstAddrPointer_PTR9), .S(P1_READY_n), .Z(_02019__PTR9) );
  MUX2_X1 U5569 ( .A(_02084__PTR42), .B(P1_P1_InstAddrPointer_PTR10), .S(P1_READY_n), .Z(_02019__PTR10) );
  MUX2_X1 U5570 ( .A(_02084__PTR43), .B(P1_P1_InstAddrPointer_PTR11), .S(P1_READY_n), .Z(_02019__PTR11) );
  MUX2_X1 U5571 ( .A(_02084__PTR44), .B(P1_P1_InstAddrPointer_PTR12), .S(P1_READY_n), .Z(_02019__PTR12) );
  MUX2_X1 U5572 ( .A(_02084__PTR45), .B(P1_P1_InstAddrPointer_PTR13), .S(P1_READY_n), .Z(_02019__PTR13) );
  MUX2_X1 U5573 ( .A(_02084__PTR46), .B(P1_P1_InstAddrPointer_PTR14), .S(P1_READY_n), .Z(_02019__PTR14) );
  MUX2_X1 U5574 ( .A(_02084__PTR47), .B(P1_P1_InstAddrPointer_PTR15), .S(P1_READY_n), .Z(_02019__PTR15) );
  MUX2_X1 U5575 ( .A(_02084__PTR48), .B(P1_P1_InstAddrPointer_PTR16), .S(P1_READY_n), .Z(_02019__PTR16) );
  MUX2_X1 U5576 ( .A(_02084__PTR49), .B(P1_P1_InstAddrPointer_PTR17), .S(P1_READY_n), .Z(_02019__PTR17) );
  MUX2_X1 U5577 ( .A(_02084__PTR50), .B(P1_P1_InstAddrPointer_PTR18), .S(P1_READY_n), .Z(_02019__PTR18) );
  MUX2_X1 U5578 ( .A(_02084__PTR51), .B(P1_P1_InstAddrPointer_PTR19), .S(P1_READY_n), .Z(_02019__PTR19) );
  MUX2_X1 U5579 ( .A(_02084__PTR52), .B(P1_P1_InstAddrPointer_PTR20), .S(P1_READY_n), .Z(_02019__PTR20) );
  MUX2_X1 U5580 ( .A(_02084__PTR53), .B(P1_P1_InstAddrPointer_PTR21), .S(P1_READY_n), .Z(_02019__PTR21) );
  MUX2_X1 U5581 ( .A(_02084__PTR54), .B(P1_P1_InstAddrPointer_PTR22), .S(P1_READY_n), .Z(_02019__PTR22) );
  MUX2_X1 U5582 ( .A(_02084__PTR55), .B(P1_P1_InstAddrPointer_PTR23), .S(P1_READY_n), .Z(_02019__PTR23) );
  MUX2_X1 U5583 ( .A(_02084__PTR56), .B(P1_P1_InstAddrPointer_PTR24), .S(P1_READY_n), .Z(_02019__PTR24) );
  MUX2_X1 U5584 ( .A(_02084__PTR57), .B(P1_P1_InstAddrPointer_PTR25), .S(P1_READY_n), .Z(_02019__PTR25) );
  MUX2_X1 U5585 ( .A(_02084__PTR58), .B(P1_P1_InstAddrPointer_PTR26), .S(P1_READY_n), .Z(_02019__PTR26) );
  MUX2_X1 U5586 ( .A(_02084__PTR59), .B(P1_P1_InstAddrPointer_PTR27), .S(P1_READY_n), .Z(_02019__PTR27) );
  MUX2_X1 U5587 ( .A(_02084__PTR60), .B(P1_P1_InstAddrPointer_PTR28), .S(P1_READY_n), .Z(_02019__PTR28) );
  MUX2_X1 U5588 ( .A(_02084__PTR61), .B(P1_P1_InstAddrPointer_PTR29), .S(P1_READY_n), .Z(_02019__PTR29) );
  MUX2_X1 U5589 ( .A(_02084__PTR62), .B(P1_P1_InstAddrPointer_PTR30), .S(P1_READY_n), .Z(_02019__PTR30) );
  MUX2_X1 U5590 ( .A(_02084__PTR63), .B(P1_P1_InstAddrPointer_PTR31), .S(P1_READY_n), .Z(_02019__PTR31) );
  MUX2_X1 U5591 ( .A(1'b0), .B(P1_P1_Flush), .S(P1_READY_n), .Z(_02018_) );
  MUX2_X1 U5592 ( .A(1'b0), .B(P1_P1_More), .S(P1_READY_n), .Z(_02017_) );
  MUX2_X1 U5593 ( .A(_02010__PTR0), .B(P1_EBX_PTR0), .S(P1_READY_n), .Z(_02015__PTR0) );
  MUX2_X1 U5594 ( .A(_02010__PTR1), .B(_02009__PTR1), .S(P1_READY_n), .Z(_02015__PTR1) );
  MUX2_X1 U5595 ( .A(_02010__PTR2), .B(_02009__PTR2), .S(P1_READY_n), .Z(_02015__PTR2) );
  MUX2_X1 U5596 ( .A(_02010__PTR3), .B(_02009__PTR3), .S(P1_READY_n), .Z(_02015__PTR3) );
  MUX2_X1 U5597 ( .A(_02010__PTR4), .B(_02009__PTR4), .S(P1_READY_n), .Z(_02015__PTR4) );
  MUX2_X1 U5598 ( .A(_02010__PTR5), .B(_02009__PTR5), .S(P1_READY_n), .Z(_02015__PTR5) );
  MUX2_X1 U5599 ( .A(_02010__PTR6), .B(_02009__PTR6), .S(P1_READY_n), .Z(_02015__PTR6) );
  MUX2_X1 U5600 ( .A(_02010__PTR7), .B(_02009__PTR7), .S(P1_READY_n), .Z(_02015__PTR7) );
  MUX2_X1 U5601 ( .A(_02010__PTR8), .B(_02009__PTR8), .S(P1_READY_n), .Z(_02015__PTR8) );
  MUX2_X1 U5602 ( .A(_02010__PTR9), .B(_02009__PTR9), .S(P1_READY_n), .Z(_02015__PTR9) );
  MUX2_X1 U5603 ( .A(_02010__PTR10), .B(_02009__PTR10), .S(P1_READY_n), .Z(_02015__PTR10) );
  MUX2_X1 U5604 ( .A(_02010__PTR11), .B(_02009__PTR11), .S(P1_READY_n), .Z(_02015__PTR11) );
  MUX2_X1 U5605 ( .A(_02010__PTR12), .B(_02009__PTR12), .S(P1_READY_n), .Z(_02015__PTR12) );
  MUX2_X1 U5606 ( .A(_02010__PTR13), .B(_02009__PTR13), .S(P1_READY_n), .Z(_02015__PTR13) );
  MUX2_X1 U5607 ( .A(_02010__PTR14), .B(_02009__PTR14), .S(P1_READY_n), .Z(_02015__PTR14) );
  MUX2_X1 U5608 ( .A(_02010__PTR15), .B(_02009__PTR15), .S(P1_READY_n), .Z(_02015__PTR15) );
  MUX2_X1 U5609 ( .A(_02010__PTR16), .B(_02009__PTR16), .S(P1_READY_n), .Z(_02015__PTR16) );
  MUX2_X1 U5610 ( .A(_02010__PTR17), .B(_02009__PTR17), .S(P1_READY_n), .Z(_02015__PTR17) );
  MUX2_X1 U5611 ( .A(_02010__PTR18), .B(_02009__PTR18), .S(P1_READY_n), .Z(_02015__PTR18) );
  MUX2_X1 U5612 ( .A(_02010__PTR19), .B(_02009__PTR19), .S(P1_READY_n), .Z(_02015__PTR19) );
  MUX2_X1 U5613 ( .A(_02010__PTR20), .B(_02009__PTR20), .S(P1_READY_n), .Z(_02015__PTR20) );
  MUX2_X1 U5614 ( .A(_02010__PTR21), .B(_02009__PTR21), .S(P1_READY_n), .Z(_02015__PTR21) );
  MUX2_X1 U5615 ( .A(_02010__PTR22), .B(_02009__PTR22), .S(P1_READY_n), .Z(_02015__PTR22) );
  MUX2_X1 U5616 ( .A(_02010__PTR23), .B(_02009__PTR23), .S(P1_READY_n), .Z(_02015__PTR23) );
  MUX2_X1 U5617 ( .A(_02010__PTR24), .B(_02009__PTR24), .S(P1_READY_n), .Z(_02015__PTR24) );
  MUX2_X1 U5618 ( .A(_02010__PTR25), .B(_02009__PTR25), .S(P1_READY_n), .Z(_02015__PTR25) );
  MUX2_X1 U5619 ( .A(_02010__PTR26), .B(_02009__PTR26), .S(P1_READY_n), .Z(_02015__PTR26) );
  MUX2_X1 U5620 ( .A(_02010__PTR27), .B(_02009__PTR27), .S(P1_READY_n), .Z(_02015__PTR27) );
  MUX2_X1 U5621 ( .A(_02010__PTR28), .B(_02009__PTR28), .S(P1_READY_n), .Z(_02015__PTR28) );
  MUX2_X1 U5622 ( .A(_02010__PTR29), .B(_02009__PTR29), .S(P1_READY_n), .Z(_02015__PTR29) );
  MUX2_X1 U5623 ( .A(_02010__PTR30), .B(_02009__PTR30), .S(P1_READY_n), .Z(_02015__PTR30) );
  MUX2_X1 U5624 ( .A(_02010__PTR31), .B(_02009__PTR31), .S(P1_READY_n), .Z(_02015__PTR31) );
  MUX2_X1 U5625 ( .A(di1_PTR0), .B(P1_P1_lWord_PTR0), .S(P1_READY_n), .Z(_02014__PTR0) );
  MUX2_X1 U5626 ( .A(di1_PTR1), .B(P1_P1_lWord_PTR1), .S(P1_READY_n), .Z(_02014__PTR1) );
  MUX2_X1 U5627 ( .A(di1_PTR2), .B(P1_P1_lWord_PTR2), .S(P1_READY_n), .Z(_02014__PTR2) );
  MUX2_X1 U5628 ( .A(di1_PTR3), .B(P1_P1_lWord_PTR3), .S(P1_READY_n), .Z(_02014__PTR3) );
  MUX2_X1 U5629 ( .A(di1_PTR4), .B(P1_P1_lWord_PTR4), .S(P1_READY_n), .Z(_02014__PTR4) );
  MUX2_X1 U5630 ( .A(di1_PTR5), .B(P1_P1_lWord_PTR5), .S(P1_READY_n), .Z(_02014__PTR5) );
  MUX2_X1 U5631 ( .A(di1_PTR6), .B(P1_P1_lWord_PTR6), .S(P1_READY_n), .Z(_02014__PTR6) );
  MUX2_X1 U5632 ( .A(di1_PTR7), .B(P1_P1_lWord_PTR7), .S(P1_READY_n), .Z(_02014__PTR7) );
  MUX2_X1 U5633 ( .A(di1_PTR8), .B(P1_P1_lWord_PTR8), .S(P1_READY_n), .Z(_02014__PTR8) );
  MUX2_X1 U5634 ( .A(di1_PTR9), .B(P1_P1_lWord_PTR9), .S(P1_READY_n), .Z(_02014__PTR9) );
  MUX2_X1 U5635 ( .A(di1_PTR10), .B(P1_P1_lWord_PTR10), .S(P1_READY_n), .Z(_02014__PTR10) );
  MUX2_X1 U5636 ( .A(di1_PTR11), .B(P1_P1_lWord_PTR11), .S(P1_READY_n), .Z(_02014__PTR11) );
  MUX2_X1 U5637 ( .A(di1_PTR12), .B(P1_P1_lWord_PTR12), .S(P1_READY_n), .Z(_02014__PTR12) );
  MUX2_X1 U5638 ( .A(di1_PTR13), .B(P1_P1_lWord_PTR13), .S(P1_READY_n), .Z(_02014__PTR13) );
  MUX2_X1 U5639 ( .A(di1_PTR14), .B(P1_P1_lWord_PTR14), .S(P1_READY_n), .Z(_02014__PTR14) );
  MUX2_X1 U5640 ( .A(di1_PTR15), .B(P1_P1_lWord_PTR15), .S(P1_READY_n), .Z(_02014__PTR15) );
  MUX2_X1 U5641 ( .A(di1_PTR0), .B(P1_P1_uWord_PTR0), .S(P1_READY_n), .Z(_02013__PTR0) );
  MUX2_X1 U5642 ( .A(di1_PTR1), .B(P1_P1_uWord_PTR1), .S(P1_READY_n), .Z(_02013__PTR1) );
  MUX2_X1 U5643 ( .A(di1_PTR2), .B(P1_P1_uWord_PTR2), .S(P1_READY_n), .Z(_02013__PTR2) );
  MUX2_X1 U5644 ( .A(di1_PTR3), .B(P1_P1_uWord_PTR3), .S(P1_READY_n), .Z(_02013__PTR3) );
  MUX2_X1 U5645 ( .A(di1_PTR4), .B(P1_P1_uWord_PTR4), .S(P1_READY_n), .Z(_02013__PTR4) );
  MUX2_X1 U5646 ( .A(di1_PTR5), .B(P1_P1_uWord_PTR5), .S(P1_READY_n), .Z(_02013__PTR5) );
  MUX2_X1 U5647 ( .A(di1_PTR6), .B(P1_P1_uWord_PTR6), .S(P1_READY_n), .Z(_02013__PTR6) );
  MUX2_X1 U5648 ( .A(di1_PTR7), .B(P1_P1_uWord_PTR7), .S(P1_READY_n), .Z(_02013__PTR7) );
  MUX2_X1 U5649 ( .A(di1_PTR8), .B(P1_P1_uWord_PTR8), .S(P1_READY_n), .Z(_02013__PTR8) );
  MUX2_X1 U5650 ( .A(di1_PTR9), .B(P1_P1_uWord_PTR9), .S(P1_READY_n), .Z(_02013__PTR9) );
  MUX2_X1 U5651 ( .A(di1_PTR10), .B(P1_P1_uWord_PTR10), .S(P1_READY_n), .Z(_02013__PTR10) );
  MUX2_X1 U5652 ( .A(di1_PTR11), .B(P1_P1_uWord_PTR11), .S(P1_READY_n), .Z(_02013__PTR11) );
  MUX2_X1 U5653 ( .A(di1_PTR12), .B(P1_P1_uWord_PTR12), .S(P1_READY_n), .Z(_02013__PTR12) );
  MUX2_X1 U5654 ( .A(di1_PTR13), .B(P1_P1_uWord_PTR13), .S(P1_READY_n), .Z(_02013__PTR13) );
  MUX2_X1 U5655 ( .A(di1_PTR14), .B(P1_P1_uWord_PTR14), .S(P1_READY_n), .Z(_02013__PTR14) );
  MUX2_X1 U5656 ( .A(P1_P1_InstAddrPointer_PTR0), .B(_02084__PTR0), .S(_01853__PTR2), .Z(_02084__PTR128) );
  MUX2_X1 U5657 ( .A(P1_P1_InstAddrPointer_PTR1), .B(_02084__PTR1), .S(_01853__PTR2), .Z(_02084__PTR129) );
  MUX2_X1 U5658 ( .A(P1_P1_InstAddrPointer_PTR2), .B(_02807__PTR2), .S(_01853__PTR2), .Z(_02084__PTR130) );
  MUX2_X1 U5659 ( .A(P1_P1_InstAddrPointer_PTR3), .B(_02807__PTR3), .S(_01853__PTR2), .Z(_02084__PTR131) );
  MUX2_X1 U5660 ( .A(P1_P1_InstAddrPointer_PTR4), .B(_02807__PTR4), .S(_01853__PTR2), .Z(_02084__PTR132) );
  MUX2_X1 U5661 ( .A(P1_P1_InstAddrPointer_PTR5), .B(_02807__PTR5), .S(_01853__PTR2), .Z(_02084__PTR133) );
  MUX2_X1 U5662 ( .A(P1_P1_InstAddrPointer_PTR6), .B(_02807__PTR6), .S(_01853__PTR2), .Z(_02084__PTR134) );
  MUX2_X1 U5663 ( .A(P1_P1_InstAddrPointer_PTR7), .B(_02807__PTR7), .S(_01853__PTR2), .Z(_02084__PTR135) );
  MUX2_X1 U5664 ( .A(P1_P1_InstAddrPointer_PTR8), .B(_02807__PTR8), .S(_01853__PTR2), .Z(_02084__PTR136) );
  MUX2_X1 U5665 ( .A(P1_P1_InstAddrPointer_PTR9), .B(_02807__PTR9), .S(_01853__PTR2), .Z(_02084__PTR137) );
  MUX2_X1 U5666 ( .A(P1_P1_InstAddrPointer_PTR10), .B(_02807__PTR10), .S(_01853__PTR2), .Z(_02084__PTR138) );
  MUX2_X1 U5667 ( .A(P1_P1_InstAddrPointer_PTR11), .B(_02807__PTR11), .S(_01853__PTR2), .Z(_02084__PTR139) );
  MUX2_X1 U5668 ( .A(P1_P1_InstAddrPointer_PTR12), .B(_02807__PTR12), .S(_01853__PTR2), .Z(_02084__PTR140) );
  MUX2_X1 U5669 ( .A(P1_P1_InstAddrPointer_PTR13), .B(_02807__PTR13), .S(_01853__PTR2), .Z(_02084__PTR141) );
  MUX2_X1 U5670 ( .A(P1_P1_InstAddrPointer_PTR14), .B(_02807__PTR14), .S(_01853__PTR2), .Z(_02084__PTR142) );
  MUX2_X1 U5671 ( .A(P1_P1_InstAddrPointer_PTR15), .B(_02807__PTR15), .S(_01853__PTR2), .Z(_02084__PTR143) );
  MUX2_X1 U5672 ( .A(P1_P1_InstAddrPointer_PTR16), .B(_02807__PTR16), .S(_01853__PTR2), .Z(_02084__PTR144) );
  MUX2_X1 U5673 ( .A(P1_P1_InstAddrPointer_PTR17), .B(_02807__PTR17), .S(_01853__PTR2), .Z(_02084__PTR145) );
  MUX2_X1 U5674 ( .A(P1_P1_InstAddrPointer_PTR18), .B(_02807__PTR18), .S(_01853__PTR2), .Z(_02084__PTR146) );
  MUX2_X1 U5675 ( .A(P1_P1_InstAddrPointer_PTR19), .B(_02807__PTR19), .S(_01853__PTR2), .Z(_02084__PTR147) );
  MUX2_X1 U5676 ( .A(P1_P1_InstAddrPointer_PTR20), .B(_02807__PTR20), .S(_01853__PTR2), .Z(_02084__PTR148) );
  MUX2_X1 U5677 ( .A(P1_P1_InstAddrPointer_PTR21), .B(_02807__PTR21), .S(_01853__PTR2), .Z(_02084__PTR149) );
  MUX2_X1 U5678 ( .A(P1_P1_InstAddrPointer_PTR22), .B(_02807__PTR22), .S(_01853__PTR2), .Z(_02084__PTR150) );
  MUX2_X1 U5679 ( .A(P1_P1_InstAddrPointer_PTR23), .B(_02807__PTR23), .S(_01853__PTR2), .Z(_02084__PTR151) );
  MUX2_X1 U5680 ( .A(P1_P1_InstAddrPointer_PTR24), .B(_02807__PTR24), .S(_01853__PTR2), .Z(_02084__PTR152) );
  MUX2_X1 U5681 ( .A(P1_P1_InstAddrPointer_PTR25), .B(_02807__PTR25), .S(_01853__PTR2), .Z(_02084__PTR153) );
  MUX2_X1 U5682 ( .A(P1_P1_InstAddrPointer_PTR26), .B(_02807__PTR26), .S(_01853__PTR2), .Z(_02084__PTR154) );
  MUX2_X1 U5683 ( .A(P1_P1_InstAddrPointer_PTR27), .B(_02807__PTR27), .S(_01853__PTR2), .Z(_02084__PTR155) );
  MUX2_X1 U5684 ( .A(P1_P1_InstAddrPointer_PTR28), .B(_02807__PTR28), .S(_01853__PTR2), .Z(_02084__PTR156) );
  MUX2_X1 U5685 ( .A(P1_P1_InstAddrPointer_PTR29), .B(_02807__PTR29), .S(_01853__PTR2), .Z(_02084__PTR157) );
  MUX2_X1 U5686 ( .A(P1_P1_InstAddrPointer_PTR30), .B(_02807__PTR30), .S(_01853__PTR2), .Z(_02084__PTR158) );
  MUX2_X1 U5687 ( .A(P1_P1_InstAddrPointer_PTR31), .B(_02807__PTR31), .S(_01853__PTR2), .Z(_02084__PTR159) );
  MUX2_X1 U5688 ( .A(P1_P1_InstAddrPointer_PTR0), .B(_02809__PTR0), .S(_01853__PTR2), .Z(_02084__PTR160) );
  MUX2_X1 U5689 ( .A(P1_P1_InstAddrPointer_PTR1), .B(_02810__PTR1), .S(_01853__PTR2), .Z(_02084__PTR161) );
  MUX2_X1 U5690 ( .A(P1_P1_InstAddrPointer_PTR2), .B(_02810__PTR2), .S(_01853__PTR2), .Z(_02084__PTR162) );
  MUX2_X1 U5691 ( .A(P1_P1_InstAddrPointer_PTR3), .B(_02810__PTR3), .S(_01853__PTR2), .Z(_02084__PTR163) );
  MUX2_X1 U5692 ( .A(P1_P1_InstAddrPointer_PTR4), .B(_02810__PTR4), .S(_01853__PTR2), .Z(_02084__PTR164) );
  MUX2_X1 U5693 ( .A(P1_P1_InstAddrPointer_PTR5), .B(_02810__PTR5), .S(_01853__PTR2), .Z(_02084__PTR165) );
  MUX2_X1 U5694 ( .A(P1_P1_InstAddrPointer_PTR6), .B(_02810__PTR6), .S(_01853__PTR2), .Z(_02084__PTR166) );
  MUX2_X1 U5695 ( .A(P1_P1_InstAddrPointer_PTR7), .B(_02810__PTR7), .S(_01853__PTR2), .Z(_02084__PTR167) );
  MUX2_X1 U5696 ( .A(P1_P1_InstAddrPointer_PTR8), .B(_02810__PTR8), .S(_01853__PTR2), .Z(_02084__PTR168) );
  MUX2_X1 U5697 ( .A(P1_P1_InstAddrPointer_PTR9), .B(_02810__PTR9), .S(_01853__PTR2), .Z(_02084__PTR169) );
  MUX2_X1 U5698 ( .A(P1_P1_InstAddrPointer_PTR10), .B(_02810__PTR10), .S(_01853__PTR2), .Z(_02084__PTR170) );
  MUX2_X1 U5699 ( .A(P1_P1_InstAddrPointer_PTR11), .B(_02810__PTR11), .S(_01853__PTR2), .Z(_02084__PTR171) );
  MUX2_X1 U5700 ( .A(P1_P1_InstAddrPointer_PTR12), .B(_02810__PTR12), .S(_01853__PTR2), .Z(_02084__PTR172) );
  MUX2_X1 U5701 ( .A(P1_P1_InstAddrPointer_PTR13), .B(_02810__PTR13), .S(_01853__PTR2), .Z(_02084__PTR173) );
  MUX2_X1 U5702 ( .A(P1_P1_InstAddrPointer_PTR14), .B(_02810__PTR14), .S(_01853__PTR2), .Z(_02084__PTR174) );
  MUX2_X1 U5703 ( .A(P1_P1_InstAddrPointer_PTR15), .B(_02810__PTR15), .S(_01853__PTR2), .Z(_02084__PTR175) );
  MUX2_X1 U5704 ( .A(P1_P1_InstAddrPointer_PTR16), .B(_02810__PTR16), .S(_01853__PTR2), .Z(_02084__PTR176) );
  MUX2_X1 U5705 ( .A(P1_P1_InstAddrPointer_PTR17), .B(_02810__PTR17), .S(_01853__PTR2), .Z(_02084__PTR177) );
  MUX2_X1 U5706 ( .A(P1_P1_InstAddrPointer_PTR18), .B(_02810__PTR18), .S(_01853__PTR2), .Z(_02084__PTR178) );
  MUX2_X1 U5707 ( .A(P1_P1_InstAddrPointer_PTR19), .B(_02810__PTR19), .S(_01853__PTR2), .Z(_02084__PTR179) );
  MUX2_X1 U5708 ( .A(P1_P1_InstAddrPointer_PTR20), .B(_02810__PTR20), .S(_01853__PTR2), .Z(_02084__PTR180) );
  MUX2_X1 U5709 ( .A(P1_P1_InstAddrPointer_PTR21), .B(_02810__PTR21), .S(_01853__PTR2), .Z(_02084__PTR181) );
  MUX2_X1 U5710 ( .A(P1_P1_InstAddrPointer_PTR22), .B(_02810__PTR22), .S(_01853__PTR2), .Z(_02084__PTR182) );
  MUX2_X1 U5711 ( .A(P1_P1_InstAddrPointer_PTR23), .B(_02810__PTR23), .S(_01853__PTR2), .Z(_02084__PTR183) );
  MUX2_X1 U5712 ( .A(P1_P1_InstAddrPointer_PTR24), .B(_02810__PTR24), .S(_01853__PTR2), .Z(_02084__PTR184) );
  MUX2_X1 U5713 ( .A(P1_P1_InstAddrPointer_PTR25), .B(_02810__PTR25), .S(_01853__PTR2), .Z(_02084__PTR185) );
  MUX2_X1 U5714 ( .A(P1_P1_InstAddrPointer_PTR26), .B(_02810__PTR26), .S(_01853__PTR2), .Z(_02084__PTR186) );
  MUX2_X1 U5715 ( .A(P1_P1_InstAddrPointer_PTR27), .B(_02810__PTR27), .S(_01853__PTR2), .Z(_02084__PTR187) );
  MUX2_X1 U5716 ( .A(P1_P1_InstAddrPointer_PTR28), .B(_02810__PTR28), .S(_01853__PTR2), .Z(_02084__PTR188) );
  MUX2_X1 U5717 ( .A(P1_P1_InstAddrPointer_PTR29), .B(_02810__PTR29), .S(_01853__PTR2), .Z(_02084__PTR189) );
  MUX2_X1 U5718 ( .A(P1_P1_InstAddrPointer_PTR30), .B(_02810__PTR30), .S(_01853__PTR2), .Z(_02084__PTR190) );
  MUX2_X1 U5719 ( .A(P1_P1_InstAddrPointer_PTR31), .B(_02810__PTR31), .S(_01853__PTR2), .Z(_02084__PTR191) );
  MUX2_X1 U5720 ( .A(P1_rEIP_PTR0), .B(_01884__PTR3), .S(_02006_), .Z(_02104__PTR32) );
  MUX2_X1 U5721 ( .A(P1_rEIP_PTR1), .B(_01884__PTR4), .S(_02006_), .Z(_02104__PTR33) );
  MUX2_X1 U5722 ( .A(P1_rEIP_PTR2), .B(_01884__PTR5), .S(_02006_), .Z(_02104__PTR34) );
  MUX2_X1 U5723 ( .A(P1_rEIP_PTR3), .B(_01884__PTR6), .S(_02006_), .Z(_02104__PTR35) );
  MUX2_X1 U5724 ( .A(P1_rEIP_PTR4), .B(_02800__PTR4), .S(_02006_), .Z(_02104__PTR36) );
  MUX2_X1 U5725 ( .A(P1_rEIP_PTR5), .B(_02799__PTR4), .S(_02006_), .Z(_02104__PTR37) );
  MUX2_X1 U5726 ( .A(P1_rEIP_PTR6), .B(1'b0), .S(_02006_), .Z(_02104__PTR38) );
  MUX2_X1 U5727 ( .A(P1_rEIP_PTR7), .B(1'b0), .S(_02006_), .Z(_02104__PTR39) );
  MUX2_X1 U5728 ( .A(P1_rEIP_PTR8), .B(1'b0), .S(_02006_), .Z(_02104__PTR40) );
  MUX2_X1 U5729 ( .A(P1_rEIP_PTR9), .B(1'b0), .S(_02006_), .Z(_02104__PTR41) );
  MUX2_X1 U5730 ( .A(P1_rEIP_PTR10), .B(1'b0), .S(_02006_), .Z(_02104__PTR42) );
  MUX2_X1 U5731 ( .A(P1_rEIP_PTR11), .B(1'b0), .S(_02006_), .Z(_02104__PTR43) );
  MUX2_X1 U5732 ( .A(P1_rEIP_PTR12), .B(1'b0), .S(_02006_), .Z(_02104__PTR44) );
  MUX2_X1 U5733 ( .A(P1_rEIP_PTR13), .B(1'b0), .S(_02006_), .Z(_02104__PTR45) );
  MUX2_X1 U5734 ( .A(P1_rEIP_PTR14), .B(1'b0), .S(_02006_), .Z(_02104__PTR46) );
  MUX2_X1 U5735 ( .A(P1_rEIP_PTR15), .B(1'b0), .S(_02006_), .Z(_02104__PTR47) );
  MUX2_X1 U5736 ( .A(P1_rEIP_PTR16), .B(1'b0), .S(_02006_), .Z(_02104__PTR48) );
  MUX2_X1 U5737 ( .A(P1_rEIP_PTR17), .B(1'b0), .S(_02006_), .Z(_02104__PTR49) );
  MUX2_X1 U5738 ( .A(P1_rEIP_PTR18), .B(1'b0), .S(_02006_), .Z(_02104__PTR50) );
  MUX2_X1 U5739 ( .A(P1_rEIP_PTR19), .B(1'b0), .S(_02006_), .Z(_02104__PTR51) );
  MUX2_X1 U5740 ( .A(P1_rEIP_PTR20), .B(1'b0), .S(_02006_), .Z(_02104__PTR52) );
  MUX2_X1 U5741 ( .A(P1_rEIP_PTR21), .B(1'b0), .S(_02006_), .Z(_02104__PTR53) );
  MUX2_X1 U5742 ( .A(P1_rEIP_PTR22), .B(1'b0), .S(_02006_), .Z(_02104__PTR54) );
  MUX2_X1 U5743 ( .A(P1_rEIP_PTR23), .B(1'b0), .S(_02006_), .Z(_02104__PTR55) );
  MUX2_X1 U5744 ( .A(P1_rEIP_PTR24), .B(1'b0), .S(_02006_), .Z(_02104__PTR56) );
  MUX2_X1 U5745 ( .A(P1_rEIP_PTR25), .B(1'b0), .S(_02006_), .Z(_02104__PTR57) );
  MUX2_X1 U5746 ( .A(P1_rEIP_PTR26), .B(1'b0), .S(_02006_), .Z(_02104__PTR58) );
  MUX2_X1 U5747 ( .A(P1_rEIP_PTR27), .B(1'b0), .S(_02006_), .Z(_02104__PTR59) );
  MUX2_X1 U5748 ( .A(P1_rEIP_PTR28), .B(1'b0), .S(_02006_), .Z(_02104__PTR60) );
  MUX2_X1 U5749 ( .A(P1_rEIP_PTR29), .B(1'b0), .S(_02006_), .Z(_02104__PTR61) );
  MUX2_X1 U5750 ( .A(P1_rEIP_PTR30), .B(1'b0), .S(_02006_), .Z(_02104__PTR62) );
  MUX2_X1 U5751 ( .A(P1_rEIP_PTR31), .B(1'b0), .S(_02006_), .Z(_02104__PTR63) );
  MUX2_X1 U5752 ( .A(P1_rEIP_PTR0), .B(_02033__PTR0), .S(_02006_), .Z(_02104__PTR64) );
  MUX2_X1 U5753 ( .A(P1_rEIP_PTR1), .B(_02033__PTR1), .S(_02006_), .Z(_02104__PTR65) );
  MUX2_X1 U5754 ( .A(P1_rEIP_PTR2), .B(_02033__PTR2), .S(_02006_), .Z(_02104__PTR66) );
  MUX2_X1 U5755 ( .A(P1_rEIP_PTR3), .B(_02033__PTR3), .S(_02006_), .Z(_02104__PTR67) );
  MUX2_X1 U5756 ( .A(P1_rEIP_PTR4), .B(_02033__PTR4), .S(_02006_), .Z(_02104__PTR68) );
  MUX2_X1 U5757 ( .A(P1_rEIP_PTR5), .B(_02033__PTR5), .S(_02006_), .Z(_02104__PTR69) );
  MUX2_X1 U5758 ( .A(P1_rEIP_PTR6), .B(_02033__PTR6), .S(_02006_), .Z(_02104__PTR70) );
  MUX2_X1 U5759 ( .A(P1_rEIP_PTR7), .B(_02033__PTR7), .S(_02006_), .Z(_02104__PTR71) );
  MUX2_X1 U5760 ( .A(P1_rEIP_PTR8), .B(_02033__PTR8), .S(_02006_), .Z(_02104__PTR72) );
  MUX2_X1 U5761 ( .A(P1_rEIP_PTR9), .B(_02033__PTR9), .S(_02006_), .Z(_02104__PTR73) );
  MUX2_X1 U5762 ( .A(P1_rEIP_PTR10), .B(_02033__PTR10), .S(_02006_), .Z(_02104__PTR74) );
  MUX2_X1 U5763 ( .A(P1_rEIP_PTR11), .B(_02033__PTR11), .S(_02006_), .Z(_02104__PTR75) );
  MUX2_X1 U5764 ( .A(P1_rEIP_PTR12), .B(_02033__PTR12), .S(_02006_), .Z(_02104__PTR76) );
  MUX2_X1 U5765 ( .A(P1_rEIP_PTR13), .B(_02033__PTR13), .S(_02006_), .Z(_02104__PTR77) );
  MUX2_X1 U5766 ( .A(P1_rEIP_PTR14), .B(_02033__PTR14), .S(_02006_), .Z(_02104__PTR78) );
  MUX2_X1 U5767 ( .A(P1_rEIP_PTR15), .B(_02033__PTR15), .S(_02006_), .Z(_02104__PTR79) );
  MUX2_X1 U5768 ( .A(P1_rEIP_PTR16), .B(_02033__PTR16), .S(_02006_), .Z(_02104__PTR80) );
  MUX2_X1 U5769 ( .A(P1_rEIP_PTR17), .B(_02033__PTR17), .S(_02006_), .Z(_02104__PTR81) );
  MUX2_X1 U5770 ( .A(P1_rEIP_PTR18), .B(_02033__PTR18), .S(_02006_), .Z(_02104__PTR82) );
  MUX2_X1 U5771 ( .A(P1_rEIP_PTR19), .B(_02033__PTR19), .S(_02006_), .Z(_02104__PTR83) );
  MUX2_X1 U5772 ( .A(P1_rEIP_PTR20), .B(_02033__PTR20), .S(_02006_), .Z(_02104__PTR84) );
  MUX2_X1 U5773 ( .A(P1_rEIP_PTR21), .B(_02033__PTR21), .S(_02006_), .Z(_02104__PTR85) );
  MUX2_X1 U5774 ( .A(P1_rEIP_PTR22), .B(_02033__PTR22), .S(_02006_), .Z(_02104__PTR86) );
  MUX2_X1 U5775 ( .A(P1_rEIP_PTR23), .B(_02033__PTR23), .S(_02006_), .Z(_02104__PTR87) );
  MUX2_X1 U5776 ( .A(P1_rEIP_PTR24), .B(_02033__PTR24), .S(_02006_), .Z(_02104__PTR88) );
  MUX2_X1 U5777 ( .A(P1_rEIP_PTR25), .B(_02033__PTR25), .S(_02006_), .Z(_02104__PTR89) );
  MUX2_X1 U5778 ( .A(P1_rEIP_PTR26), .B(_02033__PTR26), .S(_02006_), .Z(_02104__PTR90) );
  MUX2_X1 U5779 ( .A(P1_rEIP_PTR27), .B(_02033__PTR27), .S(_02006_), .Z(_02104__PTR91) );
  MUX2_X1 U5780 ( .A(P1_rEIP_PTR28), .B(_02033__PTR28), .S(_02006_), .Z(_02104__PTR92) );
  MUX2_X1 U5781 ( .A(P1_rEIP_PTR29), .B(_02033__PTR29), .S(_02006_), .Z(_02104__PTR93) );
  MUX2_X1 U5782 ( .A(P1_rEIP_PTR30), .B(_02033__PTR30), .S(_02006_), .Z(_02104__PTR94) );
  MUX2_X1 U5783 ( .A(P1_rEIP_PTR31), .B(_02033__PTR31), .S(_02006_), .Z(_02104__PTR95) );
  MUX2_X1 U5784 ( .A(P1_rEIP_PTR0), .B(_02015__PTR0), .S(_02006_), .Z(_02104__PTR96) );
  MUX2_X1 U5785 ( .A(P1_rEIP_PTR1), .B(_02015__PTR1), .S(_02006_), .Z(_02104__PTR97) );
  MUX2_X1 U5786 ( .A(P1_rEIP_PTR2), .B(_02015__PTR2), .S(_02006_), .Z(_02104__PTR98) );
  MUX2_X1 U5787 ( .A(P1_rEIP_PTR3), .B(_02015__PTR3), .S(_02006_), .Z(_02104__PTR99) );
  MUX2_X1 U5788 ( .A(P1_rEIP_PTR4), .B(_02015__PTR4), .S(_02006_), .Z(_02104__PTR100) );
  MUX2_X1 U5789 ( .A(P1_rEIP_PTR5), .B(_02015__PTR5), .S(_02006_), .Z(_02104__PTR101) );
  MUX2_X1 U5790 ( .A(P1_rEIP_PTR6), .B(_02015__PTR6), .S(_02006_), .Z(_02104__PTR102) );
  MUX2_X1 U5791 ( .A(P1_rEIP_PTR7), .B(_02015__PTR7), .S(_02006_), .Z(_02104__PTR103) );
  MUX2_X1 U5792 ( .A(P1_rEIP_PTR8), .B(_02015__PTR8), .S(_02006_), .Z(_02104__PTR104) );
  MUX2_X1 U5793 ( .A(P1_rEIP_PTR9), .B(_02015__PTR9), .S(_02006_), .Z(_02104__PTR105) );
  MUX2_X1 U5794 ( .A(P1_rEIP_PTR10), .B(_02015__PTR10), .S(_02006_), .Z(_02104__PTR106) );
  MUX2_X1 U5795 ( .A(P1_rEIP_PTR11), .B(_02015__PTR11), .S(_02006_), .Z(_02104__PTR107) );
  MUX2_X1 U5796 ( .A(P1_rEIP_PTR12), .B(_02015__PTR12), .S(_02006_), .Z(_02104__PTR108) );
  MUX2_X1 U5797 ( .A(P1_rEIP_PTR13), .B(_02015__PTR13), .S(_02006_), .Z(_02104__PTR109) );
  MUX2_X1 U5798 ( .A(P1_rEIP_PTR14), .B(_02015__PTR14), .S(_02006_), .Z(_02104__PTR110) );
  MUX2_X1 U5799 ( .A(P1_rEIP_PTR15), .B(_02015__PTR15), .S(_02006_), .Z(_02104__PTR111) );
  MUX2_X1 U5800 ( .A(P1_rEIP_PTR16), .B(_02015__PTR16), .S(_02006_), .Z(_02104__PTR112) );
  MUX2_X1 U5801 ( .A(P1_rEIP_PTR17), .B(_02015__PTR17), .S(_02006_), .Z(_02104__PTR113) );
  MUX2_X1 U5802 ( .A(P1_rEIP_PTR18), .B(_02015__PTR18), .S(_02006_), .Z(_02104__PTR114) );
  MUX2_X1 U5803 ( .A(P1_rEIP_PTR19), .B(_02015__PTR19), .S(_02006_), .Z(_02104__PTR115) );
  MUX2_X1 U5804 ( .A(P1_rEIP_PTR20), .B(_02015__PTR20), .S(_02006_), .Z(_02104__PTR116) );
  MUX2_X1 U5805 ( .A(P1_rEIP_PTR21), .B(_02015__PTR21), .S(_02006_), .Z(_02104__PTR117) );
  MUX2_X1 U5806 ( .A(P1_rEIP_PTR22), .B(_02015__PTR22), .S(_02006_), .Z(_02104__PTR118) );
  MUX2_X1 U5807 ( .A(P1_rEIP_PTR23), .B(_02015__PTR23), .S(_02006_), .Z(_02104__PTR119) );
  MUX2_X1 U5808 ( .A(P1_rEIP_PTR24), .B(_02015__PTR24), .S(_02006_), .Z(_02104__PTR120) );
  MUX2_X1 U5809 ( .A(P1_rEIP_PTR25), .B(_02015__PTR25), .S(_02006_), .Z(_02104__PTR121) );
  MUX2_X1 U5810 ( .A(P1_rEIP_PTR26), .B(_02015__PTR26), .S(_02006_), .Z(_02104__PTR122) );
  MUX2_X1 U5811 ( .A(P1_rEIP_PTR27), .B(_02015__PTR27), .S(_02006_), .Z(_02104__PTR123) );
  MUX2_X1 U5812 ( .A(P1_rEIP_PTR28), .B(_02015__PTR28), .S(_02006_), .Z(_02104__PTR124) );
  MUX2_X1 U5813 ( .A(P1_rEIP_PTR29), .B(_02015__PTR29), .S(_02006_), .Z(_02104__PTR125) );
  MUX2_X1 U5814 ( .A(P1_rEIP_PTR30), .B(_02015__PTR30), .S(_02006_), .Z(_02104__PTR126) );
  MUX2_X1 U5815 ( .A(P1_rEIP_PTR31), .B(_02015__PTR31), .S(_02006_), .Z(_02104__PTR127) );
  MUX2_X1 U5816 ( .A(P1_rEIP_PTR0), .B(P1_EBX_PTR0), .S(P1_StateBS16), .Z(_02010__PTR0) );
  MUX2_X1 U5817 ( .A(_01882__PTR7), .B(_02009__PTR1), .S(P1_StateBS16), .Z(_02010__PTR1) );
  MUX2_X1 U5818 ( .A(_02822__PTR1), .B(_02009__PTR2), .S(P1_StateBS16), .Z(_02010__PTR2) );
  MUX2_X1 U5819 ( .A(_02822__PTR2), .B(_02009__PTR3), .S(P1_StateBS16), .Z(_02010__PTR3) );
  MUX2_X1 U5820 ( .A(_02822__PTR3), .B(_02009__PTR4), .S(P1_StateBS16), .Z(_02010__PTR4) );
  MUX2_X1 U5821 ( .A(_02822__PTR4), .B(_02009__PTR5), .S(P1_StateBS16), .Z(_02010__PTR5) );
  MUX2_X1 U5822 ( .A(_02822__PTR5), .B(_02009__PTR6), .S(P1_StateBS16), .Z(_02010__PTR6) );
  MUX2_X1 U5823 ( .A(_02822__PTR6), .B(_02009__PTR7), .S(P1_StateBS16), .Z(_02010__PTR7) );
  MUX2_X1 U5824 ( .A(_02822__PTR7), .B(_02009__PTR8), .S(P1_StateBS16), .Z(_02010__PTR8) );
  MUX2_X1 U5825 ( .A(_02822__PTR8), .B(_02009__PTR9), .S(P1_StateBS16), .Z(_02010__PTR9) );
  MUX2_X1 U5826 ( .A(_02822__PTR9), .B(_02009__PTR10), .S(P1_StateBS16), .Z(_02010__PTR10) );
  MUX2_X1 U5827 ( .A(_02822__PTR10), .B(_02009__PTR11), .S(P1_StateBS16), .Z(_02010__PTR11) );
  MUX2_X1 U5828 ( .A(_02822__PTR11), .B(_02009__PTR12), .S(P1_StateBS16), .Z(_02010__PTR12) );
  MUX2_X1 U5829 ( .A(_02822__PTR12), .B(_02009__PTR13), .S(P1_StateBS16), .Z(_02010__PTR13) );
  MUX2_X1 U5830 ( .A(_02822__PTR13), .B(_02009__PTR14), .S(P1_StateBS16), .Z(_02010__PTR14) );
  MUX2_X1 U5831 ( .A(_02822__PTR14), .B(_02009__PTR15), .S(P1_StateBS16), .Z(_02010__PTR15) );
  MUX2_X1 U5832 ( .A(_02822__PTR15), .B(_02009__PTR16), .S(P1_StateBS16), .Z(_02010__PTR16) );
  MUX2_X1 U5833 ( .A(_02822__PTR16), .B(_02009__PTR17), .S(P1_StateBS16), .Z(_02010__PTR17) );
  MUX2_X1 U5834 ( .A(_02822__PTR17), .B(_02009__PTR18), .S(P1_StateBS16), .Z(_02010__PTR18) );
  MUX2_X1 U5835 ( .A(_02822__PTR18), .B(_02009__PTR19), .S(P1_StateBS16), .Z(_02010__PTR19) );
  MUX2_X1 U5836 ( .A(_02822__PTR19), .B(_02009__PTR20), .S(P1_StateBS16), .Z(_02010__PTR20) );
  MUX2_X1 U5837 ( .A(_02822__PTR20), .B(_02009__PTR21), .S(P1_StateBS16), .Z(_02010__PTR21) );
  MUX2_X1 U5838 ( .A(_02822__PTR21), .B(_02009__PTR22), .S(P1_StateBS16), .Z(_02010__PTR22) );
  MUX2_X1 U5839 ( .A(_02822__PTR22), .B(_02009__PTR23), .S(P1_StateBS16), .Z(_02010__PTR23) );
  MUX2_X1 U5840 ( .A(_02822__PTR23), .B(_02009__PTR24), .S(P1_StateBS16), .Z(_02010__PTR24) );
  MUX2_X1 U5841 ( .A(_02822__PTR24), .B(_02009__PTR25), .S(P1_StateBS16), .Z(_02010__PTR25) );
  MUX2_X1 U5842 ( .A(_02822__PTR25), .B(_02009__PTR26), .S(P1_StateBS16), .Z(_02010__PTR26) );
  MUX2_X1 U5843 ( .A(_02822__PTR26), .B(_02009__PTR27), .S(P1_StateBS16), .Z(_02010__PTR27) );
  MUX2_X1 U5844 ( .A(_02822__PTR27), .B(_02009__PTR28), .S(P1_StateBS16), .Z(_02010__PTR28) );
  MUX2_X1 U5845 ( .A(_02822__PTR28), .B(_02009__PTR29), .S(P1_StateBS16), .Z(_02010__PTR29) );
  MUX2_X1 U5846 ( .A(_02822__PTR29), .B(_02009__PTR30), .S(P1_StateBS16), .Z(_02010__PTR30) );
  MUX2_X1 U5847 ( .A(_02822__PTR30), .B(_02009__PTR31), .S(P1_StateBS16), .Z(_02010__PTR31) );
  MUX2_X1 U5848 ( .A(_02948__PTR1), .B(P1_EBX_PTR1), .S(_02733__PTR31), .Z(_02009__PTR1) );
  MUX2_X1 U5849 ( .A(_02948__PTR2), .B(P1_EBX_PTR2), .S(_02733__PTR31), .Z(_02009__PTR2) );
  MUX2_X1 U5850 ( .A(_02948__PTR3), .B(P1_EBX_PTR3), .S(_02733__PTR31), .Z(_02009__PTR3) );
  MUX2_X1 U5851 ( .A(_02948__PTR4), .B(P1_EBX_PTR4), .S(_02733__PTR31), .Z(_02009__PTR4) );
  MUX2_X1 U5852 ( .A(_02948__PTR5), .B(P1_EBX_PTR5), .S(_02733__PTR31), .Z(_02009__PTR5) );
  MUX2_X1 U5853 ( .A(_02948__PTR6), .B(P1_EBX_PTR6), .S(_02733__PTR31), .Z(_02009__PTR6) );
  MUX2_X1 U5854 ( .A(_02948__PTR7), .B(P1_EBX_PTR7), .S(_02733__PTR31), .Z(_02009__PTR7) );
  MUX2_X1 U5855 ( .A(_02948__PTR8), .B(P1_EBX_PTR8), .S(_02733__PTR31), .Z(_02009__PTR8) );
  MUX2_X1 U5856 ( .A(_02948__PTR9), .B(P1_EBX_PTR9), .S(_02733__PTR31), .Z(_02009__PTR9) );
  MUX2_X1 U5857 ( .A(_02948__PTR10), .B(P1_EBX_PTR10), .S(_02733__PTR31), .Z(_02009__PTR10) );
  MUX2_X1 U5858 ( .A(_02948__PTR11), .B(P1_EBX_PTR11), .S(_02733__PTR31), .Z(_02009__PTR11) );
  MUX2_X1 U5859 ( .A(_02948__PTR12), .B(P1_EBX_PTR12), .S(_02733__PTR31), .Z(_02009__PTR12) );
  MUX2_X1 U5860 ( .A(_02948__PTR13), .B(P1_EBX_PTR13), .S(_02733__PTR31), .Z(_02009__PTR13) );
  MUX2_X1 U5861 ( .A(_02948__PTR14), .B(P1_EBX_PTR14), .S(_02733__PTR31), .Z(_02009__PTR14) );
  MUX2_X1 U5862 ( .A(_02948__PTR15), .B(P1_EBX_PTR15), .S(_02733__PTR31), .Z(_02009__PTR15) );
  MUX2_X1 U5863 ( .A(_02948__PTR16), .B(P1_EBX_PTR16), .S(_02733__PTR31), .Z(_02009__PTR16) );
  MUX2_X1 U5864 ( .A(_02948__PTR17), .B(P1_EBX_PTR17), .S(_02733__PTR31), .Z(_02009__PTR17) );
  MUX2_X1 U5865 ( .A(_02948__PTR18), .B(P1_EBX_PTR18), .S(_02733__PTR31), .Z(_02009__PTR18) );
  MUX2_X1 U5866 ( .A(_02948__PTR19), .B(P1_EBX_PTR19), .S(_02733__PTR31), .Z(_02009__PTR19) );
  MUX2_X1 U5867 ( .A(_02948__PTR20), .B(P1_EBX_PTR20), .S(_02733__PTR31), .Z(_02009__PTR20) );
  MUX2_X1 U5868 ( .A(_02948__PTR21), .B(P1_EBX_PTR21), .S(_02733__PTR31), .Z(_02009__PTR21) );
  MUX2_X1 U5869 ( .A(_02948__PTR22), .B(P1_EBX_PTR22), .S(_02733__PTR31), .Z(_02009__PTR22) );
  MUX2_X1 U5870 ( .A(_02948__PTR23), .B(P1_EBX_PTR23), .S(_02733__PTR31), .Z(_02009__PTR23) );
  MUX2_X1 U5871 ( .A(_02948__PTR24), .B(P1_EBX_PTR24), .S(_02733__PTR31), .Z(_02009__PTR24) );
  MUX2_X1 U5872 ( .A(_02948__PTR25), .B(P1_EBX_PTR25), .S(_02733__PTR31), .Z(_02009__PTR25) );
  MUX2_X1 U5873 ( .A(_02948__PTR26), .B(P1_EBX_PTR26), .S(_02733__PTR31), .Z(_02009__PTR26) );
  MUX2_X1 U5874 ( .A(_02948__PTR27), .B(P1_EBX_PTR27), .S(_02733__PTR31), .Z(_02009__PTR27) );
  MUX2_X1 U5875 ( .A(_02948__PTR28), .B(P1_EBX_PTR28), .S(_02733__PTR31), .Z(_02009__PTR28) );
  MUX2_X1 U5876 ( .A(_02948__PTR29), .B(P1_EBX_PTR29), .S(_02733__PTR31), .Z(_02009__PTR29) );
  MUX2_X1 U5877 ( .A(_02948__PTR30), .B(P1_EBX_PTR30), .S(_02733__PTR31), .Z(_02009__PTR30) );
  MUX2_X1 U5878 ( .A(_02948__PTR31), .B(P1_EBX_PTR31), .S(_02733__PTR31), .Z(_02009__PTR31) );
  MUX2_X1 U5879 ( .A(P1_EBX_PTR0), .B(P1_P1_InstQueue_PTR0_PTR0), .S(_01853__PTR2), .Z(_02100__PTR64) );
  MUX2_X1 U5880 ( .A(P1_EBX_PTR1), .B(P1_P1_InstQueue_PTR0_PTR1), .S(_01853__PTR2), .Z(_02100__PTR65) );
  MUX2_X1 U5881 ( .A(P1_EBX_PTR2), .B(P1_P1_InstQueue_PTR0_PTR2), .S(_01853__PTR2), .Z(_02100__PTR66) );
  MUX2_X1 U5882 ( .A(P1_EBX_PTR3), .B(P1_P1_InstQueue_PTR0_PTR3), .S(_01853__PTR2), .Z(_02100__PTR67) );
  MUX2_X1 U5883 ( .A(P1_EBX_PTR4), .B(P1_P1_InstQueue_PTR0_PTR4), .S(_01853__PTR2), .Z(_02100__PTR68) );
  MUX2_X1 U5884 ( .A(P1_EBX_PTR5), .B(P1_P1_InstQueue_PTR0_PTR5), .S(_01853__PTR2), .Z(_02100__PTR69) );
  MUX2_X1 U5885 ( .A(P1_EBX_PTR6), .B(P1_P1_InstQueue_PTR0_PTR6), .S(_01853__PTR2), .Z(_02100__PTR70) );
  MUX2_X1 U5886 ( .A(P1_EBX_PTR7), .B(P1_P1_InstQueue_PTR0_PTR7), .S(_01853__PTR2), .Z(_02100__PTR71) );
  MUX2_X1 U5887 ( .A(P1_EBX_PTR8), .B(_01891__PTR0), .S(_01853__PTR2), .Z(_02100__PTR72) );
  MUX2_X1 U5888 ( .A(P1_EBX_PTR9), .B(_01891__PTR1), .S(_01853__PTR2), .Z(_02100__PTR73) );
  MUX2_X1 U5889 ( .A(P1_EBX_PTR10), .B(_01891__PTR2), .S(_01853__PTR2), .Z(_02100__PTR74) );
  MUX2_X1 U5890 ( .A(P1_EBX_PTR11), .B(_01891__PTR3), .S(_01853__PTR2), .Z(_02100__PTR75) );
  MUX2_X1 U5891 ( .A(P1_EBX_PTR12), .B(_01891__PTR4), .S(_01853__PTR2), .Z(_02100__PTR76) );
  MUX2_X1 U5892 ( .A(P1_EBX_PTR13), .B(_01891__PTR5), .S(_01853__PTR2), .Z(_02100__PTR77) );
  MUX2_X1 U5893 ( .A(P1_EBX_PTR14), .B(_01891__PTR6), .S(_01853__PTR2), .Z(_02100__PTR78) );
  MUX2_X1 U5894 ( .A(P1_EBX_PTR15), .B(_01891__PTR7), .S(_01853__PTR2), .Z(_02100__PTR79) );
  MUX2_X1 U5895 ( .A(P1_EBX_PTR16), .B(_01889__PTR0), .S(_01853__PTR2), .Z(_02100__PTR80) );
  MUX2_X1 U5896 ( .A(P1_EBX_PTR17), .B(_01889__PTR1), .S(_01853__PTR2), .Z(_02100__PTR81) );
  MUX2_X1 U5897 ( .A(P1_EBX_PTR18), .B(_01889__PTR2), .S(_01853__PTR2), .Z(_02100__PTR82) );
  MUX2_X1 U5898 ( .A(P1_EBX_PTR19), .B(_01889__PTR3), .S(_01853__PTR2), .Z(_02100__PTR83) );
  MUX2_X1 U5899 ( .A(P1_EBX_PTR20), .B(_01889__PTR4), .S(_01853__PTR2), .Z(_02100__PTR84) );
  MUX2_X1 U5900 ( .A(P1_EBX_PTR21), .B(_01889__PTR5), .S(_01853__PTR2), .Z(_02100__PTR85) );
  MUX2_X1 U5901 ( .A(P1_EBX_PTR22), .B(_01889__PTR6), .S(_01853__PTR2), .Z(_02100__PTR86) );
  MUX2_X1 U5902 ( .A(P1_EBX_PTR23), .B(_02815__PTR0), .S(_01853__PTR2), .Z(_02100__PTR87) );
  MUX2_X1 U5903 ( .A(P1_EBX_PTR24), .B(_02816__PTR1), .S(_01853__PTR2), .Z(_02100__PTR88) );
  MUX2_X1 U5904 ( .A(P1_EBX_PTR25), .B(_02816__PTR2), .S(_01853__PTR2), .Z(_02100__PTR89) );
  MUX2_X1 U5905 ( .A(P1_EBX_PTR26), .B(_02816__PTR3), .S(_01853__PTR2), .Z(_02100__PTR90) );
  MUX2_X1 U5906 ( .A(P1_EBX_PTR27), .B(_02816__PTR4), .S(_01853__PTR2), .Z(_02100__PTR91) );
  MUX2_X1 U5907 ( .A(P1_EBX_PTR28), .B(_02816__PTR5), .S(_01853__PTR2), .Z(_02100__PTR92) );
  MUX2_X1 U5908 ( .A(P1_EBX_PTR29), .B(_02816__PTR6), .S(_01853__PTR2), .Z(_02100__PTR93) );
  MUX2_X1 U5909 ( .A(P1_EBX_PTR30), .B(_02816__PTR7), .S(_01853__PTR2), .Z(_02100__PTR94) );
  MUX2_X1 U5910 ( .A(P1_EBX_PTR31), .B(_02814__PTR7), .S(_01853__PTR2), .Z(_02100__PTR95) );
  MUX2_X1 U5911 ( .A(P1_P1_InstQueueRd_Addr_PTR0), .B(_01884__PTR3), .S(_01853__PTR2), .Z(_02088__PTR25) );
  MUX2_X1 U5912 ( .A(P1_P1_InstQueueRd_Addr_PTR1), .B(_01884__PTR4), .S(_01853__PTR2), .Z(_02088__PTR26) );
  MUX2_X1 U5913 ( .A(P1_P1_InstQueueRd_Addr_PTR2), .B(_02820__PTR2), .S(_01853__PTR2), .Z(_02088__PTR27) );
  MUX2_X1 U5914 ( .A(P1_P1_InstQueueRd_Addr_PTR3), .B(_02820__PTR3), .S(_01853__PTR2), .Z(_02088__PTR28) );
  MUX2_X1 U5915 ( .A(P1_P1_InstQueueRd_Addr_PTR4), .B(1'b0), .S(_01853__PTR2), .Z(_02088__PTR29) );
  MUX2_X1 U5916 ( .A(P1_EAX_PTR0), .B(_01885__PTR0), .S(_01853__PTR2), .Z(_02096__PTR128) );
  MUX2_X1 U5917 ( .A(P1_EAX_PTR1), .B(_01885__PTR1), .S(_01853__PTR2), .Z(_02096__PTR129) );
  MUX2_X1 U5918 ( .A(P1_EAX_PTR2), .B(_01885__PTR2), .S(_01853__PTR2), .Z(_02096__PTR130) );
  MUX2_X1 U5919 ( .A(P1_EAX_PTR3), .B(_01885__PTR3), .S(_01853__PTR2), .Z(_02096__PTR131) );
  MUX2_X1 U5920 ( .A(P1_EAX_PTR4), .B(_01885__PTR4), .S(_01853__PTR2), .Z(_02096__PTR132) );
  MUX2_X1 U5921 ( .A(P1_EAX_PTR5), .B(_01885__PTR5), .S(_01853__PTR2), .Z(_02096__PTR133) );
  MUX2_X1 U5922 ( .A(P1_EAX_PTR6), .B(_01885__PTR6), .S(_01853__PTR2), .Z(_02096__PTR134) );
  MUX2_X1 U5923 ( .A(P1_EAX_PTR7), .B(_01885__PTR7), .S(_01853__PTR2), .Z(_02096__PTR135) );
  MUX2_X1 U5924 ( .A(P1_EAX_PTR8), .B(_01891__PTR0), .S(_01853__PTR2), .Z(_02096__PTR136) );
  MUX2_X1 U5925 ( .A(P1_EAX_PTR9), .B(_01891__PTR1), .S(_01853__PTR2), .Z(_02096__PTR137) );
  MUX2_X1 U5926 ( .A(P1_EAX_PTR10), .B(_01891__PTR2), .S(_01853__PTR2), .Z(_02096__PTR138) );
  MUX2_X1 U5927 ( .A(P1_EAX_PTR11), .B(_01891__PTR3), .S(_01853__PTR2), .Z(_02096__PTR139) );
  MUX2_X1 U5928 ( .A(P1_EAX_PTR12), .B(_01891__PTR4), .S(_01853__PTR2), .Z(_02096__PTR140) );
  MUX2_X1 U5929 ( .A(P1_EAX_PTR13), .B(_01891__PTR5), .S(_01853__PTR2), .Z(_02096__PTR141) );
  MUX2_X1 U5930 ( .A(P1_EAX_PTR14), .B(_01891__PTR6), .S(_01853__PTR2), .Z(_02096__PTR142) );
  MUX2_X1 U5931 ( .A(P1_EAX_PTR15), .B(_01891__PTR7), .S(_01853__PTR2), .Z(_02096__PTR143) );
  MUX2_X1 U5932 ( .A(P1_EAX_PTR16), .B(_01889__PTR0), .S(_01853__PTR2), .Z(_02096__PTR144) );
  MUX2_X1 U5933 ( .A(P1_EAX_PTR17), .B(_01889__PTR1), .S(_01853__PTR2), .Z(_02096__PTR145) );
  MUX2_X1 U5934 ( .A(P1_EAX_PTR18), .B(_01889__PTR2), .S(_01853__PTR2), .Z(_02096__PTR146) );
  MUX2_X1 U5935 ( .A(P1_EAX_PTR19), .B(_01889__PTR3), .S(_01853__PTR2), .Z(_02096__PTR147) );
  MUX2_X1 U5936 ( .A(P1_EAX_PTR20), .B(_01889__PTR4), .S(_01853__PTR2), .Z(_02096__PTR148) );
  MUX2_X1 U5937 ( .A(P1_EAX_PTR21), .B(_01889__PTR5), .S(_01853__PTR2), .Z(_02096__PTR149) );
  MUX2_X1 U5938 ( .A(P1_EAX_PTR22), .B(_01889__PTR6), .S(_01853__PTR2), .Z(_02096__PTR150) );
  MUX2_X1 U5939 ( .A(P1_EAX_PTR23), .B(_02815__PTR0), .S(_01853__PTR2), .Z(_02096__PTR151) );
  MUX2_X1 U5940 ( .A(P1_EAX_PTR24), .B(_02816__PTR1), .S(_01853__PTR2), .Z(_02096__PTR152) );
  MUX2_X1 U5941 ( .A(P1_EAX_PTR25), .B(_02816__PTR2), .S(_01853__PTR2), .Z(_02096__PTR153) );
  MUX2_X1 U5942 ( .A(P1_EAX_PTR26), .B(_02816__PTR3), .S(_01853__PTR2), .Z(_02096__PTR154) );
  MUX2_X1 U5943 ( .A(P1_EAX_PTR27), .B(_02816__PTR4), .S(_01853__PTR2), .Z(_02096__PTR155) );
  MUX2_X1 U5944 ( .A(P1_EAX_PTR28), .B(_02816__PTR5), .S(_01853__PTR2), .Z(_02096__PTR156) );
  MUX2_X1 U5945 ( .A(P1_EAX_PTR29), .B(_02816__PTR6), .S(_01853__PTR2), .Z(_02096__PTR157) );
  MUX2_X1 U5946 ( .A(P1_EAX_PTR30), .B(_02816__PTR7), .S(_01853__PTR2), .Z(_02096__PTR158) );
  MUX2_X1 U5947 ( .A(P1_EAX_PTR31), .B(_02814__PTR7), .S(_01853__PTR2), .Z(_02096__PTR159) );
  MUX2_X1 U5948 ( .A(P1_P1_PhyAddrPointer_PTR0), .B(_02809__PTR0), .S(_01853__PTR2), .Z(_02092__PTR32) );
  MUX2_X1 U5949 ( .A(P1_P1_PhyAddrPointer_PTR1), .B(_02810__PTR1), .S(_01853__PTR2), .Z(_02092__PTR33) );
  MUX2_X1 U5950 ( .A(P1_P1_PhyAddrPointer_PTR2), .B(_02810__PTR2), .S(_01853__PTR2), .Z(_02092__PTR34) );
  MUX2_X1 U5951 ( .A(P1_P1_PhyAddrPointer_PTR3), .B(_02810__PTR3), .S(_01853__PTR2), .Z(_02092__PTR35) );
  MUX2_X1 U5952 ( .A(P1_P1_PhyAddrPointer_PTR4), .B(_02810__PTR4), .S(_01853__PTR2), .Z(_02092__PTR36) );
  MUX2_X1 U5953 ( .A(P1_P1_PhyAddrPointer_PTR5), .B(_02810__PTR5), .S(_01853__PTR2), .Z(_02092__PTR37) );
  MUX2_X1 U5954 ( .A(P1_P1_PhyAddrPointer_PTR6), .B(_02810__PTR6), .S(_01853__PTR2), .Z(_02092__PTR38) );
  MUX2_X1 U5955 ( .A(P1_P1_PhyAddrPointer_PTR7), .B(_02810__PTR7), .S(_01853__PTR2), .Z(_02092__PTR39) );
  MUX2_X1 U5956 ( .A(P1_P1_PhyAddrPointer_PTR8), .B(_02810__PTR8), .S(_01853__PTR2), .Z(_02092__PTR40) );
  MUX2_X1 U5957 ( .A(P1_P1_PhyAddrPointer_PTR9), .B(_02810__PTR9), .S(_01853__PTR2), .Z(_02092__PTR41) );
  MUX2_X1 U5958 ( .A(P1_P1_PhyAddrPointer_PTR10), .B(_02810__PTR10), .S(_01853__PTR2), .Z(_02092__PTR42) );
  MUX2_X1 U5959 ( .A(P1_P1_PhyAddrPointer_PTR11), .B(_02810__PTR11), .S(_01853__PTR2), .Z(_02092__PTR43) );
  MUX2_X1 U5960 ( .A(P1_P1_PhyAddrPointer_PTR12), .B(_02810__PTR12), .S(_01853__PTR2), .Z(_02092__PTR44) );
  MUX2_X1 U5961 ( .A(P1_P1_PhyAddrPointer_PTR13), .B(_02810__PTR13), .S(_01853__PTR2), .Z(_02092__PTR45) );
  MUX2_X1 U5962 ( .A(P1_P1_PhyAddrPointer_PTR14), .B(_02810__PTR14), .S(_01853__PTR2), .Z(_02092__PTR46) );
  MUX2_X1 U5963 ( .A(P1_P1_PhyAddrPointer_PTR15), .B(_02810__PTR15), .S(_01853__PTR2), .Z(_02092__PTR47) );
  MUX2_X1 U5964 ( .A(P1_P1_PhyAddrPointer_PTR16), .B(_02810__PTR16), .S(_01853__PTR2), .Z(_02092__PTR48) );
  MUX2_X1 U5965 ( .A(P1_P1_PhyAddrPointer_PTR17), .B(_02810__PTR17), .S(_01853__PTR2), .Z(_02092__PTR49) );
  MUX2_X1 U5966 ( .A(P1_P1_PhyAddrPointer_PTR18), .B(_02810__PTR18), .S(_01853__PTR2), .Z(_02092__PTR50) );
  MUX2_X1 U5967 ( .A(P1_P1_PhyAddrPointer_PTR19), .B(_02810__PTR19), .S(_01853__PTR2), .Z(_02092__PTR51) );
  MUX2_X1 U5968 ( .A(P1_P1_PhyAddrPointer_PTR20), .B(_02810__PTR20), .S(_01853__PTR2), .Z(_02092__PTR52) );
  MUX2_X1 U5969 ( .A(P1_P1_PhyAddrPointer_PTR21), .B(_02810__PTR21), .S(_01853__PTR2), .Z(_02092__PTR53) );
  MUX2_X1 U5970 ( .A(P1_P1_PhyAddrPointer_PTR22), .B(_02810__PTR22), .S(_01853__PTR2), .Z(_02092__PTR54) );
  MUX2_X1 U5971 ( .A(P1_P1_PhyAddrPointer_PTR23), .B(_02810__PTR23), .S(_01853__PTR2), .Z(_02092__PTR55) );
  MUX2_X1 U5972 ( .A(P1_P1_PhyAddrPointer_PTR24), .B(_02810__PTR24), .S(_01853__PTR2), .Z(_02092__PTR56) );
  MUX2_X1 U5973 ( .A(P1_P1_PhyAddrPointer_PTR25), .B(_02810__PTR25), .S(_01853__PTR2), .Z(_02092__PTR57) );
  MUX2_X1 U5974 ( .A(P1_P1_PhyAddrPointer_PTR26), .B(_02810__PTR26), .S(_01853__PTR2), .Z(_02092__PTR58) );
  MUX2_X1 U5975 ( .A(P1_P1_PhyAddrPointer_PTR27), .B(_02810__PTR27), .S(_01853__PTR2), .Z(_02092__PTR59) );
  MUX2_X1 U5976 ( .A(P1_P1_PhyAddrPointer_PTR28), .B(_02810__PTR28), .S(_01853__PTR2), .Z(_02092__PTR60) );
  MUX2_X1 U5977 ( .A(P1_P1_PhyAddrPointer_PTR29), .B(_02810__PTR29), .S(_01853__PTR2), .Z(_02092__PTR61) );
  MUX2_X1 U5978 ( .A(P1_P1_PhyAddrPointer_PTR30), .B(_02810__PTR30), .S(_01853__PTR2), .Z(_02092__PTR62) );
  MUX2_X1 U5979 ( .A(P1_P1_PhyAddrPointer_PTR31), .B(_02810__PTR31), .S(_01853__PTR2), .Z(_02092__PTR63) );
  MUX2_X1 U5980 ( .A(P1_P1_InstAddrPointer_PTR1), .B(_02037__PTR1), .S(_02006_), .Z(_02084__PTR65) );
  MUX2_X1 U5981 ( .A(P1_P1_InstAddrPointer_PTR2), .B(_02037__PTR2), .S(_02006_), .Z(_02084__PTR66) );
  MUX2_X1 U5982 ( .A(P1_P1_InstAddrPointer_PTR3), .B(_02037__PTR3), .S(_02006_), .Z(_02084__PTR67) );
  MUX2_X1 U5983 ( .A(P1_P1_InstAddrPointer_PTR4), .B(_02037__PTR4), .S(_02006_), .Z(_02084__PTR68) );
  MUX2_X1 U5984 ( .A(P1_P1_InstAddrPointer_PTR5), .B(_02037__PTR5), .S(_02006_), .Z(_02084__PTR69) );
  MUX2_X1 U5985 ( .A(P1_P1_InstAddrPointer_PTR6), .B(_02037__PTR6), .S(_02006_), .Z(_02084__PTR70) );
  MUX2_X1 U5986 ( .A(P1_P1_InstAddrPointer_PTR7), .B(_02037__PTR7), .S(_02006_), .Z(_02084__PTR71) );
  MUX2_X1 U5987 ( .A(P1_P1_InstAddrPointer_PTR8), .B(_02037__PTR8), .S(_02006_), .Z(_02084__PTR72) );
  MUX2_X1 U5988 ( .A(P1_P1_InstAddrPointer_PTR9), .B(_02037__PTR9), .S(_02006_), .Z(_02084__PTR73) );
  MUX2_X1 U5989 ( .A(P1_P1_InstAddrPointer_PTR10), .B(_02037__PTR10), .S(_02006_), .Z(_02084__PTR74) );
  MUX2_X1 U5990 ( .A(P1_P1_InstAddrPointer_PTR11), .B(_02037__PTR11), .S(_02006_), .Z(_02084__PTR75) );
  MUX2_X1 U5991 ( .A(P1_P1_InstAddrPointer_PTR12), .B(_02037__PTR12), .S(_02006_), .Z(_02084__PTR76) );
  MUX2_X1 U5992 ( .A(P1_P1_InstAddrPointer_PTR13), .B(_02037__PTR13), .S(_02006_), .Z(_02084__PTR77) );
  MUX2_X1 U5993 ( .A(P1_P1_InstAddrPointer_PTR14), .B(_02037__PTR14), .S(_02006_), .Z(_02084__PTR78) );
  MUX2_X1 U5994 ( .A(P1_P1_InstAddrPointer_PTR15), .B(_02037__PTR15), .S(_02006_), .Z(_02084__PTR79) );
  MUX2_X1 U5995 ( .A(P1_P1_InstAddrPointer_PTR16), .B(_02037__PTR16), .S(_02006_), .Z(_02084__PTR80) );
  MUX2_X1 U5996 ( .A(P1_P1_InstAddrPointer_PTR17), .B(_02037__PTR17), .S(_02006_), .Z(_02084__PTR81) );
  MUX2_X1 U5997 ( .A(P1_P1_InstAddrPointer_PTR18), .B(_02037__PTR18), .S(_02006_), .Z(_02084__PTR82) );
  MUX2_X1 U5998 ( .A(P1_P1_InstAddrPointer_PTR19), .B(_02037__PTR19), .S(_02006_), .Z(_02084__PTR83) );
  MUX2_X1 U5999 ( .A(P1_P1_InstAddrPointer_PTR20), .B(_02037__PTR20), .S(_02006_), .Z(_02084__PTR84) );
  MUX2_X1 U6000 ( .A(P1_P1_InstAddrPointer_PTR21), .B(_02037__PTR21), .S(_02006_), .Z(_02084__PTR85) );
  MUX2_X1 U6001 ( .A(P1_P1_InstAddrPointer_PTR22), .B(_02037__PTR22), .S(_02006_), .Z(_02084__PTR86) );
  MUX2_X1 U6002 ( .A(P1_P1_InstAddrPointer_PTR23), .B(_02037__PTR23), .S(_02006_), .Z(_02084__PTR87) );
  MUX2_X1 U6003 ( .A(P1_P1_InstAddrPointer_PTR24), .B(_02037__PTR24), .S(_02006_), .Z(_02084__PTR88) );
  MUX2_X1 U6004 ( .A(P1_P1_InstAddrPointer_PTR25), .B(_02037__PTR25), .S(_02006_), .Z(_02084__PTR89) );
  MUX2_X1 U6005 ( .A(P1_P1_InstAddrPointer_PTR26), .B(_02037__PTR26), .S(_02006_), .Z(_02084__PTR90) );
  MUX2_X1 U6006 ( .A(P1_P1_InstAddrPointer_PTR27), .B(_02037__PTR27), .S(_02006_), .Z(_02084__PTR91) );
  MUX2_X1 U6007 ( .A(P1_P1_InstAddrPointer_PTR28), .B(_02037__PTR28), .S(_02006_), .Z(_02084__PTR92) );
  MUX2_X1 U6008 ( .A(P1_P1_InstAddrPointer_PTR29), .B(_02037__PTR29), .S(_02006_), .Z(_02084__PTR93) );
  MUX2_X1 U6009 ( .A(P1_P1_InstAddrPointer_PTR30), .B(_02037__PTR30), .S(_02006_), .Z(_02084__PTR94) );
  MUX2_X1 U6010 ( .A(P1_P1_InstAddrPointer_PTR31), .B(_02037__PTR31), .S(_02006_), .Z(_02084__PTR95) );
  MUX2_X1 U6011 ( .A(P1_P1_InstAddrPointer_PTR1), .B(_02019__PTR1), .S(_02006_), .Z(_02084__PTR97) );
  MUX2_X1 U6012 ( .A(P1_P1_InstAddrPointer_PTR2), .B(_02019__PTR2), .S(_02006_), .Z(_02084__PTR98) );
  MUX2_X1 U6013 ( .A(P1_P1_InstAddrPointer_PTR3), .B(_02019__PTR3), .S(_02006_), .Z(_02084__PTR99) );
  MUX2_X1 U6014 ( .A(P1_P1_InstAddrPointer_PTR4), .B(_02019__PTR4), .S(_02006_), .Z(_02084__PTR100) );
  MUX2_X1 U6015 ( .A(P1_P1_InstAddrPointer_PTR5), .B(_02019__PTR5), .S(_02006_), .Z(_02084__PTR101) );
  MUX2_X1 U6016 ( .A(P1_P1_InstAddrPointer_PTR6), .B(_02019__PTR6), .S(_02006_), .Z(_02084__PTR102) );
  MUX2_X1 U6017 ( .A(P1_P1_InstAddrPointer_PTR7), .B(_02019__PTR7), .S(_02006_), .Z(_02084__PTR103) );
  MUX2_X1 U6018 ( .A(P1_P1_InstAddrPointer_PTR8), .B(_02019__PTR8), .S(_02006_), .Z(_02084__PTR104) );
  MUX2_X1 U6019 ( .A(P1_P1_InstAddrPointer_PTR9), .B(_02019__PTR9), .S(_02006_), .Z(_02084__PTR105) );
  MUX2_X1 U6020 ( .A(P1_P1_InstAddrPointer_PTR10), .B(_02019__PTR10), .S(_02006_), .Z(_02084__PTR106) );
  MUX2_X1 U6021 ( .A(P1_P1_InstAddrPointer_PTR11), .B(_02019__PTR11), .S(_02006_), .Z(_02084__PTR107) );
  MUX2_X1 U6022 ( .A(P1_P1_InstAddrPointer_PTR12), .B(_02019__PTR12), .S(_02006_), .Z(_02084__PTR108) );
  MUX2_X1 U6023 ( .A(P1_P1_InstAddrPointer_PTR13), .B(_02019__PTR13), .S(_02006_), .Z(_02084__PTR109) );
  MUX2_X1 U6024 ( .A(P1_P1_InstAddrPointer_PTR14), .B(_02019__PTR14), .S(_02006_), .Z(_02084__PTR110) );
  MUX2_X1 U6025 ( .A(P1_P1_InstAddrPointer_PTR15), .B(_02019__PTR15), .S(_02006_), .Z(_02084__PTR111) );
  MUX2_X1 U6026 ( .A(P1_P1_InstAddrPointer_PTR16), .B(_02019__PTR16), .S(_02006_), .Z(_02084__PTR112) );
  MUX2_X1 U6027 ( .A(P1_P1_InstAddrPointer_PTR17), .B(_02019__PTR17), .S(_02006_), .Z(_02084__PTR113) );
  MUX2_X1 U6028 ( .A(P1_P1_InstAddrPointer_PTR18), .B(_02019__PTR18), .S(_02006_), .Z(_02084__PTR114) );
  MUX2_X1 U6029 ( .A(P1_P1_InstAddrPointer_PTR19), .B(_02019__PTR19), .S(_02006_), .Z(_02084__PTR115) );
  MUX2_X1 U6030 ( .A(P1_P1_InstAddrPointer_PTR20), .B(_02019__PTR20), .S(_02006_), .Z(_02084__PTR116) );
  MUX2_X1 U6031 ( .A(P1_P1_InstAddrPointer_PTR21), .B(_02019__PTR21), .S(_02006_), .Z(_02084__PTR117) );
  MUX2_X1 U6032 ( .A(P1_P1_InstAddrPointer_PTR22), .B(_02019__PTR22), .S(_02006_), .Z(_02084__PTR118) );
  MUX2_X1 U6033 ( .A(P1_P1_InstAddrPointer_PTR23), .B(_02019__PTR23), .S(_02006_), .Z(_02084__PTR119) );
  MUX2_X1 U6034 ( .A(P1_P1_InstAddrPointer_PTR24), .B(_02019__PTR24), .S(_02006_), .Z(_02084__PTR120) );
  MUX2_X1 U6035 ( .A(P1_P1_InstAddrPointer_PTR25), .B(_02019__PTR25), .S(_02006_), .Z(_02084__PTR121) );
  MUX2_X1 U6036 ( .A(P1_P1_InstAddrPointer_PTR26), .B(_02019__PTR26), .S(_02006_), .Z(_02084__PTR122) );
  MUX2_X1 U6037 ( .A(P1_P1_InstAddrPointer_PTR27), .B(_02019__PTR27), .S(_02006_), .Z(_02084__PTR123) );
  MUX2_X1 U6038 ( .A(P1_P1_InstAddrPointer_PTR28), .B(_02019__PTR28), .S(_02006_), .Z(_02084__PTR124) );
  MUX2_X1 U6039 ( .A(P1_P1_InstAddrPointer_PTR29), .B(_02019__PTR29), .S(_02006_), .Z(_02084__PTR125) );
  MUX2_X1 U6040 ( .A(P1_P1_InstAddrPointer_PTR30), .B(_02019__PTR30), .S(_02006_), .Z(_02084__PTR126) );
  MUX2_X1 U6041 ( .A(P1_P1_InstAddrPointer_PTR31), .B(_02019__PTR31), .S(_02006_), .Z(_02084__PTR127) );
  MUX2_X1 U6042 ( .A(P1_P1_InstAddrPointer_PTR0), .B(_01998__PTR0), .S(_01853__PTR3), .Z(_02084__PTR192) );
  MUX2_X1 U6043 ( .A(P1_P1_InstAddrPointer_PTR1), .B(_01998__PTR1), .S(_01853__PTR3), .Z(_02084__PTR193) );
  MUX2_X1 U6044 ( .A(P1_P1_InstAddrPointer_PTR2), .B(_01998__PTR2), .S(_01853__PTR3), .Z(_02084__PTR194) );
  MUX2_X1 U6045 ( .A(P1_P1_InstAddrPointer_PTR3), .B(_01998__PTR3), .S(_01853__PTR3), .Z(_02084__PTR195) );
  MUX2_X1 U6046 ( .A(P1_P1_InstAddrPointer_PTR4), .B(_01998__PTR4), .S(_01853__PTR3), .Z(_02084__PTR196) );
  MUX2_X1 U6047 ( .A(P1_P1_InstAddrPointer_PTR5), .B(_01998__PTR5), .S(_01853__PTR3), .Z(_02084__PTR197) );
  MUX2_X1 U6048 ( .A(P1_P1_InstAddrPointer_PTR6), .B(_01998__PTR6), .S(_01853__PTR3), .Z(_02084__PTR198) );
  MUX2_X1 U6049 ( .A(P1_P1_InstAddrPointer_PTR7), .B(_01998__PTR7), .S(_01853__PTR3), .Z(_02084__PTR199) );
  MUX2_X1 U6050 ( .A(P1_P1_InstAddrPointer_PTR8), .B(_01998__PTR8), .S(_01853__PTR3), .Z(_02084__PTR200) );
  MUX2_X1 U6051 ( .A(P1_P1_InstAddrPointer_PTR9), .B(_01998__PTR9), .S(_01853__PTR3), .Z(_02084__PTR201) );
  MUX2_X1 U6052 ( .A(P1_P1_InstAddrPointer_PTR10), .B(_01998__PTR10), .S(_01853__PTR3), .Z(_02084__PTR202) );
  MUX2_X1 U6053 ( .A(P1_P1_InstAddrPointer_PTR11), .B(_01998__PTR11), .S(_01853__PTR3), .Z(_02084__PTR203) );
  MUX2_X1 U6054 ( .A(P1_P1_InstAddrPointer_PTR12), .B(_01998__PTR12), .S(_01853__PTR3), .Z(_02084__PTR204) );
  MUX2_X1 U6055 ( .A(P1_P1_InstAddrPointer_PTR13), .B(_01998__PTR13), .S(_01853__PTR3), .Z(_02084__PTR205) );
  MUX2_X1 U6056 ( .A(P1_P1_InstAddrPointer_PTR14), .B(_01998__PTR14), .S(_01853__PTR3), .Z(_02084__PTR206) );
  MUX2_X1 U6057 ( .A(P1_P1_InstAddrPointer_PTR15), .B(_01998__PTR15), .S(_01853__PTR3), .Z(_02084__PTR207) );
  MUX2_X1 U6058 ( .A(P1_P1_InstAddrPointer_PTR16), .B(_01998__PTR16), .S(_01853__PTR3), .Z(_02084__PTR208) );
  MUX2_X1 U6059 ( .A(P1_P1_InstAddrPointer_PTR17), .B(_01998__PTR17), .S(_01853__PTR3), .Z(_02084__PTR209) );
  MUX2_X1 U6060 ( .A(P1_P1_InstAddrPointer_PTR18), .B(_01998__PTR18), .S(_01853__PTR3), .Z(_02084__PTR210) );
  MUX2_X1 U6061 ( .A(P1_P1_InstAddrPointer_PTR19), .B(_01998__PTR19), .S(_01853__PTR3), .Z(_02084__PTR211) );
  MUX2_X1 U6062 ( .A(P1_P1_InstAddrPointer_PTR20), .B(_01998__PTR20), .S(_01853__PTR3), .Z(_02084__PTR212) );
  MUX2_X1 U6063 ( .A(P1_P1_InstAddrPointer_PTR21), .B(_01998__PTR21), .S(_01853__PTR3), .Z(_02084__PTR213) );
  MUX2_X1 U6064 ( .A(P1_P1_InstAddrPointer_PTR22), .B(_01998__PTR22), .S(_01853__PTR3), .Z(_02084__PTR214) );
  MUX2_X1 U6065 ( .A(P1_P1_InstAddrPointer_PTR23), .B(_01998__PTR23), .S(_01853__PTR3), .Z(_02084__PTR215) );
  MUX2_X1 U6066 ( .A(P1_P1_InstAddrPointer_PTR24), .B(_01998__PTR24), .S(_01853__PTR3), .Z(_02084__PTR216) );
  MUX2_X1 U6067 ( .A(P1_P1_InstAddrPointer_PTR25), .B(_01998__PTR25), .S(_01853__PTR3), .Z(_02084__PTR217) );
  MUX2_X1 U6068 ( .A(P1_P1_InstAddrPointer_PTR26), .B(_01998__PTR26), .S(_01853__PTR3), .Z(_02084__PTR218) );
  MUX2_X1 U6069 ( .A(P1_P1_InstAddrPointer_PTR27), .B(_01998__PTR27), .S(_01853__PTR3), .Z(_02084__PTR219) );
  MUX2_X1 U6070 ( .A(P1_P1_InstAddrPointer_PTR28), .B(_01998__PTR28), .S(_01853__PTR3), .Z(_02084__PTR220) );
  MUX2_X1 U6071 ( .A(P1_P1_InstAddrPointer_PTR29), .B(_01998__PTR29), .S(_01853__PTR3), .Z(_02084__PTR221) );
  MUX2_X1 U6072 ( .A(P1_P1_InstAddrPointer_PTR30), .B(_01998__PTR30), .S(_01853__PTR3), .Z(_02084__PTR222) );
  MUX2_X1 U6073 ( .A(P1_P1_InstAddrPointer_PTR31), .B(_01998__PTR31), .S(_01853__PTR3), .Z(_02084__PTR223) );
  MUX2_X1 U6074 ( .A(P1_P1_PhyAddrPointer_PTR0), .B(_01998__PTR0), .S(_01853__PTR3), .Z(_02092__PTR64) );
  MUX2_X1 U6075 ( .A(P1_P1_PhyAddrPointer_PTR1), .B(_01998__PTR1), .S(_01853__PTR3), .Z(_02092__PTR65) );
  MUX2_X1 U6076 ( .A(P1_P1_PhyAddrPointer_PTR2), .B(_01998__PTR2), .S(_01853__PTR3), .Z(_02092__PTR66) );
  MUX2_X1 U6077 ( .A(P1_P1_PhyAddrPointer_PTR3), .B(_01998__PTR3), .S(_01853__PTR3), .Z(_02092__PTR67) );
  MUX2_X1 U6078 ( .A(P1_P1_PhyAddrPointer_PTR4), .B(_01998__PTR4), .S(_01853__PTR3), .Z(_02092__PTR68) );
  MUX2_X1 U6079 ( .A(P1_P1_PhyAddrPointer_PTR5), .B(_01998__PTR5), .S(_01853__PTR3), .Z(_02092__PTR69) );
  MUX2_X1 U6080 ( .A(P1_P1_PhyAddrPointer_PTR6), .B(_01998__PTR6), .S(_01853__PTR3), .Z(_02092__PTR70) );
  MUX2_X1 U6081 ( .A(P1_P1_PhyAddrPointer_PTR7), .B(_01998__PTR7), .S(_01853__PTR3), .Z(_02092__PTR71) );
  MUX2_X1 U6082 ( .A(P1_P1_PhyAddrPointer_PTR8), .B(_01998__PTR8), .S(_01853__PTR3), .Z(_02092__PTR72) );
  MUX2_X1 U6083 ( .A(P1_P1_PhyAddrPointer_PTR9), .B(_01998__PTR9), .S(_01853__PTR3), .Z(_02092__PTR73) );
  MUX2_X1 U6084 ( .A(P1_P1_PhyAddrPointer_PTR10), .B(_01998__PTR10), .S(_01853__PTR3), .Z(_02092__PTR74) );
  MUX2_X1 U6085 ( .A(P1_P1_PhyAddrPointer_PTR11), .B(_01998__PTR11), .S(_01853__PTR3), .Z(_02092__PTR75) );
  MUX2_X1 U6086 ( .A(P1_P1_PhyAddrPointer_PTR12), .B(_01998__PTR12), .S(_01853__PTR3), .Z(_02092__PTR76) );
  MUX2_X1 U6087 ( .A(P1_P1_PhyAddrPointer_PTR13), .B(_01998__PTR13), .S(_01853__PTR3), .Z(_02092__PTR77) );
  MUX2_X1 U6088 ( .A(P1_P1_PhyAddrPointer_PTR14), .B(_01998__PTR14), .S(_01853__PTR3), .Z(_02092__PTR78) );
  MUX2_X1 U6089 ( .A(P1_P1_PhyAddrPointer_PTR15), .B(_01998__PTR15), .S(_01853__PTR3), .Z(_02092__PTR79) );
  MUX2_X1 U6090 ( .A(P1_P1_PhyAddrPointer_PTR16), .B(_01998__PTR16), .S(_01853__PTR3), .Z(_02092__PTR80) );
  MUX2_X1 U6091 ( .A(P1_P1_PhyAddrPointer_PTR17), .B(_01998__PTR17), .S(_01853__PTR3), .Z(_02092__PTR81) );
  MUX2_X1 U6092 ( .A(P1_P1_PhyAddrPointer_PTR18), .B(_01998__PTR18), .S(_01853__PTR3), .Z(_02092__PTR82) );
  MUX2_X1 U6093 ( .A(P1_P1_PhyAddrPointer_PTR19), .B(_01998__PTR19), .S(_01853__PTR3), .Z(_02092__PTR83) );
  MUX2_X1 U6094 ( .A(P1_P1_PhyAddrPointer_PTR20), .B(_01998__PTR20), .S(_01853__PTR3), .Z(_02092__PTR84) );
  MUX2_X1 U6095 ( .A(P1_P1_PhyAddrPointer_PTR21), .B(_01998__PTR21), .S(_01853__PTR3), .Z(_02092__PTR85) );
  MUX2_X1 U6096 ( .A(P1_P1_PhyAddrPointer_PTR22), .B(_01998__PTR22), .S(_01853__PTR3), .Z(_02092__PTR86) );
  MUX2_X1 U6097 ( .A(P1_P1_PhyAddrPointer_PTR23), .B(_01998__PTR23), .S(_01853__PTR3), .Z(_02092__PTR87) );
  MUX2_X1 U6098 ( .A(P1_P1_PhyAddrPointer_PTR24), .B(_01998__PTR24), .S(_01853__PTR3), .Z(_02092__PTR88) );
  MUX2_X1 U6099 ( .A(P1_P1_PhyAddrPointer_PTR25), .B(_01998__PTR25), .S(_01853__PTR3), .Z(_02092__PTR89) );
  MUX2_X1 U6100 ( .A(P1_P1_PhyAddrPointer_PTR26), .B(_01998__PTR26), .S(_01853__PTR3), .Z(_02092__PTR90) );
  MUX2_X1 U6101 ( .A(P1_P1_PhyAddrPointer_PTR27), .B(_01998__PTR27), .S(_01853__PTR3), .Z(_02092__PTR91) );
  MUX2_X1 U6102 ( .A(P1_P1_PhyAddrPointer_PTR28), .B(_01998__PTR28), .S(_01853__PTR3), .Z(_02092__PTR92) );
  MUX2_X1 U6103 ( .A(P1_P1_PhyAddrPointer_PTR29), .B(_01998__PTR29), .S(_01853__PTR3), .Z(_02092__PTR93) );
  MUX2_X1 U6104 ( .A(P1_P1_PhyAddrPointer_PTR30), .B(_01998__PTR30), .S(_01853__PTR3), .Z(_02092__PTR94) );
  MUX2_X1 U6105 ( .A(P1_P1_PhyAddrPointer_PTR31), .B(_01998__PTR31), .S(_01853__PTR3), .Z(_02092__PTR95) );
  MUX2_X1 U6106 ( .A(_02939__PTR0), .B(_02803__PTR0), .S(_02724__PTR7), .Z(_01998__PTR0) );
  MUX2_X1 U6107 ( .A(_02939__PTR1), .B(_02804__PTR1), .S(_02724__PTR7), .Z(_01998__PTR1) );
  MUX2_X1 U6108 ( .A(_02939__PTR2), .B(_02804__PTR2), .S(_02724__PTR7), .Z(_01998__PTR2) );
  MUX2_X1 U6109 ( .A(_02939__PTR3), .B(_02804__PTR3), .S(_02724__PTR7), .Z(_01998__PTR3) );
  MUX2_X1 U6110 ( .A(_02939__PTR4), .B(_02804__PTR4), .S(_02724__PTR7), .Z(_01998__PTR4) );
  MUX2_X1 U6111 ( .A(_02939__PTR5), .B(_02804__PTR5), .S(_02724__PTR7), .Z(_01998__PTR5) );
  MUX2_X1 U6112 ( .A(_02939__PTR6), .B(_02804__PTR6), .S(_02724__PTR7), .Z(_01998__PTR6) );
  MUX2_X1 U6113 ( .A(_02939__PTR7), .B(_02804__PTR7), .S(_02724__PTR7), .Z(_01998__PTR7) );
  MUX2_X1 U6114 ( .A(_02939__PTR8), .B(_02804__PTR8), .S(_02724__PTR7), .Z(_01998__PTR8) );
  MUX2_X1 U6115 ( .A(_02939__PTR9), .B(_02804__PTR9), .S(_02724__PTR7), .Z(_01998__PTR9) );
  MUX2_X1 U6116 ( .A(_02939__PTR10), .B(_02804__PTR10), .S(_02724__PTR7), .Z(_01998__PTR10) );
  MUX2_X1 U6117 ( .A(_02939__PTR11), .B(_02804__PTR11), .S(_02724__PTR7), .Z(_01998__PTR11) );
  MUX2_X1 U6118 ( .A(_02939__PTR12), .B(_02804__PTR12), .S(_02724__PTR7), .Z(_01998__PTR12) );
  MUX2_X1 U6119 ( .A(_02939__PTR13), .B(_02804__PTR13), .S(_02724__PTR7), .Z(_01998__PTR13) );
  MUX2_X1 U6120 ( .A(_02939__PTR14), .B(_02804__PTR14), .S(_02724__PTR7), .Z(_01998__PTR14) );
  MUX2_X1 U6121 ( .A(_02939__PTR15), .B(_02804__PTR15), .S(_02724__PTR7), .Z(_01998__PTR15) );
  MUX2_X1 U6122 ( .A(_02939__PTR16), .B(_02804__PTR16), .S(_02724__PTR7), .Z(_01998__PTR16) );
  MUX2_X1 U6123 ( .A(_02939__PTR17), .B(_02804__PTR17), .S(_02724__PTR7), .Z(_01998__PTR17) );
  MUX2_X1 U6124 ( .A(_02939__PTR18), .B(_02804__PTR18), .S(_02724__PTR7), .Z(_01998__PTR18) );
  MUX2_X1 U6125 ( .A(_02939__PTR19), .B(_02804__PTR19), .S(_02724__PTR7), .Z(_01998__PTR19) );
  MUX2_X1 U6126 ( .A(_02939__PTR20), .B(_02804__PTR20), .S(_02724__PTR7), .Z(_01998__PTR20) );
  MUX2_X1 U6127 ( .A(_02939__PTR21), .B(_02804__PTR21), .S(_02724__PTR7), .Z(_01998__PTR21) );
  MUX2_X1 U6128 ( .A(_02939__PTR22), .B(_02804__PTR22), .S(_02724__PTR7), .Z(_01998__PTR22) );
  MUX2_X1 U6129 ( .A(_02939__PTR23), .B(_02804__PTR23), .S(_02724__PTR7), .Z(_01998__PTR23) );
  MUX2_X1 U6130 ( .A(_02939__PTR24), .B(_02804__PTR24), .S(_02724__PTR7), .Z(_01998__PTR24) );
  MUX2_X1 U6131 ( .A(_02939__PTR25), .B(_02804__PTR25), .S(_02724__PTR7), .Z(_01998__PTR25) );
  MUX2_X1 U6132 ( .A(_02939__PTR26), .B(_02804__PTR26), .S(_02724__PTR7), .Z(_01998__PTR26) );
  MUX2_X1 U6133 ( .A(_02939__PTR27), .B(_02804__PTR27), .S(_02724__PTR7), .Z(_01998__PTR27) );
  MUX2_X1 U6134 ( .A(_02939__PTR28), .B(_02804__PTR28), .S(_02724__PTR7), .Z(_01998__PTR28) );
  MUX2_X1 U6135 ( .A(_02939__PTR29), .B(_02804__PTR29), .S(_02724__PTR7), .Z(_01998__PTR29) );
  MUX2_X1 U6136 ( .A(_02939__PTR30), .B(_02804__PTR30), .S(_02724__PTR7), .Z(_01998__PTR30) );
  MUX2_X1 U6137 ( .A(_02939__PTR31), .B(_02804__PTR31), .S(_02724__PTR7), .Z(_01998__PTR31) );
  MUX2_X1 U6138 ( .A(P1_P1_PhyAddrPointer_PTR0), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR128) );
  MUX2_X1 U6139 ( .A(_01996__PTR1), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR129) );
  MUX2_X1 U6140 ( .A(_01996__PTR2), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR130) );
  MUX2_X1 U6141 ( .A(_01996__PTR3), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR131) );
  MUX2_X1 U6142 ( .A(_01996__PTR4), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR132) );
  MUX2_X1 U6143 ( .A(_01996__PTR5), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR133) );
  MUX2_X1 U6144 ( .A(_01996__PTR6), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR134) );
  MUX2_X1 U6145 ( .A(_01996__PTR7), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR135) );
  MUX2_X1 U6146 ( .A(_01996__PTR8), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR136) );
  MUX2_X1 U6147 ( .A(_01996__PTR9), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR137) );
  MUX2_X1 U6148 ( .A(_01996__PTR10), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR138) );
  MUX2_X1 U6149 ( .A(_01996__PTR11), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR139) );
  MUX2_X1 U6150 ( .A(_01996__PTR12), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR140) );
  MUX2_X1 U6151 ( .A(_01996__PTR13), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR141) );
  MUX2_X1 U6152 ( .A(_01996__PTR14), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR142) );
  MUX2_X1 U6153 ( .A(_01996__PTR15), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR143) );
  MUX2_X1 U6154 ( .A(_01996__PTR16), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR144) );
  MUX2_X1 U6155 ( .A(_01996__PTR17), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR145) );
  MUX2_X1 U6156 ( .A(_01996__PTR18), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR146) );
  MUX2_X1 U6157 ( .A(_01996__PTR19), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR147) );
  MUX2_X1 U6158 ( .A(_01996__PTR20), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR148) );
  MUX2_X1 U6159 ( .A(_01996__PTR21), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR149) );
  MUX2_X1 U6160 ( .A(_01996__PTR22), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR150) );
  MUX2_X1 U6161 ( .A(_01996__PTR23), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR151) );
  MUX2_X1 U6162 ( .A(_01996__PTR24), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR152) );
  MUX2_X1 U6163 ( .A(_01996__PTR25), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR153) );
  MUX2_X1 U6164 ( .A(_01996__PTR26), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR154) );
  MUX2_X1 U6165 ( .A(_01996__PTR27), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR155) );
  MUX2_X1 U6166 ( .A(_01996__PTR28), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR156) );
  MUX2_X1 U6167 ( .A(_01996__PTR29), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR157) );
  MUX2_X1 U6168 ( .A(_01996__PTR30), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR158) );
  MUX2_X1 U6169 ( .A(_01996__PTR31), .B(1'b0), .S(P1_StateBS16), .Z(_01896__PTR160) );
  MUX2_X1 U6170 ( .A(_01892__PTR129), .B(1'b0), .S(P1_StateBS16), .Z(_01892__PTR65) );
  MUX2_X1 U6171 ( .A(_01892__PTR130), .B(_02795__PTR0), .S(P1_StateBS16), .Z(_01892__PTR66) );
  MUX2_X1 U6172 ( .A(_01892__PTR131), .B(_02796__PTR1), .S(P1_StateBS16), .Z(_01892__PTR67) );
  MUX2_X1 U6173 ( .A(_01892__PTR132), .B(_02796__PTR2), .S(P1_StateBS16), .Z(_01892__PTR68) );
  MUX2_X1 U6174 ( .A(_01892__PTR133), .B(_02796__PTR3), .S(P1_StateBS16), .Z(_01892__PTR69) );
  MUX2_X1 U6175 ( .A(_01892__PTR134), .B(_02796__PTR4), .S(P1_StateBS16), .Z(_01892__PTR70) );
  MUX2_X1 U6176 ( .A(_01892__PTR135), .B(_02796__PTR5), .S(P1_StateBS16), .Z(_01892__PTR71) );
  MUX2_X1 U6177 ( .A(_01892__PTR136), .B(_02796__PTR6), .S(P1_StateBS16), .Z(_01892__PTR72) );
  MUX2_X1 U6178 ( .A(_01892__PTR137), .B(_02796__PTR7), .S(P1_StateBS16), .Z(_01892__PTR73) );
  MUX2_X1 U6179 ( .A(_01892__PTR138), .B(_02796__PTR8), .S(P1_StateBS16), .Z(_01892__PTR74) );
  MUX2_X1 U6180 ( .A(_01892__PTR139), .B(_02796__PTR9), .S(P1_StateBS16), .Z(_01892__PTR75) );
  MUX2_X1 U6181 ( .A(_01892__PTR140), .B(_02796__PTR10), .S(P1_StateBS16), .Z(_01892__PTR76) );
  MUX2_X1 U6182 ( .A(_01892__PTR141), .B(_02796__PTR11), .S(P1_StateBS16), .Z(_01892__PTR77) );
  MUX2_X1 U6183 ( .A(_01892__PTR142), .B(_02796__PTR12), .S(P1_StateBS16), .Z(_01892__PTR78) );
  MUX2_X1 U6184 ( .A(_01892__PTR143), .B(_02796__PTR13), .S(P1_StateBS16), .Z(_01892__PTR79) );
  MUX2_X1 U6185 ( .A(_01892__PTR144), .B(_02796__PTR14), .S(P1_StateBS16), .Z(_01892__PTR80) );
  MUX2_X1 U6186 ( .A(_01892__PTR145), .B(_02796__PTR15), .S(P1_StateBS16), .Z(_01892__PTR81) );
  MUX2_X1 U6187 ( .A(_01892__PTR146), .B(_02796__PTR16), .S(P1_StateBS16), .Z(_01892__PTR82) );
  MUX2_X1 U6188 ( .A(_01892__PTR147), .B(_02796__PTR17), .S(P1_StateBS16), .Z(_01892__PTR83) );
  MUX2_X1 U6189 ( .A(_01892__PTR148), .B(_02796__PTR18), .S(P1_StateBS16), .Z(_01892__PTR84) );
  MUX2_X1 U6190 ( .A(_01892__PTR149), .B(_02796__PTR19), .S(P1_StateBS16), .Z(_01892__PTR85) );
  MUX2_X1 U6191 ( .A(_01892__PTR150), .B(_02796__PTR20), .S(P1_StateBS16), .Z(_01892__PTR86) );
  MUX2_X1 U6192 ( .A(_01892__PTR151), .B(_02796__PTR21), .S(P1_StateBS16), .Z(_01892__PTR87) );
  MUX2_X1 U6193 ( .A(_01892__PTR152), .B(_02796__PTR22), .S(P1_StateBS16), .Z(_01892__PTR88) );
  MUX2_X1 U6194 ( .A(_01892__PTR153), .B(_02796__PTR23), .S(P1_StateBS16), .Z(_01892__PTR89) );
  MUX2_X1 U6195 ( .A(_01892__PTR154), .B(_02796__PTR24), .S(P1_StateBS16), .Z(_01892__PTR90) );
  MUX2_X1 U6196 ( .A(_01892__PTR155), .B(_02796__PTR25), .S(P1_StateBS16), .Z(_01892__PTR91) );
  MUX2_X1 U6197 ( .A(_01892__PTR156), .B(_02796__PTR26), .S(P1_StateBS16), .Z(_01892__PTR92) );
  MUX2_X1 U6198 ( .A(_01892__PTR157), .B(_02796__PTR27), .S(P1_StateBS16), .Z(_01892__PTR93) );
  MUX2_X1 U6199 ( .A(_01892__PTR158), .B(_02796__PTR28), .S(P1_StateBS16), .Z(_01892__PTR94) );
  MUX2_X1 U6200 ( .A(_01892__PTR159), .B(_02796__PTR29), .S(P1_StateBS16), .Z(_01892__PTR95) );
  MUX2_X1 U6201 ( .A(_01838__PTR1), .B(_02791__PTR1), .S(P1_StateBS16), .Z(_01930__PTR17) );
  MUX2_X1 U6202 ( .A(_01838__PTR2), .B(_02791__PTR2), .S(P1_StateBS16), .Z(_01930__PTR18) );
  MUX2_X1 U6203 ( .A(_01838__PTR3), .B(_02791__PTR3), .S(P1_StateBS16), .Z(_01930__PTR19) );
  MUX2_X1 U6204 ( .A(_01928__PTR32), .B(_01995__PTR0), .S(P1_StateBS16), .Z(_01928__PTR16) );
  MUX2_X1 U6205 ( .A(_01928__PTR33), .B(_01995__PTR1), .S(P1_StateBS16), .Z(_01928__PTR17) );
  MUX2_X1 U6206 ( .A(_01928__PTR34), .B(_01995__PTR2), .S(P1_StateBS16), .Z(_01928__PTR18) );
  MUX2_X1 U6207 ( .A(_01928__PTR35), .B(_01995__PTR3), .S(P1_StateBS16), .Z(_01928__PTR19) );
  MUX2_X1 U6208 ( .A(_01928__PTR36), .B(_01995__PTR4), .S(P1_StateBS16), .Z(_01928__PTR20) );
  MUX2_X1 U6209 ( .A(_01928__PTR37), .B(_01995__PTR5), .S(P1_StateBS16), .Z(_01928__PTR21) );
  MUX2_X1 U6210 ( .A(_01928__PTR38), .B(_01995__PTR6), .S(P1_StateBS16), .Z(_01928__PTR22) );
  MUX2_X1 U6211 ( .A(_01928__PTR39), .B(_01995__PTR7), .S(P1_StateBS16), .Z(_01928__PTR23) );
  MUX2_X1 U6212 ( .A(_01926__PTR32), .B(_01994__PTR0), .S(P1_StateBS16), .Z(_01926__PTR16) );
  MUX2_X1 U6213 ( .A(_01926__PTR33), .B(_01994__PTR1), .S(P1_StateBS16), .Z(_01926__PTR17) );
  MUX2_X1 U6214 ( .A(_01926__PTR34), .B(_01994__PTR2), .S(P1_StateBS16), .Z(_01926__PTR18) );
  MUX2_X1 U6215 ( .A(_01926__PTR35), .B(_01994__PTR3), .S(P1_StateBS16), .Z(_01926__PTR19) );
  MUX2_X1 U6216 ( .A(_01926__PTR36), .B(_01994__PTR4), .S(P1_StateBS16), .Z(_01926__PTR20) );
  MUX2_X1 U6217 ( .A(_01926__PTR37), .B(_01994__PTR5), .S(P1_StateBS16), .Z(_01926__PTR21) );
  MUX2_X1 U6218 ( .A(_01926__PTR38), .B(_01994__PTR6), .S(P1_StateBS16), .Z(_01926__PTR22) );
  MUX2_X1 U6219 ( .A(_01926__PTR39), .B(_01994__PTR7), .S(P1_StateBS16), .Z(_01926__PTR23) );
  MUX2_X1 U6220 ( .A(_01924__PTR32), .B(_01993__PTR0), .S(P1_StateBS16), .Z(_01924__PTR16) );
  MUX2_X1 U6221 ( .A(_01924__PTR33), .B(_01993__PTR1), .S(P1_StateBS16), .Z(_01924__PTR17) );
  MUX2_X1 U6222 ( .A(_01924__PTR34), .B(_01993__PTR2), .S(P1_StateBS16), .Z(_01924__PTR18) );
  MUX2_X1 U6223 ( .A(_01924__PTR35), .B(_01993__PTR3), .S(P1_StateBS16), .Z(_01924__PTR19) );
  MUX2_X1 U6224 ( .A(_01924__PTR36), .B(_01993__PTR4), .S(P1_StateBS16), .Z(_01924__PTR20) );
  MUX2_X1 U6225 ( .A(_01924__PTR37), .B(_01993__PTR5), .S(P1_StateBS16), .Z(_01924__PTR21) );
  MUX2_X1 U6226 ( .A(_01924__PTR38), .B(_01993__PTR6), .S(P1_StateBS16), .Z(_01924__PTR22) );
  MUX2_X1 U6227 ( .A(_01924__PTR39), .B(_01993__PTR7), .S(P1_StateBS16), .Z(_01924__PTR23) );
  MUX2_X1 U6228 ( .A(_01922__PTR32), .B(_01992__PTR0), .S(P1_StateBS16), .Z(_01922__PTR16) );
  MUX2_X1 U6229 ( .A(_01922__PTR33), .B(_01992__PTR1), .S(P1_StateBS16), .Z(_01922__PTR17) );
  MUX2_X1 U6230 ( .A(_01922__PTR34), .B(_01992__PTR2), .S(P1_StateBS16), .Z(_01922__PTR18) );
  MUX2_X1 U6231 ( .A(_01922__PTR35), .B(_01992__PTR3), .S(P1_StateBS16), .Z(_01922__PTR19) );
  MUX2_X1 U6232 ( .A(_01922__PTR36), .B(_01992__PTR4), .S(P1_StateBS16), .Z(_01922__PTR20) );
  MUX2_X1 U6233 ( .A(_01922__PTR37), .B(_01992__PTR5), .S(P1_StateBS16), .Z(_01922__PTR21) );
  MUX2_X1 U6234 ( .A(_01922__PTR38), .B(_01992__PTR6), .S(P1_StateBS16), .Z(_01922__PTR22) );
  MUX2_X1 U6235 ( .A(_01922__PTR39), .B(_01992__PTR7), .S(P1_StateBS16), .Z(_01922__PTR23) );
  MUX2_X1 U6236 ( .A(_01920__PTR32), .B(_01991__PTR0), .S(P1_StateBS16), .Z(_01920__PTR16) );
  MUX2_X1 U6237 ( .A(_01920__PTR33), .B(_01991__PTR1), .S(P1_StateBS16), .Z(_01920__PTR17) );
  MUX2_X1 U6238 ( .A(_01920__PTR34), .B(_01991__PTR2), .S(P1_StateBS16), .Z(_01920__PTR18) );
  MUX2_X1 U6239 ( .A(_01920__PTR35), .B(_01991__PTR3), .S(P1_StateBS16), .Z(_01920__PTR19) );
  MUX2_X1 U6240 ( .A(_01920__PTR36), .B(_01991__PTR4), .S(P1_StateBS16), .Z(_01920__PTR20) );
  MUX2_X1 U6241 ( .A(_01920__PTR37), .B(_01991__PTR5), .S(P1_StateBS16), .Z(_01920__PTR21) );
  MUX2_X1 U6242 ( .A(_01920__PTR38), .B(_01991__PTR6), .S(P1_StateBS16), .Z(_01920__PTR22) );
  MUX2_X1 U6243 ( .A(_01920__PTR39), .B(_01991__PTR7), .S(P1_StateBS16), .Z(_01920__PTR23) );
  MUX2_X1 U6244 ( .A(_01918__PTR32), .B(_01990__PTR0), .S(P1_StateBS16), .Z(_01918__PTR16) );
  MUX2_X1 U6245 ( .A(_01918__PTR33), .B(_01990__PTR1), .S(P1_StateBS16), .Z(_01918__PTR17) );
  MUX2_X1 U6246 ( .A(_01918__PTR34), .B(_01990__PTR2), .S(P1_StateBS16), .Z(_01918__PTR18) );
  MUX2_X1 U6247 ( .A(_01918__PTR35), .B(_01990__PTR3), .S(P1_StateBS16), .Z(_01918__PTR19) );
  MUX2_X1 U6248 ( .A(_01918__PTR36), .B(_01990__PTR4), .S(P1_StateBS16), .Z(_01918__PTR20) );
  MUX2_X1 U6249 ( .A(_01918__PTR37), .B(_01990__PTR5), .S(P1_StateBS16), .Z(_01918__PTR21) );
  MUX2_X1 U6250 ( .A(_01918__PTR38), .B(_01990__PTR6), .S(P1_StateBS16), .Z(_01918__PTR22) );
  MUX2_X1 U6251 ( .A(_01918__PTR39), .B(_01990__PTR7), .S(P1_StateBS16), .Z(_01918__PTR23) );
  MUX2_X1 U6252 ( .A(_01916__PTR32), .B(_01989__PTR0), .S(P1_StateBS16), .Z(_01916__PTR16) );
  MUX2_X1 U6253 ( .A(_01916__PTR33), .B(_01989__PTR1), .S(P1_StateBS16), .Z(_01916__PTR17) );
  MUX2_X1 U6254 ( .A(_01916__PTR34), .B(_01989__PTR2), .S(P1_StateBS16), .Z(_01916__PTR18) );
  MUX2_X1 U6255 ( .A(_01916__PTR35), .B(_01989__PTR3), .S(P1_StateBS16), .Z(_01916__PTR19) );
  MUX2_X1 U6256 ( .A(_01916__PTR36), .B(_01989__PTR4), .S(P1_StateBS16), .Z(_01916__PTR20) );
  MUX2_X1 U6257 ( .A(_01916__PTR37), .B(_01989__PTR5), .S(P1_StateBS16), .Z(_01916__PTR21) );
  MUX2_X1 U6258 ( .A(_01916__PTR38), .B(_01989__PTR6), .S(P1_StateBS16), .Z(_01916__PTR22) );
  MUX2_X1 U6259 ( .A(_01916__PTR39), .B(_01989__PTR7), .S(P1_StateBS16), .Z(_01916__PTR23) );
  MUX2_X1 U6260 ( .A(_01914__PTR32), .B(_01988__PTR0), .S(P1_StateBS16), .Z(_01914__PTR16) );
  MUX2_X1 U6261 ( .A(_01914__PTR33), .B(_01988__PTR1), .S(P1_StateBS16), .Z(_01914__PTR17) );
  MUX2_X1 U6262 ( .A(_01914__PTR34), .B(_01988__PTR2), .S(P1_StateBS16), .Z(_01914__PTR18) );
  MUX2_X1 U6263 ( .A(_01914__PTR35), .B(_01988__PTR3), .S(P1_StateBS16), .Z(_01914__PTR19) );
  MUX2_X1 U6264 ( .A(_01914__PTR36), .B(_01988__PTR4), .S(P1_StateBS16), .Z(_01914__PTR20) );
  MUX2_X1 U6265 ( .A(_01914__PTR37), .B(_01988__PTR5), .S(P1_StateBS16), .Z(_01914__PTR21) );
  MUX2_X1 U6266 ( .A(_01914__PTR38), .B(_01988__PTR6), .S(P1_StateBS16), .Z(_01914__PTR22) );
  MUX2_X1 U6267 ( .A(_01914__PTR39), .B(_01988__PTR7), .S(P1_StateBS16), .Z(_01914__PTR23) );
  MUX2_X1 U6268 ( .A(_01912__PTR32), .B(_01987__PTR0), .S(P1_StateBS16), .Z(_01912__PTR16) );
  MUX2_X1 U6269 ( .A(_01912__PTR33), .B(_01987__PTR1), .S(P1_StateBS16), .Z(_01912__PTR17) );
  MUX2_X1 U6270 ( .A(_01912__PTR34), .B(_01987__PTR2), .S(P1_StateBS16), .Z(_01912__PTR18) );
  MUX2_X1 U6271 ( .A(_01912__PTR35), .B(_01987__PTR3), .S(P1_StateBS16), .Z(_01912__PTR19) );
  MUX2_X1 U6272 ( .A(_01912__PTR36), .B(_01987__PTR4), .S(P1_StateBS16), .Z(_01912__PTR20) );
  MUX2_X1 U6273 ( .A(_01912__PTR37), .B(_01987__PTR5), .S(P1_StateBS16), .Z(_01912__PTR21) );
  MUX2_X1 U6274 ( .A(_01912__PTR38), .B(_01987__PTR6), .S(P1_StateBS16), .Z(_01912__PTR22) );
  MUX2_X1 U6275 ( .A(_01912__PTR39), .B(_01987__PTR7), .S(P1_StateBS16), .Z(_01912__PTR23) );
  MUX2_X1 U6276 ( .A(_01910__PTR32), .B(_01986__PTR0), .S(P1_StateBS16), .Z(_01910__PTR16) );
  MUX2_X1 U6277 ( .A(_01910__PTR33), .B(_01986__PTR1), .S(P1_StateBS16), .Z(_01910__PTR17) );
  MUX2_X1 U6278 ( .A(_01910__PTR34), .B(_01986__PTR2), .S(P1_StateBS16), .Z(_01910__PTR18) );
  MUX2_X1 U6279 ( .A(_01910__PTR35), .B(_01986__PTR3), .S(P1_StateBS16), .Z(_01910__PTR19) );
  MUX2_X1 U6280 ( .A(_01910__PTR36), .B(_01986__PTR4), .S(P1_StateBS16), .Z(_01910__PTR20) );
  MUX2_X1 U6281 ( .A(_01910__PTR37), .B(_01986__PTR5), .S(P1_StateBS16), .Z(_01910__PTR21) );
  MUX2_X1 U6282 ( .A(_01910__PTR38), .B(_01986__PTR6), .S(P1_StateBS16), .Z(_01910__PTR22) );
  MUX2_X1 U6283 ( .A(_01910__PTR39), .B(_01986__PTR7), .S(P1_StateBS16), .Z(_01910__PTR23) );
  MUX2_X1 U6284 ( .A(_01908__PTR32), .B(_01985__PTR0), .S(P1_StateBS16), .Z(_01908__PTR16) );
  MUX2_X1 U6285 ( .A(_01908__PTR33), .B(_01985__PTR1), .S(P1_StateBS16), .Z(_01908__PTR17) );
  MUX2_X1 U6286 ( .A(_01908__PTR34), .B(_01985__PTR2), .S(P1_StateBS16), .Z(_01908__PTR18) );
  MUX2_X1 U6287 ( .A(_01908__PTR35), .B(_01985__PTR3), .S(P1_StateBS16), .Z(_01908__PTR19) );
  MUX2_X1 U6288 ( .A(_01908__PTR36), .B(_01985__PTR4), .S(P1_StateBS16), .Z(_01908__PTR20) );
  MUX2_X1 U6289 ( .A(_01908__PTR37), .B(_01985__PTR5), .S(P1_StateBS16), .Z(_01908__PTR21) );
  MUX2_X1 U6290 ( .A(_01908__PTR38), .B(_01985__PTR6), .S(P1_StateBS16), .Z(_01908__PTR22) );
  MUX2_X1 U6291 ( .A(_01908__PTR39), .B(_01985__PTR7), .S(P1_StateBS16), .Z(_01908__PTR23) );
  MUX2_X1 U6292 ( .A(_01906__PTR32), .B(_01984__PTR0), .S(P1_StateBS16), .Z(_01906__PTR16) );
  MUX2_X1 U6293 ( .A(_01906__PTR33), .B(_01984__PTR1), .S(P1_StateBS16), .Z(_01906__PTR17) );
  MUX2_X1 U6294 ( .A(_01906__PTR34), .B(_01984__PTR2), .S(P1_StateBS16), .Z(_01906__PTR18) );
  MUX2_X1 U6295 ( .A(_01906__PTR35), .B(_01984__PTR3), .S(P1_StateBS16), .Z(_01906__PTR19) );
  MUX2_X1 U6296 ( .A(_01906__PTR36), .B(_01984__PTR4), .S(P1_StateBS16), .Z(_01906__PTR20) );
  MUX2_X1 U6297 ( .A(_01906__PTR37), .B(_01984__PTR5), .S(P1_StateBS16), .Z(_01906__PTR21) );
  MUX2_X1 U6298 ( .A(_01906__PTR38), .B(_01984__PTR6), .S(P1_StateBS16), .Z(_01906__PTR22) );
  MUX2_X1 U6299 ( .A(_01906__PTR39), .B(_01984__PTR7), .S(P1_StateBS16), .Z(_01906__PTR23) );
  MUX2_X1 U6300 ( .A(_01904__PTR32), .B(_01983__PTR0), .S(P1_StateBS16), .Z(_01904__PTR16) );
  MUX2_X1 U6301 ( .A(_01904__PTR33), .B(_01983__PTR1), .S(P1_StateBS16), .Z(_01904__PTR17) );
  MUX2_X1 U6302 ( .A(_01904__PTR34), .B(_01983__PTR2), .S(P1_StateBS16), .Z(_01904__PTR18) );
  MUX2_X1 U6303 ( .A(_01904__PTR35), .B(_01983__PTR3), .S(P1_StateBS16), .Z(_01904__PTR19) );
  MUX2_X1 U6304 ( .A(_01904__PTR36), .B(_01983__PTR4), .S(P1_StateBS16), .Z(_01904__PTR20) );
  MUX2_X1 U6305 ( .A(_01904__PTR37), .B(_01983__PTR5), .S(P1_StateBS16), .Z(_01904__PTR21) );
  MUX2_X1 U6306 ( .A(_01904__PTR38), .B(_01983__PTR6), .S(P1_StateBS16), .Z(_01904__PTR22) );
  MUX2_X1 U6307 ( .A(_01904__PTR39), .B(_01983__PTR7), .S(P1_StateBS16), .Z(_01904__PTR23) );
  MUX2_X1 U6308 ( .A(_01902__PTR32), .B(_01982__PTR0), .S(P1_StateBS16), .Z(_01902__PTR16) );
  MUX2_X1 U6309 ( .A(_01902__PTR33), .B(_01982__PTR1), .S(P1_StateBS16), .Z(_01902__PTR17) );
  MUX2_X1 U6310 ( .A(_01902__PTR34), .B(_01982__PTR2), .S(P1_StateBS16), .Z(_01902__PTR18) );
  MUX2_X1 U6311 ( .A(_01902__PTR35), .B(_01982__PTR3), .S(P1_StateBS16), .Z(_01902__PTR19) );
  MUX2_X1 U6312 ( .A(_01902__PTR36), .B(_01982__PTR4), .S(P1_StateBS16), .Z(_01902__PTR20) );
  MUX2_X1 U6313 ( .A(_01902__PTR37), .B(_01982__PTR5), .S(P1_StateBS16), .Z(_01902__PTR21) );
  MUX2_X1 U6314 ( .A(_01902__PTR38), .B(_01982__PTR6), .S(P1_StateBS16), .Z(_01902__PTR22) );
  MUX2_X1 U6315 ( .A(_01902__PTR39), .B(_01982__PTR7), .S(P1_StateBS16), .Z(_01902__PTR23) );
  MUX2_X1 U6316 ( .A(_01900__PTR32), .B(_01981__PTR0), .S(P1_StateBS16), .Z(_01900__PTR16) );
  MUX2_X1 U6317 ( .A(_01900__PTR33), .B(_01981__PTR1), .S(P1_StateBS16), .Z(_01900__PTR17) );
  MUX2_X1 U6318 ( .A(_01900__PTR34), .B(_01981__PTR2), .S(P1_StateBS16), .Z(_01900__PTR18) );
  MUX2_X1 U6319 ( .A(_01900__PTR35), .B(_01981__PTR3), .S(P1_StateBS16), .Z(_01900__PTR19) );
  MUX2_X1 U6320 ( .A(_01900__PTR36), .B(_01981__PTR4), .S(P1_StateBS16), .Z(_01900__PTR20) );
  MUX2_X1 U6321 ( .A(_01900__PTR37), .B(_01981__PTR5), .S(P1_StateBS16), .Z(_01900__PTR21) );
  MUX2_X1 U6322 ( .A(_01900__PTR38), .B(_01981__PTR6), .S(P1_StateBS16), .Z(_01900__PTR22) );
  MUX2_X1 U6323 ( .A(_01900__PTR39), .B(_01981__PTR7), .S(P1_StateBS16), .Z(_01900__PTR23) );
  MUX2_X1 U6324 ( .A(_01898__PTR32), .B(_01980__PTR0), .S(P1_StateBS16), .Z(_01898__PTR16) );
  MUX2_X1 U6325 ( .A(_01898__PTR33), .B(_01980__PTR1), .S(P1_StateBS16), .Z(_01898__PTR17) );
  MUX2_X1 U6326 ( .A(_01898__PTR34), .B(_01980__PTR2), .S(P1_StateBS16), .Z(_01898__PTR18) );
  MUX2_X1 U6327 ( .A(_01898__PTR35), .B(_01980__PTR3), .S(P1_StateBS16), .Z(_01898__PTR19) );
  MUX2_X1 U6328 ( .A(_01898__PTR36), .B(_01980__PTR4), .S(P1_StateBS16), .Z(_01898__PTR20) );
  MUX2_X1 U6329 ( .A(_01898__PTR37), .B(_01980__PTR5), .S(P1_StateBS16), .Z(_01898__PTR21) );
  MUX2_X1 U6330 ( .A(_01898__PTR38), .B(_01980__PTR6), .S(P1_StateBS16), .Z(_01898__PTR22) );
  MUX2_X1 U6331 ( .A(_01898__PTR39), .B(_01980__PTR7), .S(P1_StateBS16), .Z(_01898__PTR23) );
  MUX2_X1 U6332 ( .A(_02946__PTR1), .B(_01892__PTR129), .S(_02714__PTR31), .Z(_01996__PTR1) );
  MUX2_X1 U6333 ( .A(_02946__PTR2), .B(_01892__PTR130), .S(_02714__PTR31), .Z(_01996__PTR2) );
  MUX2_X1 U6334 ( .A(_02946__PTR3), .B(_01892__PTR131), .S(_02714__PTR31), .Z(_01996__PTR3) );
  MUX2_X1 U6335 ( .A(_02946__PTR4), .B(_01892__PTR132), .S(_02714__PTR31), .Z(_01996__PTR4) );
  MUX2_X1 U6336 ( .A(_02946__PTR5), .B(_01892__PTR133), .S(_02714__PTR31), .Z(_01996__PTR5) );
  MUX2_X1 U6337 ( .A(_02946__PTR6), .B(_01892__PTR134), .S(_02714__PTR31), .Z(_01996__PTR6) );
  MUX2_X1 U6338 ( .A(_02946__PTR7), .B(_01892__PTR135), .S(_02714__PTR31), .Z(_01996__PTR7) );
  MUX2_X1 U6339 ( .A(_02946__PTR8), .B(_01892__PTR136), .S(_02714__PTR31), .Z(_01996__PTR8) );
  MUX2_X1 U6340 ( .A(_02946__PTR9), .B(_01892__PTR137), .S(_02714__PTR31), .Z(_01996__PTR9) );
  MUX2_X1 U6341 ( .A(_02946__PTR10), .B(_01892__PTR138), .S(_02714__PTR31), .Z(_01996__PTR10) );
  MUX2_X1 U6342 ( .A(_02946__PTR11), .B(_01892__PTR139), .S(_02714__PTR31), .Z(_01996__PTR11) );
  MUX2_X1 U6343 ( .A(_02946__PTR12), .B(_01892__PTR140), .S(_02714__PTR31), .Z(_01996__PTR12) );
  MUX2_X1 U6344 ( .A(_02946__PTR13), .B(_01892__PTR141), .S(_02714__PTR31), .Z(_01996__PTR13) );
  MUX2_X1 U6345 ( .A(_02946__PTR14), .B(_01892__PTR142), .S(_02714__PTR31), .Z(_01996__PTR14) );
  MUX2_X1 U6346 ( .A(_02946__PTR15), .B(_01892__PTR143), .S(_02714__PTR31), .Z(_01996__PTR15) );
  MUX2_X1 U6347 ( .A(_02946__PTR16), .B(_01892__PTR144), .S(_02714__PTR31), .Z(_01996__PTR16) );
  MUX2_X1 U6348 ( .A(_02946__PTR17), .B(_01892__PTR145), .S(_02714__PTR31), .Z(_01996__PTR17) );
  MUX2_X1 U6349 ( .A(_02946__PTR18), .B(_01892__PTR146), .S(_02714__PTR31), .Z(_01996__PTR18) );
  MUX2_X1 U6350 ( .A(_02946__PTR19), .B(_01892__PTR147), .S(_02714__PTR31), .Z(_01996__PTR19) );
  MUX2_X1 U6351 ( .A(_02946__PTR20), .B(_01892__PTR148), .S(_02714__PTR31), .Z(_01996__PTR20) );
  MUX2_X1 U6352 ( .A(_02946__PTR21), .B(_01892__PTR149), .S(_02714__PTR31), .Z(_01996__PTR21) );
  MUX2_X1 U6353 ( .A(_02946__PTR22), .B(_01892__PTR150), .S(_02714__PTR31), .Z(_01996__PTR22) );
  MUX2_X1 U6354 ( .A(_02946__PTR23), .B(_01892__PTR151), .S(_02714__PTR31), .Z(_01996__PTR23) );
  MUX2_X1 U6355 ( .A(_02946__PTR24), .B(_01892__PTR152), .S(_02714__PTR31), .Z(_01996__PTR24) );
  MUX2_X1 U6356 ( .A(_02946__PTR25), .B(_01892__PTR153), .S(_02714__PTR31), .Z(_01996__PTR25) );
  MUX2_X1 U6357 ( .A(_02946__PTR26), .B(_01892__PTR154), .S(_02714__PTR31), .Z(_01996__PTR26) );
  MUX2_X1 U6358 ( .A(_02946__PTR27), .B(_01892__PTR155), .S(_02714__PTR31), .Z(_01996__PTR27) );
  MUX2_X1 U6359 ( .A(_02946__PTR28), .B(_01892__PTR156), .S(_02714__PTR31), .Z(_01996__PTR28) );
  MUX2_X1 U6360 ( .A(_02946__PTR29), .B(_01892__PTR157), .S(_02714__PTR31), .Z(_01996__PTR29) );
  MUX2_X1 U6361 ( .A(_02946__PTR30), .B(_01892__PTR158), .S(_02714__PTR31), .Z(_01996__PTR30) );
  MUX2_X1 U6362 ( .A(_02946__PTR31), .B(_01892__PTR159), .S(_02714__PTR31), .Z(_01996__PTR31) );
  MUX2_X1 U6363 ( .A(_01978__PTR0), .B(_02788__PTR0), .S(_01841__PTR0), .Z(_01995__PTR0) );
  MUX2_X1 U6364 ( .A(_01978__PTR1), .B(_02789__PTR1), .S(_01841__PTR0), .Z(_01995__PTR1) );
  MUX2_X1 U6365 ( .A(_01978__PTR2), .B(_02789__PTR2), .S(_01841__PTR0), .Z(_01995__PTR2) );
  MUX2_X1 U6366 ( .A(_01978__PTR3), .B(_02789__PTR3), .S(_01841__PTR0), .Z(_01995__PTR3) );
  MUX2_X1 U6367 ( .A(_01978__PTR4), .B(_02789__PTR4), .S(_01841__PTR0), .Z(_01995__PTR4) );
  MUX2_X1 U6368 ( .A(_01978__PTR5), .B(_02789__PTR5), .S(_01841__PTR0), .Z(_01995__PTR5) );
  MUX2_X1 U6369 ( .A(_01978__PTR6), .B(_02789__PTR6), .S(_01841__PTR0), .Z(_01995__PTR6) );
  MUX2_X1 U6370 ( .A(_01978__PTR7), .B(_02789__PTR7), .S(_01841__PTR0), .Z(_01995__PTR7) );
  MUX2_X1 U6371 ( .A(_01977__PTR0), .B(_02788__PTR0), .S(_01841__PTR1), .Z(_01994__PTR0) );
  MUX2_X1 U6372 ( .A(_01977__PTR1), .B(_02789__PTR1), .S(_01841__PTR1), .Z(_01994__PTR1) );
  MUX2_X1 U6373 ( .A(_01977__PTR2), .B(_02789__PTR2), .S(_01841__PTR1), .Z(_01994__PTR2) );
  MUX2_X1 U6374 ( .A(_01977__PTR3), .B(_02789__PTR3), .S(_01841__PTR1), .Z(_01994__PTR3) );
  MUX2_X1 U6375 ( .A(_01977__PTR4), .B(_02789__PTR4), .S(_01841__PTR1), .Z(_01994__PTR4) );
  MUX2_X1 U6376 ( .A(_01977__PTR5), .B(_02789__PTR5), .S(_01841__PTR1), .Z(_01994__PTR5) );
  MUX2_X1 U6377 ( .A(_01977__PTR6), .B(_02789__PTR6), .S(_01841__PTR1), .Z(_01994__PTR6) );
  MUX2_X1 U6378 ( .A(_01977__PTR7), .B(_02789__PTR7), .S(_01841__PTR1), .Z(_01994__PTR7) );
  MUX2_X1 U6379 ( .A(_01976__PTR0), .B(_02788__PTR0), .S(_01841__PTR2), .Z(_01993__PTR0) );
  MUX2_X1 U6380 ( .A(_01976__PTR1), .B(_02789__PTR1), .S(_01841__PTR2), .Z(_01993__PTR1) );
  MUX2_X1 U6381 ( .A(_01976__PTR2), .B(_02789__PTR2), .S(_01841__PTR2), .Z(_01993__PTR2) );
  MUX2_X1 U6382 ( .A(_01976__PTR3), .B(_02789__PTR3), .S(_01841__PTR2), .Z(_01993__PTR3) );
  MUX2_X1 U6383 ( .A(_01976__PTR4), .B(_02789__PTR4), .S(_01841__PTR2), .Z(_01993__PTR4) );
  MUX2_X1 U6384 ( .A(_01976__PTR5), .B(_02789__PTR5), .S(_01841__PTR2), .Z(_01993__PTR5) );
  MUX2_X1 U6385 ( .A(_01976__PTR6), .B(_02789__PTR6), .S(_01841__PTR2), .Z(_01993__PTR6) );
  MUX2_X1 U6386 ( .A(_01976__PTR7), .B(_02789__PTR7), .S(_01841__PTR2), .Z(_01993__PTR7) );
  MUX2_X1 U6387 ( .A(_01975__PTR0), .B(_02788__PTR0), .S(_01841__PTR3), .Z(_01992__PTR0) );
  MUX2_X1 U6388 ( .A(_01975__PTR1), .B(_02789__PTR1), .S(_01841__PTR3), .Z(_01992__PTR1) );
  MUX2_X1 U6389 ( .A(_01975__PTR2), .B(_02789__PTR2), .S(_01841__PTR3), .Z(_01992__PTR2) );
  MUX2_X1 U6390 ( .A(_01975__PTR3), .B(_02789__PTR3), .S(_01841__PTR3), .Z(_01992__PTR3) );
  MUX2_X1 U6391 ( .A(_01975__PTR4), .B(_02789__PTR4), .S(_01841__PTR3), .Z(_01992__PTR4) );
  MUX2_X1 U6392 ( .A(_01975__PTR5), .B(_02789__PTR5), .S(_01841__PTR3), .Z(_01992__PTR5) );
  MUX2_X1 U6393 ( .A(_01975__PTR6), .B(_02789__PTR6), .S(_01841__PTR3), .Z(_01992__PTR6) );
  MUX2_X1 U6394 ( .A(_01975__PTR7), .B(_02789__PTR7), .S(_01841__PTR3), .Z(_01992__PTR7) );
  MUX2_X1 U6395 ( .A(_01974__PTR0), .B(_02788__PTR0), .S(_01841__PTR4), .Z(_01991__PTR0) );
  MUX2_X1 U6396 ( .A(_01974__PTR1), .B(_02789__PTR1), .S(_01841__PTR4), .Z(_01991__PTR1) );
  MUX2_X1 U6397 ( .A(_01974__PTR2), .B(_02789__PTR2), .S(_01841__PTR4), .Z(_01991__PTR2) );
  MUX2_X1 U6398 ( .A(_01974__PTR3), .B(_02789__PTR3), .S(_01841__PTR4), .Z(_01991__PTR3) );
  MUX2_X1 U6399 ( .A(_01974__PTR4), .B(_02789__PTR4), .S(_01841__PTR4), .Z(_01991__PTR4) );
  MUX2_X1 U6400 ( .A(_01974__PTR5), .B(_02789__PTR5), .S(_01841__PTR4), .Z(_01991__PTR5) );
  MUX2_X1 U6401 ( .A(_01974__PTR6), .B(_02789__PTR6), .S(_01841__PTR4), .Z(_01991__PTR6) );
  MUX2_X1 U6402 ( .A(_01974__PTR7), .B(_02789__PTR7), .S(_01841__PTR4), .Z(_01991__PTR7) );
  MUX2_X1 U6403 ( .A(_01973__PTR0), .B(_02788__PTR0), .S(_01841__PTR5), .Z(_01990__PTR0) );
  MUX2_X1 U6404 ( .A(_01973__PTR1), .B(_02789__PTR1), .S(_01841__PTR5), .Z(_01990__PTR1) );
  MUX2_X1 U6405 ( .A(_01973__PTR2), .B(_02789__PTR2), .S(_01841__PTR5), .Z(_01990__PTR2) );
  MUX2_X1 U6406 ( .A(_01973__PTR3), .B(_02789__PTR3), .S(_01841__PTR5), .Z(_01990__PTR3) );
  MUX2_X1 U6407 ( .A(_01973__PTR4), .B(_02789__PTR4), .S(_01841__PTR5), .Z(_01990__PTR4) );
  MUX2_X1 U6408 ( .A(_01973__PTR5), .B(_02789__PTR5), .S(_01841__PTR5), .Z(_01990__PTR5) );
  MUX2_X1 U6409 ( .A(_01973__PTR6), .B(_02789__PTR6), .S(_01841__PTR5), .Z(_01990__PTR6) );
  MUX2_X1 U6410 ( .A(_01973__PTR7), .B(_02789__PTR7), .S(_01841__PTR5), .Z(_01990__PTR7) );
  MUX2_X1 U6411 ( .A(_01972__PTR0), .B(_02788__PTR0), .S(_01841__PTR6), .Z(_01989__PTR0) );
  MUX2_X1 U6412 ( .A(_01972__PTR1), .B(_02789__PTR1), .S(_01841__PTR6), .Z(_01989__PTR1) );
  MUX2_X1 U6413 ( .A(_01972__PTR2), .B(_02789__PTR2), .S(_01841__PTR6), .Z(_01989__PTR2) );
  MUX2_X1 U6414 ( .A(_01972__PTR3), .B(_02789__PTR3), .S(_01841__PTR6), .Z(_01989__PTR3) );
  MUX2_X1 U6415 ( .A(_01972__PTR4), .B(_02789__PTR4), .S(_01841__PTR6), .Z(_01989__PTR4) );
  MUX2_X1 U6416 ( .A(_01972__PTR5), .B(_02789__PTR5), .S(_01841__PTR6), .Z(_01989__PTR5) );
  MUX2_X1 U6417 ( .A(_01972__PTR6), .B(_02789__PTR6), .S(_01841__PTR6), .Z(_01989__PTR6) );
  MUX2_X1 U6418 ( .A(_01972__PTR7), .B(_02789__PTR7), .S(_01841__PTR6), .Z(_01989__PTR7) );
  MUX2_X1 U6419 ( .A(_01971__PTR0), .B(_02788__PTR0), .S(_01841__PTR7), .Z(_01988__PTR0) );
  MUX2_X1 U6420 ( .A(_01971__PTR1), .B(_02789__PTR1), .S(_01841__PTR7), .Z(_01988__PTR1) );
  MUX2_X1 U6421 ( .A(_01971__PTR2), .B(_02789__PTR2), .S(_01841__PTR7), .Z(_01988__PTR2) );
  MUX2_X1 U6422 ( .A(_01971__PTR3), .B(_02789__PTR3), .S(_01841__PTR7), .Z(_01988__PTR3) );
  MUX2_X1 U6423 ( .A(_01971__PTR4), .B(_02789__PTR4), .S(_01841__PTR7), .Z(_01988__PTR4) );
  MUX2_X1 U6424 ( .A(_01971__PTR5), .B(_02789__PTR5), .S(_01841__PTR7), .Z(_01988__PTR5) );
  MUX2_X1 U6425 ( .A(_01971__PTR6), .B(_02789__PTR6), .S(_01841__PTR7), .Z(_01988__PTR6) );
  MUX2_X1 U6426 ( .A(_01971__PTR7), .B(_02789__PTR7), .S(_01841__PTR7), .Z(_01988__PTR7) );
  MUX2_X1 U6427 ( .A(_01970__PTR0), .B(_02788__PTR0), .S(_01841__PTR8), .Z(_01987__PTR0) );
  MUX2_X1 U6428 ( .A(_01970__PTR1), .B(_02789__PTR1), .S(_01841__PTR8), .Z(_01987__PTR1) );
  MUX2_X1 U6429 ( .A(_01970__PTR2), .B(_02789__PTR2), .S(_01841__PTR8), .Z(_01987__PTR2) );
  MUX2_X1 U6430 ( .A(_01970__PTR3), .B(_02789__PTR3), .S(_01841__PTR8), .Z(_01987__PTR3) );
  MUX2_X1 U6431 ( .A(_01970__PTR4), .B(_02789__PTR4), .S(_01841__PTR8), .Z(_01987__PTR4) );
  MUX2_X1 U6432 ( .A(_01970__PTR5), .B(_02789__PTR5), .S(_01841__PTR8), .Z(_01987__PTR5) );
  MUX2_X1 U6433 ( .A(_01970__PTR6), .B(_02789__PTR6), .S(_01841__PTR8), .Z(_01987__PTR6) );
  MUX2_X1 U6434 ( .A(_01970__PTR7), .B(_02789__PTR7), .S(_01841__PTR8), .Z(_01987__PTR7) );
  MUX2_X1 U6435 ( .A(_01969__PTR0), .B(_02788__PTR0), .S(_01841__PTR9), .Z(_01986__PTR0) );
  MUX2_X1 U6436 ( .A(_01969__PTR1), .B(_02789__PTR1), .S(_01841__PTR9), .Z(_01986__PTR1) );
  MUX2_X1 U6437 ( .A(_01969__PTR2), .B(_02789__PTR2), .S(_01841__PTR9), .Z(_01986__PTR2) );
  MUX2_X1 U6438 ( .A(_01969__PTR3), .B(_02789__PTR3), .S(_01841__PTR9), .Z(_01986__PTR3) );
  MUX2_X1 U6439 ( .A(_01969__PTR4), .B(_02789__PTR4), .S(_01841__PTR9), .Z(_01986__PTR4) );
  MUX2_X1 U6440 ( .A(_01969__PTR5), .B(_02789__PTR5), .S(_01841__PTR9), .Z(_01986__PTR5) );
  MUX2_X1 U6441 ( .A(_01969__PTR6), .B(_02789__PTR6), .S(_01841__PTR9), .Z(_01986__PTR6) );
  MUX2_X1 U6442 ( .A(_01969__PTR7), .B(_02789__PTR7), .S(_01841__PTR9), .Z(_01986__PTR7) );
  MUX2_X1 U6443 ( .A(_01968__PTR0), .B(_02788__PTR0), .S(_01841__PTR10), .Z(_01985__PTR0) );
  MUX2_X1 U6444 ( .A(_01968__PTR1), .B(_02789__PTR1), .S(_01841__PTR10), .Z(_01985__PTR1) );
  MUX2_X1 U6445 ( .A(_01968__PTR2), .B(_02789__PTR2), .S(_01841__PTR10), .Z(_01985__PTR2) );
  MUX2_X1 U6446 ( .A(_01968__PTR3), .B(_02789__PTR3), .S(_01841__PTR10), .Z(_01985__PTR3) );
  MUX2_X1 U6447 ( .A(_01968__PTR4), .B(_02789__PTR4), .S(_01841__PTR10), .Z(_01985__PTR4) );
  MUX2_X1 U6448 ( .A(_01968__PTR5), .B(_02789__PTR5), .S(_01841__PTR10), .Z(_01985__PTR5) );
  MUX2_X1 U6449 ( .A(_01968__PTR6), .B(_02789__PTR6), .S(_01841__PTR10), .Z(_01985__PTR6) );
  MUX2_X1 U6450 ( .A(_01968__PTR7), .B(_02789__PTR7), .S(_01841__PTR10), .Z(_01985__PTR7) );
  MUX2_X1 U6451 ( .A(_01967__PTR0), .B(_02788__PTR0), .S(_01841__PTR11), .Z(_01984__PTR0) );
  MUX2_X1 U6452 ( .A(_01967__PTR1), .B(_02789__PTR1), .S(_01841__PTR11), .Z(_01984__PTR1) );
  MUX2_X1 U6453 ( .A(_01967__PTR2), .B(_02789__PTR2), .S(_01841__PTR11), .Z(_01984__PTR2) );
  MUX2_X1 U6454 ( .A(_01967__PTR3), .B(_02789__PTR3), .S(_01841__PTR11), .Z(_01984__PTR3) );
  MUX2_X1 U6455 ( .A(_01967__PTR4), .B(_02789__PTR4), .S(_01841__PTR11), .Z(_01984__PTR4) );
  MUX2_X1 U6456 ( .A(_01967__PTR5), .B(_02789__PTR5), .S(_01841__PTR11), .Z(_01984__PTR5) );
  MUX2_X1 U6457 ( .A(_01967__PTR6), .B(_02789__PTR6), .S(_01841__PTR11), .Z(_01984__PTR6) );
  MUX2_X1 U6458 ( .A(_01967__PTR7), .B(_02789__PTR7), .S(_01841__PTR11), .Z(_01984__PTR7) );
  MUX2_X1 U6459 ( .A(_01966__PTR0), .B(_02788__PTR0), .S(_01841__PTR12), .Z(_01983__PTR0) );
  MUX2_X1 U6460 ( .A(_01966__PTR1), .B(_02789__PTR1), .S(_01841__PTR12), .Z(_01983__PTR1) );
  MUX2_X1 U6461 ( .A(_01966__PTR2), .B(_02789__PTR2), .S(_01841__PTR12), .Z(_01983__PTR2) );
  MUX2_X1 U6462 ( .A(_01966__PTR3), .B(_02789__PTR3), .S(_01841__PTR12), .Z(_01983__PTR3) );
  MUX2_X1 U6463 ( .A(_01966__PTR4), .B(_02789__PTR4), .S(_01841__PTR12), .Z(_01983__PTR4) );
  MUX2_X1 U6464 ( .A(_01966__PTR5), .B(_02789__PTR5), .S(_01841__PTR12), .Z(_01983__PTR5) );
  MUX2_X1 U6465 ( .A(_01966__PTR6), .B(_02789__PTR6), .S(_01841__PTR12), .Z(_01983__PTR6) );
  MUX2_X1 U6466 ( .A(_01966__PTR7), .B(_02789__PTR7), .S(_01841__PTR12), .Z(_01983__PTR7) );
  MUX2_X1 U6467 ( .A(_01965__PTR0), .B(_02788__PTR0), .S(_01841__PTR13), .Z(_01982__PTR0) );
  MUX2_X1 U6468 ( .A(_01965__PTR1), .B(_02789__PTR1), .S(_01841__PTR13), .Z(_01982__PTR1) );
  MUX2_X1 U6469 ( .A(_01965__PTR2), .B(_02789__PTR2), .S(_01841__PTR13), .Z(_01982__PTR2) );
  MUX2_X1 U6470 ( .A(_01965__PTR3), .B(_02789__PTR3), .S(_01841__PTR13), .Z(_01982__PTR3) );
  MUX2_X1 U6471 ( .A(_01965__PTR4), .B(_02789__PTR4), .S(_01841__PTR13), .Z(_01982__PTR4) );
  MUX2_X1 U6472 ( .A(_01965__PTR5), .B(_02789__PTR5), .S(_01841__PTR13), .Z(_01982__PTR5) );
  MUX2_X1 U6473 ( .A(_01965__PTR6), .B(_02789__PTR6), .S(_01841__PTR13), .Z(_01982__PTR6) );
  MUX2_X1 U6474 ( .A(_01965__PTR7), .B(_02789__PTR7), .S(_01841__PTR13), .Z(_01982__PTR7) );
  MUX2_X1 U6475 ( .A(_01964__PTR0), .B(_02788__PTR0), .S(_01841__PTR14), .Z(_01981__PTR0) );
  MUX2_X1 U6476 ( .A(_01964__PTR1), .B(_02789__PTR1), .S(_01841__PTR14), .Z(_01981__PTR1) );
  MUX2_X1 U6477 ( .A(_01964__PTR2), .B(_02789__PTR2), .S(_01841__PTR14), .Z(_01981__PTR2) );
  MUX2_X1 U6478 ( .A(_01964__PTR3), .B(_02789__PTR3), .S(_01841__PTR14), .Z(_01981__PTR3) );
  MUX2_X1 U6479 ( .A(_01964__PTR4), .B(_02789__PTR4), .S(_01841__PTR14), .Z(_01981__PTR4) );
  MUX2_X1 U6480 ( .A(_01964__PTR5), .B(_02789__PTR5), .S(_01841__PTR14), .Z(_01981__PTR5) );
  MUX2_X1 U6481 ( .A(_01964__PTR6), .B(_02789__PTR6), .S(_01841__PTR14), .Z(_01981__PTR6) );
  MUX2_X1 U6482 ( .A(_01964__PTR7), .B(_02789__PTR7), .S(_01841__PTR14), .Z(_01981__PTR7) );
  MUX2_X1 U6483 ( .A(_01963__PTR0), .B(_02788__PTR0), .S(_01841__PTR15), .Z(_01980__PTR0) );
  MUX2_X1 U6484 ( .A(_01963__PTR1), .B(_02789__PTR1), .S(_01841__PTR15), .Z(_01980__PTR1) );
  MUX2_X1 U6485 ( .A(_01963__PTR2), .B(_02789__PTR2), .S(_01841__PTR15), .Z(_01980__PTR2) );
  MUX2_X1 U6486 ( .A(_01963__PTR3), .B(_02789__PTR3), .S(_01841__PTR15), .Z(_01980__PTR3) );
  MUX2_X1 U6487 ( .A(_01963__PTR4), .B(_02789__PTR4), .S(_01841__PTR15), .Z(_01980__PTR4) );
  MUX2_X1 U6488 ( .A(_01963__PTR5), .B(_02789__PTR5), .S(_01841__PTR15), .Z(_01980__PTR5) );
  MUX2_X1 U6489 ( .A(_01963__PTR6), .B(_02789__PTR6), .S(_01841__PTR15), .Z(_01980__PTR6) );
  MUX2_X1 U6490 ( .A(_01963__PTR7), .B(_02789__PTR7), .S(_01841__PTR15), .Z(_01980__PTR7) );
  MUX2_X1 U6491 ( .A(_01928__PTR32), .B(_02783__PTR0), .S(_01839__PTR0), .Z(_01978__PTR0) );
  MUX2_X1 U6492 ( .A(_01928__PTR33), .B(_02784__PTR1), .S(_01839__PTR0), .Z(_01978__PTR1) );
  MUX2_X1 U6493 ( .A(_01928__PTR34), .B(_02784__PTR2), .S(_01839__PTR0), .Z(_01978__PTR2) );
  MUX2_X1 U6494 ( .A(_01928__PTR35), .B(_02784__PTR3), .S(_01839__PTR0), .Z(_01978__PTR3) );
  MUX2_X1 U6495 ( .A(_01928__PTR36), .B(_02784__PTR4), .S(_01839__PTR0), .Z(_01978__PTR4) );
  MUX2_X1 U6496 ( .A(_01928__PTR37), .B(_02784__PTR5), .S(_01839__PTR0), .Z(_01978__PTR5) );
  MUX2_X1 U6497 ( .A(_01928__PTR38), .B(_02784__PTR6), .S(_01839__PTR0), .Z(_01978__PTR6) );
  MUX2_X1 U6498 ( .A(_01928__PTR39), .B(_02784__PTR7), .S(_01839__PTR0), .Z(_01978__PTR7) );
  MUX2_X1 U6499 ( .A(_01926__PTR32), .B(_02783__PTR0), .S(_01839__PTR1), .Z(_01977__PTR0) );
  MUX2_X1 U6500 ( .A(_01926__PTR33), .B(_02784__PTR1), .S(_01839__PTR1), .Z(_01977__PTR1) );
  MUX2_X1 U6501 ( .A(_01926__PTR34), .B(_02784__PTR2), .S(_01839__PTR1), .Z(_01977__PTR2) );
  MUX2_X1 U6502 ( .A(_01926__PTR35), .B(_02784__PTR3), .S(_01839__PTR1), .Z(_01977__PTR3) );
  MUX2_X1 U6503 ( .A(_01926__PTR36), .B(_02784__PTR4), .S(_01839__PTR1), .Z(_01977__PTR4) );
  MUX2_X1 U6504 ( .A(_01926__PTR37), .B(_02784__PTR5), .S(_01839__PTR1), .Z(_01977__PTR5) );
  MUX2_X1 U6505 ( .A(_01926__PTR38), .B(_02784__PTR6), .S(_01839__PTR1), .Z(_01977__PTR6) );
  MUX2_X1 U6506 ( .A(_01926__PTR39), .B(_02784__PTR7), .S(_01839__PTR1), .Z(_01977__PTR7) );
  MUX2_X1 U6507 ( .A(_01924__PTR32), .B(_02783__PTR0), .S(_01839__PTR2), .Z(_01976__PTR0) );
  MUX2_X1 U6508 ( .A(_01924__PTR33), .B(_02784__PTR1), .S(_01839__PTR2), .Z(_01976__PTR1) );
  MUX2_X1 U6509 ( .A(_01924__PTR34), .B(_02784__PTR2), .S(_01839__PTR2), .Z(_01976__PTR2) );
  MUX2_X1 U6510 ( .A(_01924__PTR35), .B(_02784__PTR3), .S(_01839__PTR2), .Z(_01976__PTR3) );
  MUX2_X1 U6511 ( .A(_01924__PTR36), .B(_02784__PTR4), .S(_01839__PTR2), .Z(_01976__PTR4) );
  MUX2_X1 U6512 ( .A(_01924__PTR37), .B(_02784__PTR5), .S(_01839__PTR2), .Z(_01976__PTR5) );
  MUX2_X1 U6513 ( .A(_01924__PTR38), .B(_02784__PTR6), .S(_01839__PTR2), .Z(_01976__PTR6) );
  MUX2_X1 U6514 ( .A(_01924__PTR39), .B(_02784__PTR7), .S(_01839__PTR2), .Z(_01976__PTR7) );
  MUX2_X1 U6515 ( .A(_01922__PTR32), .B(_02783__PTR0), .S(_01839__PTR3), .Z(_01975__PTR0) );
  MUX2_X1 U6516 ( .A(_01922__PTR33), .B(_02784__PTR1), .S(_01839__PTR3), .Z(_01975__PTR1) );
  MUX2_X1 U6517 ( .A(_01922__PTR34), .B(_02784__PTR2), .S(_01839__PTR3), .Z(_01975__PTR2) );
  MUX2_X1 U6518 ( .A(_01922__PTR35), .B(_02784__PTR3), .S(_01839__PTR3), .Z(_01975__PTR3) );
  MUX2_X1 U6519 ( .A(_01922__PTR36), .B(_02784__PTR4), .S(_01839__PTR3), .Z(_01975__PTR4) );
  MUX2_X1 U6520 ( .A(_01922__PTR37), .B(_02784__PTR5), .S(_01839__PTR3), .Z(_01975__PTR5) );
  MUX2_X1 U6521 ( .A(_01922__PTR38), .B(_02784__PTR6), .S(_01839__PTR3), .Z(_01975__PTR6) );
  MUX2_X1 U6522 ( .A(_01922__PTR39), .B(_02784__PTR7), .S(_01839__PTR3), .Z(_01975__PTR7) );
  MUX2_X1 U6523 ( .A(_01920__PTR32), .B(_02783__PTR0), .S(_01839__PTR4), .Z(_01974__PTR0) );
  MUX2_X1 U6524 ( .A(_01920__PTR33), .B(_02784__PTR1), .S(_01839__PTR4), .Z(_01974__PTR1) );
  MUX2_X1 U6525 ( .A(_01920__PTR34), .B(_02784__PTR2), .S(_01839__PTR4), .Z(_01974__PTR2) );
  MUX2_X1 U6526 ( .A(_01920__PTR35), .B(_02784__PTR3), .S(_01839__PTR4), .Z(_01974__PTR3) );
  MUX2_X1 U6527 ( .A(_01920__PTR36), .B(_02784__PTR4), .S(_01839__PTR4), .Z(_01974__PTR4) );
  MUX2_X1 U6528 ( .A(_01920__PTR37), .B(_02784__PTR5), .S(_01839__PTR4), .Z(_01974__PTR5) );
  MUX2_X1 U6529 ( .A(_01920__PTR38), .B(_02784__PTR6), .S(_01839__PTR4), .Z(_01974__PTR6) );
  MUX2_X1 U6530 ( .A(_01920__PTR39), .B(_02784__PTR7), .S(_01839__PTR4), .Z(_01974__PTR7) );
  MUX2_X1 U6531 ( .A(_01918__PTR32), .B(_02783__PTR0), .S(_01839__PTR5), .Z(_01973__PTR0) );
  MUX2_X1 U6532 ( .A(_01918__PTR33), .B(_02784__PTR1), .S(_01839__PTR5), .Z(_01973__PTR1) );
  MUX2_X1 U6533 ( .A(_01918__PTR34), .B(_02784__PTR2), .S(_01839__PTR5), .Z(_01973__PTR2) );
  MUX2_X1 U6534 ( .A(_01918__PTR35), .B(_02784__PTR3), .S(_01839__PTR5), .Z(_01973__PTR3) );
  MUX2_X1 U6535 ( .A(_01918__PTR36), .B(_02784__PTR4), .S(_01839__PTR5), .Z(_01973__PTR4) );
  MUX2_X1 U6536 ( .A(_01918__PTR37), .B(_02784__PTR5), .S(_01839__PTR5), .Z(_01973__PTR5) );
  MUX2_X1 U6537 ( .A(_01918__PTR38), .B(_02784__PTR6), .S(_01839__PTR5), .Z(_01973__PTR6) );
  MUX2_X1 U6538 ( .A(_01918__PTR39), .B(_02784__PTR7), .S(_01839__PTR5), .Z(_01973__PTR7) );
  MUX2_X1 U6539 ( .A(_01916__PTR32), .B(_02783__PTR0), .S(_01839__PTR6), .Z(_01972__PTR0) );
  MUX2_X1 U6540 ( .A(_01916__PTR33), .B(_02784__PTR1), .S(_01839__PTR6), .Z(_01972__PTR1) );
  MUX2_X1 U6541 ( .A(_01916__PTR34), .B(_02784__PTR2), .S(_01839__PTR6), .Z(_01972__PTR2) );
  MUX2_X1 U6542 ( .A(_01916__PTR35), .B(_02784__PTR3), .S(_01839__PTR6), .Z(_01972__PTR3) );
  MUX2_X1 U6543 ( .A(_01916__PTR36), .B(_02784__PTR4), .S(_01839__PTR6), .Z(_01972__PTR4) );
  MUX2_X1 U6544 ( .A(_01916__PTR37), .B(_02784__PTR5), .S(_01839__PTR6), .Z(_01972__PTR5) );
  MUX2_X1 U6545 ( .A(_01916__PTR38), .B(_02784__PTR6), .S(_01839__PTR6), .Z(_01972__PTR6) );
  MUX2_X1 U6546 ( .A(_01916__PTR39), .B(_02784__PTR7), .S(_01839__PTR6), .Z(_01972__PTR7) );
  MUX2_X1 U6547 ( .A(_01914__PTR32), .B(_02783__PTR0), .S(_01839__PTR7), .Z(_01971__PTR0) );
  MUX2_X1 U6548 ( .A(_01914__PTR33), .B(_02784__PTR1), .S(_01839__PTR7), .Z(_01971__PTR1) );
  MUX2_X1 U6549 ( .A(_01914__PTR34), .B(_02784__PTR2), .S(_01839__PTR7), .Z(_01971__PTR2) );
  MUX2_X1 U6550 ( .A(_01914__PTR35), .B(_02784__PTR3), .S(_01839__PTR7), .Z(_01971__PTR3) );
  MUX2_X1 U6551 ( .A(_01914__PTR36), .B(_02784__PTR4), .S(_01839__PTR7), .Z(_01971__PTR4) );
  MUX2_X1 U6552 ( .A(_01914__PTR37), .B(_02784__PTR5), .S(_01839__PTR7), .Z(_01971__PTR5) );
  MUX2_X1 U6553 ( .A(_01914__PTR38), .B(_02784__PTR6), .S(_01839__PTR7), .Z(_01971__PTR6) );
  MUX2_X1 U6554 ( .A(_01914__PTR39), .B(_02784__PTR7), .S(_01839__PTR7), .Z(_01971__PTR7) );
  MUX2_X1 U6555 ( .A(_01912__PTR32), .B(_02783__PTR0), .S(_01839__PTR8), .Z(_01970__PTR0) );
  MUX2_X1 U6556 ( .A(_01912__PTR33), .B(_02784__PTR1), .S(_01839__PTR8), .Z(_01970__PTR1) );
  MUX2_X1 U6557 ( .A(_01912__PTR34), .B(_02784__PTR2), .S(_01839__PTR8), .Z(_01970__PTR2) );
  MUX2_X1 U6558 ( .A(_01912__PTR35), .B(_02784__PTR3), .S(_01839__PTR8), .Z(_01970__PTR3) );
  MUX2_X1 U6559 ( .A(_01912__PTR36), .B(_02784__PTR4), .S(_01839__PTR8), .Z(_01970__PTR4) );
  MUX2_X1 U6560 ( .A(_01912__PTR37), .B(_02784__PTR5), .S(_01839__PTR8), .Z(_01970__PTR5) );
  MUX2_X1 U6561 ( .A(_01912__PTR38), .B(_02784__PTR6), .S(_01839__PTR8), .Z(_01970__PTR6) );
  MUX2_X1 U6562 ( .A(_01912__PTR39), .B(_02784__PTR7), .S(_01839__PTR8), .Z(_01970__PTR7) );
  MUX2_X1 U6563 ( .A(_01910__PTR32), .B(_02783__PTR0), .S(_01839__PTR9), .Z(_01969__PTR0) );
  MUX2_X1 U6564 ( .A(_01910__PTR33), .B(_02784__PTR1), .S(_01839__PTR9), .Z(_01969__PTR1) );
  MUX2_X1 U6565 ( .A(_01910__PTR34), .B(_02784__PTR2), .S(_01839__PTR9), .Z(_01969__PTR2) );
  MUX2_X1 U6566 ( .A(_01910__PTR35), .B(_02784__PTR3), .S(_01839__PTR9), .Z(_01969__PTR3) );
  MUX2_X1 U6567 ( .A(_01910__PTR36), .B(_02784__PTR4), .S(_01839__PTR9), .Z(_01969__PTR4) );
  MUX2_X1 U6568 ( .A(_01910__PTR37), .B(_02784__PTR5), .S(_01839__PTR9), .Z(_01969__PTR5) );
  MUX2_X1 U6569 ( .A(_01910__PTR38), .B(_02784__PTR6), .S(_01839__PTR9), .Z(_01969__PTR6) );
  MUX2_X1 U6570 ( .A(_01910__PTR39), .B(_02784__PTR7), .S(_01839__PTR9), .Z(_01969__PTR7) );
  MUX2_X1 U6571 ( .A(_01908__PTR32), .B(_02783__PTR0), .S(_01839__PTR10), .Z(_01968__PTR0) );
  MUX2_X1 U6572 ( .A(_01908__PTR33), .B(_02784__PTR1), .S(_01839__PTR10), .Z(_01968__PTR1) );
  MUX2_X1 U6573 ( .A(_01908__PTR34), .B(_02784__PTR2), .S(_01839__PTR10), .Z(_01968__PTR2) );
  MUX2_X1 U6574 ( .A(_01908__PTR35), .B(_02784__PTR3), .S(_01839__PTR10), .Z(_01968__PTR3) );
  MUX2_X1 U6575 ( .A(_01908__PTR36), .B(_02784__PTR4), .S(_01839__PTR10), .Z(_01968__PTR4) );
  MUX2_X1 U6576 ( .A(_01908__PTR37), .B(_02784__PTR5), .S(_01839__PTR10), .Z(_01968__PTR5) );
  MUX2_X1 U6577 ( .A(_01908__PTR38), .B(_02784__PTR6), .S(_01839__PTR10), .Z(_01968__PTR6) );
  MUX2_X1 U6578 ( .A(_01908__PTR39), .B(_02784__PTR7), .S(_01839__PTR10), .Z(_01968__PTR7) );
  MUX2_X1 U6579 ( .A(_01906__PTR32), .B(_02783__PTR0), .S(_01839__PTR11), .Z(_01967__PTR0) );
  MUX2_X1 U6580 ( .A(_01906__PTR33), .B(_02784__PTR1), .S(_01839__PTR11), .Z(_01967__PTR1) );
  MUX2_X1 U6581 ( .A(_01906__PTR34), .B(_02784__PTR2), .S(_01839__PTR11), .Z(_01967__PTR2) );
  MUX2_X1 U6582 ( .A(_01906__PTR35), .B(_02784__PTR3), .S(_01839__PTR11), .Z(_01967__PTR3) );
  MUX2_X1 U6583 ( .A(_01906__PTR36), .B(_02784__PTR4), .S(_01839__PTR11), .Z(_01967__PTR4) );
  MUX2_X1 U6584 ( .A(_01906__PTR37), .B(_02784__PTR5), .S(_01839__PTR11), .Z(_01967__PTR5) );
  MUX2_X1 U6585 ( .A(_01906__PTR38), .B(_02784__PTR6), .S(_01839__PTR11), .Z(_01967__PTR6) );
  MUX2_X1 U6586 ( .A(_01906__PTR39), .B(_02784__PTR7), .S(_01839__PTR11), .Z(_01967__PTR7) );
  MUX2_X1 U6587 ( .A(_01904__PTR32), .B(_02783__PTR0), .S(_01839__PTR12), .Z(_01966__PTR0) );
  MUX2_X1 U6588 ( .A(_01904__PTR33), .B(_02784__PTR1), .S(_01839__PTR12), .Z(_01966__PTR1) );
  MUX2_X1 U6589 ( .A(_01904__PTR34), .B(_02784__PTR2), .S(_01839__PTR12), .Z(_01966__PTR2) );
  MUX2_X1 U6590 ( .A(_01904__PTR35), .B(_02784__PTR3), .S(_01839__PTR12), .Z(_01966__PTR3) );
  MUX2_X1 U6591 ( .A(_01904__PTR36), .B(_02784__PTR4), .S(_01839__PTR12), .Z(_01966__PTR4) );
  MUX2_X1 U6592 ( .A(_01904__PTR37), .B(_02784__PTR5), .S(_01839__PTR12), .Z(_01966__PTR5) );
  MUX2_X1 U6593 ( .A(_01904__PTR38), .B(_02784__PTR6), .S(_01839__PTR12), .Z(_01966__PTR6) );
  MUX2_X1 U6594 ( .A(_01904__PTR39), .B(_02784__PTR7), .S(_01839__PTR12), .Z(_01966__PTR7) );
  MUX2_X1 U6595 ( .A(_01902__PTR32), .B(_02783__PTR0), .S(_01839__PTR13), .Z(_01965__PTR0) );
  MUX2_X1 U6596 ( .A(_01902__PTR33), .B(_02784__PTR1), .S(_01839__PTR13), .Z(_01965__PTR1) );
  MUX2_X1 U6597 ( .A(_01902__PTR34), .B(_02784__PTR2), .S(_01839__PTR13), .Z(_01965__PTR2) );
  MUX2_X1 U6598 ( .A(_01902__PTR35), .B(_02784__PTR3), .S(_01839__PTR13), .Z(_01965__PTR3) );
  MUX2_X1 U6599 ( .A(_01902__PTR36), .B(_02784__PTR4), .S(_01839__PTR13), .Z(_01965__PTR4) );
  MUX2_X1 U6600 ( .A(_01902__PTR37), .B(_02784__PTR5), .S(_01839__PTR13), .Z(_01965__PTR5) );
  MUX2_X1 U6601 ( .A(_01902__PTR38), .B(_02784__PTR6), .S(_01839__PTR13), .Z(_01965__PTR6) );
  MUX2_X1 U6602 ( .A(_01902__PTR39), .B(_02784__PTR7), .S(_01839__PTR13), .Z(_01965__PTR7) );
  MUX2_X1 U6603 ( .A(_01900__PTR32), .B(_02783__PTR0), .S(_01839__PTR14), .Z(_01964__PTR0) );
  MUX2_X1 U6604 ( .A(_01900__PTR33), .B(_02784__PTR1), .S(_01839__PTR14), .Z(_01964__PTR1) );
  MUX2_X1 U6605 ( .A(_01900__PTR34), .B(_02784__PTR2), .S(_01839__PTR14), .Z(_01964__PTR2) );
  MUX2_X1 U6606 ( .A(_01900__PTR35), .B(_02784__PTR3), .S(_01839__PTR14), .Z(_01964__PTR3) );
  MUX2_X1 U6607 ( .A(_01900__PTR36), .B(_02784__PTR4), .S(_01839__PTR14), .Z(_01964__PTR4) );
  MUX2_X1 U6608 ( .A(_01900__PTR37), .B(_02784__PTR5), .S(_01839__PTR14), .Z(_01964__PTR5) );
  MUX2_X1 U6609 ( .A(_01900__PTR38), .B(_02784__PTR6), .S(_01839__PTR14), .Z(_01964__PTR6) );
  MUX2_X1 U6610 ( .A(_01900__PTR39), .B(_02784__PTR7), .S(_01839__PTR14), .Z(_01964__PTR7) );
  MUX2_X1 U6611 ( .A(_01898__PTR32), .B(_02783__PTR0), .S(_01839__PTR15), .Z(_01963__PTR0) );
  MUX2_X1 U6612 ( .A(_01898__PTR33), .B(_02784__PTR1), .S(_01839__PTR15), .Z(_01963__PTR1) );
  MUX2_X1 U6613 ( .A(_01898__PTR34), .B(_02784__PTR2), .S(_01839__PTR15), .Z(_01963__PTR2) );
  MUX2_X1 U6614 ( .A(_01898__PTR35), .B(_02784__PTR3), .S(_01839__PTR15), .Z(_01963__PTR3) );
  MUX2_X1 U6615 ( .A(_01898__PTR36), .B(_02784__PTR4), .S(_01839__PTR15), .Z(_01963__PTR4) );
  MUX2_X1 U6616 ( .A(_01898__PTR37), .B(_02784__PTR5), .S(_01839__PTR15), .Z(_01963__PTR5) );
  MUX2_X1 U6617 ( .A(_01898__PTR38), .B(_02784__PTR6), .S(_01839__PTR15), .Z(_01963__PTR6) );
  MUX2_X1 U6618 ( .A(_01898__PTR39), .B(_02784__PTR7), .S(_01839__PTR15), .Z(_01963__PTR7) );
  MUX2_X1 U6619 ( .A(_01962__PTR0), .B(di1_PTR0), .S(_01837__PTR0), .Z(_01928__PTR32) );
  MUX2_X1 U6620 ( .A(_01962__PTR1), .B(di1_PTR1), .S(_01837__PTR0), .Z(_01928__PTR33) );
  MUX2_X1 U6621 ( .A(_01962__PTR2), .B(di1_PTR2), .S(_01837__PTR0), .Z(_01928__PTR34) );
  MUX2_X1 U6622 ( .A(_01962__PTR3), .B(di1_PTR3), .S(_01837__PTR0), .Z(_01928__PTR35) );
  MUX2_X1 U6623 ( .A(_01962__PTR4), .B(di1_PTR4), .S(_01837__PTR0), .Z(_01928__PTR36) );
  MUX2_X1 U6624 ( .A(_01962__PTR5), .B(di1_PTR5), .S(_01837__PTR0), .Z(_01928__PTR37) );
  MUX2_X1 U6625 ( .A(_01962__PTR6), .B(di1_PTR6), .S(_01837__PTR0), .Z(_01928__PTR38) );
  MUX2_X1 U6626 ( .A(_01962__PTR7), .B(di1_PTR7), .S(_01837__PTR0), .Z(_01928__PTR39) );
  MUX2_X1 U6627 ( .A(_01961__PTR0), .B(di1_PTR0), .S(_01837__PTR1), .Z(_01926__PTR32) );
  MUX2_X1 U6628 ( .A(_01961__PTR1), .B(di1_PTR1), .S(_01837__PTR1), .Z(_01926__PTR33) );
  MUX2_X1 U6629 ( .A(_01961__PTR2), .B(di1_PTR2), .S(_01837__PTR1), .Z(_01926__PTR34) );
  MUX2_X1 U6630 ( .A(_01961__PTR3), .B(di1_PTR3), .S(_01837__PTR1), .Z(_01926__PTR35) );
  MUX2_X1 U6631 ( .A(_01961__PTR4), .B(di1_PTR4), .S(_01837__PTR1), .Z(_01926__PTR36) );
  MUX2_X1 U6632 ( .A(_01961__PTR5), .B(di1_PTR5), .S(_01837__PTR1), .Z(_01926__PTR37) );
  MUX2_X1 U6633 ( .A(_01961__PTR6), .B(di1_PTR6), .S(_01837__PTR1), .Z(_01926__PTR38) );
  MUX2_X1 U6634 ( .A(_01961__PTR7), .B(di1_PTR7), .S(_01837__PTR1), .Z(_01926__PTR39) );
  MUX2_X1 U6635 ( .A(_01960__PTR0), .B(di1_PTR0), .S(_01837__PTR2), .Z(_01924__PTR32) );
  MUX2_X1 U6636 ( .A(_01960__PTR1), .B(di1_PTR1), .S(_01837__PTR2), .Z(_01924__PTR33) );
  MUX2_X1 U6637 ( .A(_01960__PTR2), .B(di1_PTR2), .S(_01837__PTR2), .Z(_01924__PTR34) );
  MUX2_X1 U6638 ( .A(_01960__PTR3), .B(di1_PTR3), .S(_01837__PTR2), .Z(_01924__PTR35) );
  MUX2_X1 U6639 ( .A(_01960__PTR4), .B(di1_PTR4), .S(_01837__PTR2), .Z(_01924__PTR36) );
  MUX2_X1 U6640 ( .A(_01960__PTR5), .B(di1_PTR5), .S(_01837__PTR2), .Z(_01924__PTR37) );
  MUX2_X1 U6641 ( .A(_01960__PTR6), .B(di1_PTR6), .S(_01837__PTR2), .Z(_01924__PTR38) );
  MUX2_X1 U6642 ( .A(_01960__PTR7), .B(di1_PTR7), .S(_01837__PTR2), .Z(_01924__PTR39) );
  MUX2_X1 U6643 ( .A(_01959__PTR0), .B(di1_PTR0), .S(_01837__PTR3), .Z(_01922__PTR32) );
  MUX2_X1 U6644 ( .A(_01959__PTR1), .B(di1_PTR1), .S(_01837__PTR3), .Z(_01922__PTR33) );
  MUX2_X1 U6645 ( .A(_01959__PTR2), .B(di1_PTR2), .S(_01837__PTR3), .Z(_01922__PTR34) );
  MUX2_X1 U6646 ( .A(_01959__PTR3), .B(di1_PTR3), .S(_01837__PTR3), .Z(_01922__PTR35) );
  MUX2_X1 U6647 ( .A(_01959__PTR4), .B(di1_PTR4), .S(_01837__PTR3), .Z(_01922__PTR36) );
  MUX2_X1 U6648 ( .A(_01959__PTR5), .B(di1_PTR5), .S(_01837__PTR3), .Z(_01922__PTR37) );
  MUX2_X1 U6649 ( .A(_01959__PTR6), .B(di1_PTR6), .S(_01837__PTR3), .Z(_01922__PTR38) );
  MUX2_X1 U6650 ( .A(_01959__PTR7), .B(di1_PTR7), .S(_01837__PTR3), .Z(_01922__PTR39) );
  MUX2_X1 U6651 ( .A(_01958__PTR0), .B(di1_PTR0), .S(_01837__PTR4), .Z(_01920__PTR32) );
  MUX2_X1 U6652 ( .A(_01958__PTR1), .B(di1_PTR1), .S(_01837__PTR4), .Z(_01920__PTR33) );
  MUX2_X1 U6653 ( .A(_01958__PTR2), .B(di1_PTR2), .S(_01837__PTR4), .Z(_01920__PTR34) );
  MUX2_X1 U6654 ( .A(_01958__PTR3), .B(di1_PTR3), .S(_01837__PTR4), .Z(_01920__PTR35) );
  MUX2_X1 U6655 ( .A(_01958__PTR4), .B(di1_PTR4), .S(_01837__PTR4), .Z(_01920__PTR36) );
  MUX2_X1 U6656 ( .A(_01958__PTR5), .B(di1_PTR5), .S(_01837__PTR4), .Z(_01920__PTR37) );
  MUX2_X1 U6657 ( .A(_01958__PTR6), .B(di1_PTR6), .S(_01837__PTR4), .Z(_01920__PTR38) );
  MUX2_X1 U6658 ( .A(_01958__PTR7), .B(di1_PTR7), .S(_01837__PTR4), .Z(_01920__PTR39) );
  MUX2_X1 U6659 ( .A(_01957__PTR0), .B(di1_PTR0), .S(_01837__PTR5), .Z(_01918__PTR32) );
  MUX2_X1 U6660 ( .A(_01957__PTR1), .B(di1_PTR1), .S(_01837__PTR5), .Z(_01918__PTR33) );
  MUX2_X1 U6661 ( .A(_01957__PTR2), .B(di1_PTR2), .S(_01837__PTR5), .Z(_01918__PTR34) );
  MUX2_X1 U6662 ( .A(_01957__PTR3), .B(di1_PTR3), .S(_01837__PTR5), .Z(_01918__PTR35) );
  MUX2_X1 U6663 ( .A(_01957__PTR4), .B(di1_PTR4), .S(_01837__PTR5), .Z(_01918__PTR36) );
  MUX2_X1 U6664 ( .A(_01957__PTR5), .B(di1_PTR5), .S(_01837__PTR5), .Z(_01918__PTR37) );
  MUX2_X1 U6665 ( .A(_01957__PTR6), .B(di1_PTR6), .S(_01837__PTR5), .Z(_01918__PTR38) );
  MUX2_X1 U6666 ( .A(_01957__PTR7), .B(di1_PTR7), .S(_01837__PTR5), .Z(_01918__PTR39) );
  MUX2_X1 U6667 ( .A(_01956__PTR0), .B(di1_PTR0), .S(_01837__PTR6), .Z(_01916__PTR32) );
  MUX2_X1 U6668 ( .A(_01956__PTR1), .B(di1_PTR1), .S(_01837__PTR6), .Z(_01916__PTR33) );
  MUX2_X1 U6669 ( .A(_01956__PTR2), .B(di1_PTR2), .S(_01837__PTR6), .Z(_01916__PTR34) );
  MUX2_X1 U6670 ( .A(_01956__PTR3), .B(di1_PTR3), .S(_01837__PTR6), .Z(_01916__PTR35) );
  MUX2_X1 U6671 ( .A(_01956__PTR4), .B(di1_PTR4), .S(_01837__PTR6), .Z(_01916__PTR36) );
  MUX2_X1 U6672 ( .A(_01956__PTR5), .B(di1_PTR5), .S(_01837__PTR6), .Z(_01916__PTR37) );
  MUX2_X1 U6673 ( .A(_01956__PTR6), .B(di1_PTR6), .S(_01837__PTR6), .Z(_01916__PTR38) );
  MUX2_X1 U6674 ( .A(_01956__PTR7), .B(di1_PTR7), .S(_01837__PTR6), .Z(_01916__PTR39) );
  MUX2_X1 U6675 ( .A(_01955__PTR0), .B(di1_PTR0), .S(_01837__PTR7), .Z(_01914__PTR32) );
  MUX2_X1 U6676 ( .A(_01955__PTR1), .B(di1_PTR1), .S(_01837__PTR7), .Z(_01914__PTR33) );
  MUX2_X1 U6677 ( .A(_01955__PTR2), .B(di1_PTR2), .S(_01837__PTR7), .Z(_01914__PTR34) );
  MUX2_X1 U6678 ( .A(_01955__PTR3), .B(di1_PTR3), .S(_01837__PTR7), .Z(_01914__PTR35) );
  MUX2_X1 U6679 ( .A(_01955__PTR4), .B(di1_PTR4), .S(_01837__PTR7), .Z(_01914__PTR36) );
  MUX2_X1 U6680 ( .A(_01955__PTR5), .B(di1_PTR5), .S(_01837__PTR7), .Z(_01914__PTR37) );
  MUX2_X1 U6681 ( .A(_01955__PTR6), .B(di1_PTR6), .S(_01837__PTR7), .Z(_01914__PTR38) );
  MUX2_X1 U6682 ( .A(_01955__PTR7), .B(di1_PTR7), .S(_01837__PTR7), .Z(_01914__PTR39) );
  MUX2_X1 U6683 ( .A(_01954__PTR0), .B(di1_PTR0), .S(_01837__PTR8), .Z(_01912__PTR32) );
  MUX2_X1 U6684 ( .A(_01954__PTR1), .B(di1_PTR1), .S(_01837__PTR8), .Z(_01912__PTR33) );
  MUX2_X1 U6685 ( .A(_01954__PTR2), .B(di1_PTR2), .S(_01837__PTR8), .Z(_01912__PTR34) );
  MUX2_X1 U6686 ( .A(_01954__PTR3), .B(di1_PTR3), .S(_01837__PTR8), .Z(_01912__PTR35) );
  MUX2_X1 U6687 ( .A(_01954__PTR4), .B(di1_PTR4), .S(_01837__PTR8), .Z(_01912__PTR36) );
  MUX2_X1 U6688 ( .A(_01954__PTR5), .B(di1_PTR5), .S(_01837__PTR8), .Z(_01912__PTR37) );
  MUX2_X1 U6689 ( .A(_01954__PTR6), .B(di1_PTR6), .S(_01837__PTR8), .Z(_01912__PTR38) );
  MUX2_X1 U6690 ( .A(_01954__PTR7), .B(di1_PTR7), .S(_01837__PTR8), .Z(_01912__PTR39) );
  MUX2_X1 U6691 ( .A(_01953__PTR0), .B(di1_PTR0), .S(_01837__PTR9), .Z(_01910__PTR32) );
  MUX2_X1 U6692 ( .A(_01953__PTR1), .B(di1_PTR1), .S(_01837__PTR9), .Z(_01910__PTR33) );
  MUX2_X1 U6693 ( .A(_01953__PTR2), .B(di1_PTR2), .S(_01837__PTR9), .Z(_01910__PTR34) );
  MUX2_X1 U6694 ( .A(_01953__PTR3), .B(di1_PTR3), .S(_01837__PTR9), .Z(_01910__PTR35) );
  MUX2_X1 U6695 ( .A(_01953__PTR4), .B(di1_PTR4), .S(_01837__PTR9), .Z(_01910__PTR36) );
  MUX2_X1 U6696 ( .A(_01953__PTR5), .B(di1_PTR5), .S(_01837__PTR9), .Z(_01910__PTR37) );
  MUX2_X1 U6697 ( .A(_01953__PTR6), .B(di1_PTR6), .S(_01837__PTR9), .Z(_01910__PTR38) );
  MUX2_X1 U6698 ( .A(_01953__PTR7), .B(di1_PTR7), .S(_01837__PTR9), .Z(_01910__PTR39) );
  MUX2_X1 U6699 ( .A(_01952__PTR0), .B(di1_PTR0), .S(_01837__PTR10), .Z(_01908__PTR32) );
  MUX2_X1 U6700 ( .A(_01952__PTR1), .B(di1_PTR1), .S(_01837__PTR10), .Z(_01908__PTR33) );
  MUX2_X1 U6701 ( .A(_01952__PTR2), .B(di1_PTR2), .S(_01837__PTR10), .Z(_01908__PTR34) );
  MUX2_X1 U6702 ( .A(_01952__PTR3), .B(di1_PTR3), .S(_01837__PTR10), .Z(_01908__PTR35) );
  MUX2_X1 U6703 ( .A(_01952__PTR4), .B(di1_PTR4), .S(_01837__PTR10), .Z(_01908__PTR36) );
  MUX2_X1 U6704 ( .A(_01952__PTR5), .B(di1_PTR5), .S(_01837__PTR10), .Z(_01908__PTR37) );
  MUX2_X1 U6705 ( .A(_01952__PTR6), .B(di1_PTR6), .S(_01837__PTR10), .Z(_01908__PTR38) );
  MUX2_X1 U6706 ( .A(_01952__PTR7), .B(di1_PTR7), .S(_01837__PTR10), .Z(_01908__PTR39) );
  MUX2_X1 U6707 ( .A(_01951__PTR0), .B(di1_PTR0), .S(_01837__PTR11), .Z(_01906__PTR32) );
  MUX2_X1 U6708 ( .A(_01951__PTR1), .B(di1_PTR1), .S(_01837__PTR11), .Z(_01906__PTR33) );
  MUX2_X1 U6709 ( .A(_01951__PTR2), .B(di1_PTR2), .S(_01837__PTR11), .Z(_01906__PTR34) );
  MUX2_X1 U6710 ( .A(_01951__PTR3), .B(di1_PTR3), .S(_01837__PTR11), .Z(_01906__PTR35) );
  MUX2_X1 U6711 ( .A(_01951__PTR4), .B(di1_PTR4), .S(_01837__PTR11), .Z(_01906__PTR36) );
  MUX2_X1 U6712 ( .A(_01951__PTR5), .B(di1_PTR5), .S(_01837__PTR11), .Z(_01906__PTR37) );
  MUX2_X1 U6713 ( .A(_01951__PTR6), .B(di1_PTR6), .S(_01837__PTR11), .Z(_01906__PTR38) );
  MUX2_X1 U6714 ( .A(_01951__PTR7), .B(di1_PTR7), .S(_01837__PTR11), .Z(_01906__PTR39) );
  MUX2_X1 U6715 ( .A(_01950__PTR0), .B(di1_PTR0), .S(_01837__PTR12), .Z(_01904__PTR32) );
  MUX2_X1 U6716 ( .A(_01950__PTR1), .B(di1_PTR1), .S(_01837__PTR12), .Z(_01904__PTR33) );
  MUX2_X1 U6717 ( .A(_01950__PTR2), .B(di1_PTR2), .S(_01837__PTR12), .Z(_01904__PTR34) );
  MUX2_X1 U6718 ( .A(_01950__PTR3), .B(di1_PTR3), .S(_01837__PTR12), .Z(_01904__PTR35) );
  MUX2_X1 U6719 ( .A(_01950__PTR4), .B(di1_PTR4), .S(_01837__PTR12), .Z(_01904__PTR36) );
  MUX2_X1 U6720 ( .A(_01950__PTR5), .B(di1_PTR5), .S(_01837__PTR12), .Z(_01904__PTR37) );
  MUX2_X1 U6721 ( .A(_01950__PTR6), .B(di1_PTR6), .S(_01837__PTR12), .Z(_01904__PTR38) );
  MUX2_X1 U6722 ( .A(_01950__PTR7), .B(di1_PTR7), .S(_01837__PTR12), .Z(_01904__PTR39) );
  MUX2_X1 U6723 ( .A(_01949__PTR0), .B(di1_PTR0), .S(_01837__PTR13), .Z(_01902__PTR32) );
  MUX2_X1 U6724 ( .A(_01949__PTR1), .B(di1_PTR1), .S(_01837__PTR13), .Z(_01902__PTR33) );
  MUX2_X1 U6725 ( .A(_01949__PTR2), .B(di1_PTR2), .S(_01837__PTR13), .Z(_01902__PTR34) );
  MUX2_X1 U6726 ( .A(_01949__PTR3), .B(di1_PTR3), .S(_01837__PTR13), .Z(_01902__PTR35) );
  MUX2_X1 U6727 ( .A(_01949__PTR4), .B(di1_PTR4), .S(_01837__PTR13), .Z(_01902__PTR36) );
  MUX2_X1 U6728 ( .A(_01949__PTR5), .B(di1_PTR5), .S(_01837__PTR13), .Z(_01902__PTR37) );
  MUX2_X1 U6729 ( .A(_01949__PTR6), .B(di1_PTR6), .S(_01837__PTR13), .Z(_01902__PTR38) );
  MUX2_X1 U6730 ( .A(_01949__PTR7), .B(di1_PTR7), .S(_01837__PTR13), .Z(_01902__PTR39) );
  MUX2_X1 U6731 ( .A(_01948__PTR0), .B(di1_PTR0), .S(_01837__PTR14), .Z(_01900__PTR32) );
  MUX2_X1 U6732 ( .A(_01948__PTR1), .B(di1_PTR1), .S(_01837__PTR14), .Z(_01900__PTR33) );
  MUX2_X1 U6733 ( .A(_01948__PTR2), .B(di1_PTR2), .S(_01837__PTR14), .Z(_01900__PTR34) );
  MUX2_X1 U6734 ( .A(_01948__PTR3), .B(di1_PTR3), .S(_01837__PTR14), .Z(_01900__PTR35) );
  MUX2_X1 U6735 ( .A(_01948__PTR4), .B(di1_PTR4), .S(_01837__PTR14), .Z(_01900__PTR36) );
  MUX2_X1 U6736 ( .A(_01948__PTR5), .B(di1_PTR5), .S(_01837__PTR14), .Z(_01900__PTR37) );
  MUX2_X1 U6737 ( .A(_01948__PTR6), .B(di1_PTR6), .S(_01837__PTR14), .Z(_01900__PTR38) );
  MUX2_X1 U6738 ( .A(_01948__PTR7), .B(di1_PTR7), .S(_01837__PTR14), .Z(_01900__PTR39) );
  MUX2_X1 U6739 ( .A(_01947__PTR0), .B(di1_PTR0), .S(_01837__PTR15), .Z(_01898__PTR32) );
  MUX2_X1 U6740 ( .A(_01947__PTR1), .B(di1_PTR1), .S(_01837__PTR15), .Z(_01898__PTR33) );
  MUX2_X1 U6741 ( .A(_01947__PTR2), .B(di1_PTR2), .S(_01837__PTR15), .Z(_01898__PTR34) );
  MUX2_X1 U6742 ( .A(_01947__PTR3), .B(di1_PTR3), .S(_01837__PTR15), .Z(_01898__PTR35) );
  MUX2_X1 U6743 ( .A(_01947__PTR4), .B(di1_PTR4), .S(_01837__PTR15), .Z(_01898__PTR36) );
  MUX2_X1 U6744 ( .A(_01947__PTR5), .B(di1_PTR5), .S(_01837__PTR15), .Z(_01898__PTR37) );
  MUX2_X1 U6745 ( .A(_01947__PTR6), .B(di1_PTR6), .S(_01837__PTR15), .Z(_01898__PTR38) );
  MUX2_X1 U6746 ( .A(_01947__PTR7), .B(di1_PTR7), .S(_01837__PTR15), .Z(_01898__PTR39) );
  MUX2_X1 U6747 ( .A(P1_P1_InstQueue_PTR0_PTR0), .B(di1_PTR0), .S(_01835__PTR0), .Z(_01962__PTR0) );
  MUX2_X1 U6748 ( .A(P1_P1_InstQueue_PTR0_PTR1), .B(di1_PTR1), .S(_01835__PTR0), .Z(_01962__PTR1) );
  MUX2_X1 U6749 ( .A(P1_P1_InstQueue_PTR0_PTR2), .B(di1_PTR2), .S(_01835__PTR0), .Z(_01962__PTR2) );
  MUX2_X1 U6750 ( .A(P1_P1_InstQueue_PTR0_PTR3), .B(di1_PTR3), .S(_01835__PTR0), .Z(_01962__PTR3) );
  MUX2_X1 U6751 ( .A(P1_P1_InstQueue_PTR0_PTR4), .B(di1_PTR4), .S(_01835__PTR0), .Z(_01962__PTR4) );
  MUX2_X1 U6752 ( .A(P1_P1_InstQueue_PTR0_PTR5), .B(di1_PTR5), .S(_01835__PTR0), .Z(_01962__PTR5) );
  MUX2_X1 U6753 ( .A(P1_P1_InstQueue_PTR0_PTR6), .B(di1_PTR6), .S(_01835__PTR0), .Z(_01962__PTR6) );
  MUX2_X1 U6754 ( .A(P1_P1_InstQueue_PTR0_PTR7), .B(di1_PTR7), .S(_01835__PTR0), .Z(_01962__PTR7) );
  MUX2_X1 U6755 ( .A(P1_P1_InstQueue_PTR1_PTR0), .B(di1_PTR0), .S(_01835__PTR1), .Z(_01961__PTR0) );
  MUX2_X1 U6756 ( .A(P1_P1_InstQueue_PTR1_PTR1), .B(di1_PTR1), .S(_01835__PTR1), .Z(_01961__PTR1) );
  MUX2_X1 U6757 ( .A(P1_P1_InstQueue_PTR1_PTR2), .B(di1_PTR2), .S(_01835__PTR1), .Z(_01961__PTR2) );
  MUX2_X1 U6758 ( .A(P1_P1_InstQueue_PTR1_PTR3), .B(di1_PTR3), .S(_01835__PTR1), .Z(_01961__PTR3) );
  MUX2_X1 U6759 ( .A(P1_P1_InstQueue_PTR1_PTR4), .B(di1_PTR4), .S(_01835__PTR1), .Z(_01961__PTR4) );
  MUX2_X1 U6760 ( .A(P1_P1_InstQueue_PTR1_PTR5), .B(di1_PTR5), .S(_01835__PTR1), .Z(_01961__PTR5) );
  MUX2_X1 U6761 ( .A(P1_P1_InstQueue_PTR1_PTR6), .B(di1_PTR6), .S(_01835__PTR1), .Z(_01961__PTR6) );
  MUX2_X1 U6762 ( .A(P1_P1_InstQueue_PTR1_PTR7), .B(di1_PTR7), .S(_01835__PTR1), .Z(_01961__PTR7) );
  MUX2_X1 U6763 ( .A(P1_P1_InstQueue_PTR2_PTR0), .B(di1_PTR0), .S(_01835__PTR2), .Z(_01960__PTR0) );
  MUX2_X1 U6764 ( .A(P1_P1_InstQueue_PTR2_PTR1), .B(di1_PTR1), .S(_01835__PTR2), .Z(_01960__PTR1) );
  MUX2_X1 U6765 ( .A(P1_P1_InstQueue_PTR2_PTR2), .B(di1_PTR2), .S(_01835__PTR2), .Z(_01960__PTR2) );
  MUX2_X1 U6766 ( .A(P1_P1_InstQueue_PTR2_PTR3), .B(di1_PTR3), .S(_01835__PTR2), .Z(_01960__PTR3) );
  MUX2_X1 U6767 ( .A(P1_P1_InstQueue_PTR2_PTR4), .B(di1_PTR4), .S(_01835__PTR2), .Z(_01960__PTR4) );
  MUX2_X1 U6768 ( .A(P1_P1_InstQueue_PTR2_PTR5), .B(di1_PTR5), .S(_01835__PTR2), .Z(_01960__PTR5) );
  MUX2_X1 U6769 ( .A(P1_P1_InstQueue_PTR2_PTR6), .B(di1_PTR6), .S(_01835__PTR2), .Z(_01960__PTR6) );
  MUX2_X1 U6770 ( .A(P1_P1_InstQueue_PTR2_PTR7), .B(di1_PTR7), .S(_01835__PTR2), .Z(_01960__PTR7) );
  MUX2_X1 U6771 ( .A(P1_P1_InstQueue_PTR3_PTR0), .B(di1_PTR0), .S(_01835__PTR3), .Z(_01959__PTR0) );
  MUX2_X1 U6772 ( .A(P1_P1_InstQueue_PTR3_PTR1), .B(di1_PTR1), .S(_01835__PTR3), .Z(_01959__PTR1) );
  MUX2_X1 U6773 ( .A(P1_P1_InstQueue_PTR3_PTR2), .B(di1_PTR2), .S(_01835__PTR3), .Z(_01959__PTR2) );
  MUX2_X1 U6774 ( .A(P1_P1_InstQueue_PTR3_PTR3), .B(di1_PTR3), .S(_01835__PTR3), .Z(_01959__PTR3) );
  MUX2_X1 U6775 ( .A(P1_P1_InstQueue_PTR3_PTR4), .B(di1_PTR4), .S(_01835__PTR3), .Z(_01959__PTR4) );
  MUX2_X1 U6776 ( .A(P1_P1_InstQueue_PTR3_PTR5), .B(di1_PTR5), .S(_01835__PTR3), .Z(_01959__PTR5) );
  MUX2_X1 U6777 ( .A(P1_P1_InstQueue_PTR3_PTR6), .B(di1_PTR6), .S(_01835__PTR3), .Z(_01959__PTR6) );
  MUX2_X1 U6778 ( .A(P1_P1_InstQueue_PTR3_PTR7), .B(di1_PTR7), .S(_01835__PTR3), .Z(_01959__PTR7) );
  MUX2_X1 U6779 ( .A(P1_P1_InstQueue_PTR4_PTR0), .B(di1_PTR0), .S(_01835__PTR4), .Z(_01958__PTR0) );
  MUX2_X1 U6780 ( .A(P1_P1_InstQueue_PTR4_PTR1), .B(di1_PTR1), .S(_01835__PTR4), .Z(_01958__PTR1) );
  MUX2_X1 U6781 ( .A(P1_P1_InstQueue_PTR4_PTR2), .B(di1_PTR2), .S(_01835__PTR4), .Z(_01958__PTR2) );
  MUX2_X1 U6782 ( .A(P1_P1_InstQueue_PTR4_PTR3), .B(di1_PTR3), .S(_01835__PTR4), .Z(_01958__PTR3) );
  MUX2_X1 U6783 ( .A(P1_P1_InstQueue_PTR4_PTR4), .B(di1_PTR4), .S(_01835__PTR4), .Z(_01958__PTR4) );
  MUX2_X1 U6784 ( .A(P1_P1_InstQueue_PTR4_PTR5), .B(di1_PTR5), .S(_01835__PTR4), .Z(_01958__PTR5) );
  MUX2_X1 U6785 ( .A(P1_P1_InstQueue_PTR4_PTR6), .B(di1_PTR6), .S(_01835__PTR4), .Z(_01958__PTR6) );
  MUX2_X1 U6786 ( .A(P1_P1_InstQueue_PTR4_PTR7), .B(di1_PTR7), .S(_01835__PTR4), .Z(_01958__PTR7) );
  MUX2_X1 U6787 ( .A(P1_P1_InstQueue_PTR5_PTR0), .B(di1_PTR0), .S(_01835__PTR5), .Z(_01957__PTR0) );
  MUX2_X1 U6788 ( .A(P1_P1_InstQueue_PTR5_PTR1), .B(di1_PTR1), .S(_01835__PTR5), .Z(_01957__PTR1) );
  MUX2_X1 U6789 ( .A(P1_P1_InstQueue_PTR5_PTR2), .B(di1_PTR2), .S(_01835__PTR5), .Z(_01957__PTR2) );
  MUX2_X1 U6790 ( .A(P1_P1_InstQueue_PTR5_PTR3), .B(di1_PTR3), .S(_01835__PTR5), .Z(_01957__PTR3) );
  MUX2_X1 U6791 ( .A(P1_P1_InstQueue_PTR5_PTR4), .B(di1_PTR4), .S(_01835__PTR5), .Z(_01957__PTR4) );
  MUX2_X1 U6792 ( .A(P1_P1_InstQueue_PTR5_PTR5), .B(di1_PTR5), .S(_01835__PTR5), .Z(_01957__PTR5) );
  MUX2_X1 U6793 ( .A(P1_P1_InstQueue_PTR5_PTR6), .B(di1_PTR6), .S(_01835__PTR5), .Z(_01957__PTR6) );
  MUX2_X1 U6794 ( .A(P1_P1_InstQueue_PTR5_PTR7), .B(di1_PTR7), .S(_01835__PTR5), .Z(_01957__PTR7) );
  MUX2_X1 U6795 ( .A(P1_P1_InstQueue_PTR6_PTR0), .B(di1_PTR0), .S(_01835__PTR6), .Z(_01956__PTR0) );
  MUX2_X1 U6796 ( .A(P1_P1_InstQueue_PTR6_PTR1), .B(di1_PTR1), .S(_01835__PTR6), .Z(_01956__PTR1) );
  MUX2_X1 U6797 ( .A(P1_P1_InstQueue_PTR6_PTR2), .B(di1_PTR2), .S(_01835__PTR6), .Z(_01956__PTR2) );
  MUX2_X1 U6798 ( .A(P1_P1_InstQueue_PTR6_PTR3), .B(di1_PTR3), .S(_01835__PTR6), .Z(_01956__PTR3) );
  MUX2_X1 U6799 ( .A(P1_P1_InstQueue_PTR6_PTR4), .B(di1_PTR4), .S(_01835__PTR6), .Z(_01956__PTR4) );
  MUX2_X1 U6800 ( .A(P1_P1_InstQueue_PTR6_PTR5), .B(di1_PTR5), .S(_01835__PTR6), .Z(_01956__PTR5) );
  MUX2_X1 U6801 ( .A(P1_P1_InstQueue_PTR6_PTR6), .B(di1_PTR6), .S(_01835__PTR6), .Z(_01956__PTR6) );
  MUX2_X1 U6802 ( .A(P1_P1_InstQueue_PTR6_PTR7), .B(di1_PTR7), .S(_01835__PTR6), .Z(_01956__PTR7) );
  MUX2_X1 U6803 ( .A(P1_P1_InstQueue_PTR7_PTR0), .B(di1_PTR0), .S(_01835__PTR7), .Z(_01955__PTR0) );
  MUX2_X1 U6804 ( .A(P1_P1_InstQueue_PTR7_PTR1), .B(di1_PTR1), .S(_01835__PTR7), .Z(_01955__PTR1) );
  MUX2_X1 U6805 ( .A(P1_P1_InstQueue_PTR7_PTR2), .B(di1_PTR2), .S(_01835__PTR7), .Z(_01955__PTR2) );
  MUX2_X1 U6806 ( .A(P1_P1_InstQueue_PTR7_PTR3), .B(di1_PTR3), .S(_01835__PTR7), .Z(_01955__PTR3) );
  MUX2_X1 U6807 ( .A(P1_P1_InstQueue_PTR7_PTR4), .B(di1_PTR4), .S(_01835__PTR7), .Z(_01955__PTR4) );
  MUX2_X1 U6808 ( .A(P1_P1_InstQueue_PTR7_PTR5), .B(di1_PTR5), .S(_01835__PTR7), .Z(_01955__PTR5) );
  MUX2_X1 U6809 ( .A(P1_P1_InstQueue_PTR7_PTR6), .B(di1_PTR6), .S(_01835__PTR7), .Z(_01955__PTR6) );
  MUX2_X1 U6810 ( .A(P1_P1_InstQueue_PTR7_PTR7), .B(di1_PTR7), .S(_01835__PTR7), .Z(_01955__PTR7) );
  MUX2_X1 U6811 ( .A(P1_P1_InstQueue_PTR8_PTR0), .B(di1_PTR0), .S(_01835__PTR8), .Z(_01954__PTR0) );
  MUX2_X1 U6812 ( .A(P1_P1_InstQueue_PTR8_PTR1), .B(di1_PTR1), .S(_01835__PTR8), .Z(_01954__PTR1) );
  MUX2_X1 U6813 ( .A(P1_P1_InstQueue_PTR8_PTR2), .B(di1_PTR2), .S(_01835__PTR8), .Z(_01954__PTR2) );
  MUX2_X1 U6814 ( .A(P1_P1_InstQueue_PTR8_PTR3), .B(di1_PTR3), .S(_01835__PTR8), .Z(_01954__PTR3) );
  MUX2_X1 U6815 ( .A(P1_P1_InstQueue_PTR8_PTR4), .B(di1_PTR4), .S(_01835__PTR8), .Z(_01954__PTR4) );
  MUX2_X1 U6816 ( .A(P1_P1_InstQueue_PTR8_PTR5), .B(di1_PTR5), .S(_01835__PTR8), .Z(_01954__PTR5) );
  MUX2_X1 U6817 ( .A(P1_P1_InstQueue_PTR8_PTR6), .B(di1_PTR6), .S(_01835__PTR8), .Z(_01954__PTR6) );
  MUX2_X1 U6818 ( .A(P1_P1_InstQueue_PTR8_PTR7), .B(di1_PTR7), .S(_01835__PTR8), .Z(_01954__PTR7) );
  MUX2_X1 U6819 ( .A(P1_P1_InstQueue_PTR9_PTR0), .B(di1_PTR0), .S(_01835__PTR9), .Z(_01953__PTR0) );
  MUX2_X1 U6820 ( .A(P1_P1_InstQueue_PTR9_PTR1), .B(di1_PTR1), .S(_01835__PTR9), .Z(_01953__PTR1) );
  MUX2_X1 U6821 ( .A(P1_P1_InstQueue_PTR9_PTR2), .B(di1_PTR2), .S(_01835__PTR9), .Z(_01953__PTR2) );
  MUX2_X1 U6822 ( .A(P1_P1_InstQueue_PTR9_PTR3), .B(di1_PTR3), .S(_01835__PTR9), .Z(_01953__PTR3) );
  MUX2_X1 U6823 ( .A(P1_P1_InstQueue_PTR9_PTR4), .B(di1_PTR4), .S(_01835__PTR9), .Z(_01953__PTR4) );
  MUX2_X1 U6824 ( .A(P1_P1_InstQueue_PTR9_PTR5), .B(di1_PTR5), .S(_01835__PTR9), .Z(_01953__PTR5) );
  MUX2_X1 U6825 ( .A(P1_P1_InstQueue_PTR9_PTR6), .B(di1_PTR6), .S(_01835__PTR9), .Z(_01953__PTR6) );
  MUX2_X1 U6826 ( .A(P1_P1_InstQueue_PTR9_PTR7), .B(di1_PTR7), .S(_01835__PTR9), .Z(_01953__PTR7) );
  MUX2_X1 U6827 ( .A(P1_P1_InstQueue_PTR10_PTR0), .B(di1_PTR0), .S(_01835__PTR10), .Z(_01952__PTR0) );
  MUX2_X1 U6828 ( .A(P1_P1_InstQueue_PTR10_PTR1), .B(di1_PTR1), .S(_01835__PTR10), .Z(_01952__PTR1) );
  MUX2_X1 U6829 ( .A(P1_P1_InstQueue_PTR10_PTR2), .B(di1_PTR2), .S(_01835__PTR10), .Z(_01952__PTR2) );
  MUX2_X1 U6830 ( .A(P1_P1_InstQueue_PTR10_PTR3), .B(di1_PTR3), .S(_01835__PTR10), .Z(_01952__PTR3) );
  MUX2_X1 U6831 ( .A(P1_P1_InstQueue_PTR10_PTR4), .B(di1_PTR4), .S(_01835__PTR10), .Z(_01952__PTR4) );
  MUX2_X1 U6832 ( .A(P1_P1_InstQueue_PTR10_PTR5), .B(di1_PTR5), .S(_01835__PTR10), .Z(_01952__PTR5) );
  MUX2_X1 U6833 ( .A(P1_P1_InstQueue_PTR10_PTR6), .B(di1_PTR6), .S(_01835__PTR10), .Z(_01952__PTR6) );
  MUX2_X1 U6834 ( .A(P1_P1_InstQueue_PTR10_PTR7), .B(di1_PTR7), .S(_01835__PTR10), .Z(_01952__PTR7) );
  MUX2_X1 U6835 ( .A(P1_P1_InstQueue_PTR11_PTR0), .B(di1_PTR0), .S(_01835__PTR11), .Z(_01951__PTR0) );
  MUX2_X1 U6836 ( .A(P1_P1_InstQueue_PTR11_PTR1), .B(di1_PTR1), .S(_01835__PTR11), .Z(_01951__PTR1) );
  MUX2_X1 U6837 ( .A(P1_P1_InstQueue_PTR11_PTR2), .B(di1_PTR2), .S(_01835__PTR11), .Z(_01951__PTR2) );
  MUX2_X1 U6838 ( .A(P1_P1_InstQueue_PTR11_PTR3), .B(di1_PTR3), .S(_01835__PTR11), .Z(_01951__PTR3) );
  MUX2_X1 U6839 ( .A(P1_P1_InstQueue_PTR11_PTR4), .B(di1_PTR4), .S(_01835__PTR11), .Z(_01951__PTR4) );
  MUX2_X1 U6840 ( .A(P1_P1_InstQueue_PTR11_PTR5), .B(di1_PTR5), .S(_01835__PTR11), .Z(_01951__PTR5) );
  MUX2_X1 U6841 ( .A(P1_P1_InstQueue_PTR11_PTR6), .B(di1_PTR6), .S(_01835__PTR11), .Z(_01951__PTR6) );
  MUX2_X1 U6842 ( .A(P1_P1_InstQueue_PTR11_PTR7), .B(di1_PTR7), .S(_01835__PTR11), .Z(_01951__PTR7) );
  MUX2_X1 U6843 ( .A(P1_P1_InstQueue_PTR12_PTR0), .B(di1_PTR0), .S(_01835__PTR12), .Z(_01950__PTR0) );
  MUX2_X1 U6844 ( .A(P1_P1_InstQueue_PTR12_PTR1), .B(di1_PTR1), .S(_01835__PTR12), .Z(_01950__PTR1) );
  MUX2_X1 U6845 ( .A(P1_P1_InstQueue_PTR12_PTR2), .B(di1_PTR2), .S(_01835__PTR12), .Z(_01950__PTR2) );
  MUX2_X1 U6846 ( .A(P1_P1_InstQueue_PTR12_PTR3), .B(di1_PTR3), .S(_01835__PTR12), .Z(_01950__PTR3) );
  MUX2_X1 U6847 ( .A(P1_P1_InstQueue_PTR12_PTR4), .B(di1_PTR4), .S(_01835__PTR12), .Z(_01950__PTR4) );
  MUX2_X1 U6848 ( .A(P1_P1_InstQueue_PTR12_PTR5), .B(di1_PTR5), .S(_01835__PTR12), .Z(_01950__PTR5) );
  MUX2_X1 U6849 ( .A(P1_P1_InstQueue_PTR12_PTR6), .B(di1_PTR6), .S(_01835__PTR12), .Z(_01950__PTR6) );
  MUX2_X1 U6850 ( .A(P1_P1_InstQueue_PTR12_PTR7), .B(di1_PTR7), .S(_01835__PTR12), .Z(_01950__PTR7) );
  MUX2_X1 U6851 ( .A(P1_P1_InstQueue_PTR13_PTR0), .B(di1_PTR0), .S(_01835__PTR13), .Z(_01949__PTR0) );
  MUX2_X1 U6852 ( .A(P1_P1_InstQueue_PTR13_PTR1), .B(di1_PTR1), .S(_01835__PTR13), .Z(_01949__PTR1) );
  MUX2_X1 U6853 ( .A(P1_P1_InstQueue_PTR13_PTR2), .B(di1_PTR2), .S(_01835__PTR13), .Z(_01949__PTR2) );
  MUX2_X1 U6854 ( .A(P1_P1_InstQueue_PTR13_PTR3), .B(di1_PTR3), .S(_01835__PTR13), .Z(_01949__PTR3) );
  MUX2_X1 U6855 ( .A(P1_P1_InstQueue_PTR13_PTR4), .B(di1_PTR4), .S(_01835__PTR13), .Z(_01949__PTR4) );
  MUX2_X1 U6856 ( .A(P1_P1_InstQueue_PTR13_PTR5), .B(di1_PTR5), .S(_01835__PTR13), .Z(_01949__PTR5) );
  MUX2_X1 U6857 ( .A(P1_P1_InstQueue_PTR13_PTR6), .B(di1_PTR6), .S(_01835__PTR13), .Z(_01949__PTR6) );
  MUX2_X1 U6858 ( .A(P1_P1_InstQueue_PTR13_PTR7), .B(di1_PTR7), .S(_01835__PTR13), .Z(_01949__PTR7) );
  MUX2_X1 U6859 ( .A(P1_P1_InstQueue_PTR14_PTR0), .B(di1_PTR0), .S(_01835__PTR14), .Z(_01948__PTR0) );
  MUX2_X1 U6860 ( .A(P1_P1_InstQueue_PTR14_PTR1), .B(di1_PTR1), .S(_01835__PTR14), .Z(_01948__PTR1) );
  MUX2_X1 U6861 ( .A(P1_P1_InstQueue_PTR14_PTR2), .B(di1_PTR2), .S(_01835__PTR14), .Z(_01948__PTR2) );
  MUX2_X1 U6862 ( .A(P1_P1_InstQueue_PTR14_PTR3), .B(di1_PTR3), .S(_01835__PTR14), .Z(_01948__PTR3) );
  MUX2_X1 U6863 ( .A(P1_P1_InstQueue_PTR14_PTR4), .B(di1_PTR4), .S(_01835__PTR14), .Z(_01948__PTR4) );
  MUX2_X1 U6864 ( .A(P1_P1_InstQueue_PTR14_PTR5), .B(di1_PTR5), .S(_01835__PTR14), .Z(_01948__PTR5) );
  MUX2_X1 U6865 ( .A(P1_P1_InstQueue_PTR14_PTR6), .B(di1_PTR6), .S(_01835__PTR14), .Z(_01948__PTR6) );
  MUX2_X1 U6866 ( .A(P1_P1_InstQueue_PTR14_PTR7), .B(di1_PTR7), .S(_01835__PTR14), .Z(_01948__PTR7) );
  MUX2_X1 U6867 ( .A(P1_P1_InstQueue_PTR15_PTR0), .B(di1_PTR0), .S(_01835__PTR15), .Z(_01947__PTR0) );
  MUX2_X1 U6868 ( .A(P1_P1_InstQueue_PTR15_PTR1), .B(di1_PTR1), .S(_01835__PTR15), .Z(_01947__PTR1) );
  MUX2_X1 U6869 ( .A(P1_P1_InstQueue_PTR15_PTR2), .B(di1_PTR2), .S(_01835__PTR15), .Z(_01947__PTR2) );
  MUX2_X1 U6870 ( .A(P1_P1_InstQueue_PTR15_PTR3), .B(di1_PTR3), .S(_01835__PTR15), .Z(_01947__PTR3) );
  MUX2_X1 U6871 ( .A(P1_P1_InstQueue_PTR15_PTR4), .B(di1_PTR4), .S(_01835__PTR15), .Z(_01947__PTR4) );
  MUX2_X1 U6872 ( .A(P1_P1_InstQueue_PTR15_PTR5), .B(di1_PTR5), .S(_01835__PTR15), .Z(_01947__PTR5) );
  MUX2_X1 U6873 ( .A(P1_P1_InstQueue_PTR15_PTR6), .B(di1_PTR6), .S(_01835__PTR15), .Z(_01947__PTR6) );
  MUX2_X1 U6874 ( .A(P1_P1_InstQueue_PTR15_PTR7), .B(di1_PTR7), .S(_01835__PTR15), .Z(_01947__PTR7) );
  MUX2_X1 U6875 ( .A(_01946__PTR0), .B(1'b0), .S(_01941_), .Z(_01876__PTR28) );
  MUX2_X1 U6876 ( .A(_01946__PTR1), .B(1'b1), .S(_01941_), .Z(_01876__PTR29) );
  MUX2_X1 U6877 ( .A(_01946__PTR2), .B(1'b1), .S(_01941_), .Z(_01876__PTR30) );
  MUX2_X1 U6878 ( .A(_01945__PTR0), .B(1'b1), .S(_01942_), .Z(_01946__PTR0) );
  MUX2_X1 U6879 ( .A(_01945__PTR1), .B(1'b0), .S(_01942_), .Z(_01946__PTR1) );
  MUX2_X1 U6880 ( .A(_01945__PTR2), .B(1'b1), .S(_01942_), .Z(_01946__PTR2) );
  INV_X1 U6881 ( .A(_01769__PTR4), .ZN(_01945__PTR0) );
  MUX2_X1 U6882 ( .A(_01944__PTR2), .B(1'b1), .S(_01769__PTR4), .Z(_01945__PTR1) );
  MUX2_X1 U6883 ( .A(_01944__PTR2), .B(1'b0), .S(_01769__PTR4), .Z(_01945__PTR2) );
  INV_X1 U6884 ( .A(_01943_), .ZN(_01944__PTR2) );
  MUX2_X1 U6885 ( .A(P1_EAX_PTR16), .B(_02044__PTR16), .S(_02006_), .Z(_02096__PTR80) );
  MUX2_X1 U6886 ( .A(P1_EAX_PTR17), .B(_02044__PTR17), .S(_02006_), .Z(_02096__PTR81) );
  MUX2_X1 U6887 ( .A(P1_EAX_PTR18), .B(_02044__PTR18), .S(_02006_), .Z(_02096__PTR82) );
  MUX2_X1 U6888 ( .A(P1_EAX_PTR19), .B(_02044__PTR19), .S(_02006_), .Z(_02096__PTR83) );
  MUX2_X1 U6889 ( .A(P1_EAX_PTR20), .B(_02044__PTR20), .S(_02006_), .Z(_02096__PTR84) );
  MUX2_X1 U6890 ( .A(P1_EAX_PTR21), .B(_02044__PTR21), .S(_02006_), .Z(_02096__PTR85) );
  MUX2_X1 U6891 ( .A(P1_EAX_PTR22), .B(_02044__PTR22), .S(_02006_), .Z(_02096__PTR86) );
  MUX2_X1 U6892 ( .A(P1_EAX_PTR23), .B(_02044__PTR23), .S(_02006_), .Z(_02096__PTR87) );
  MUX2_X1 U6893 ( .A(P1_EAX_PTR24), .B(_02044__PTR24), .S(_02006_), .Z(_02096__PTR88) );
  MUX2_X1 U6894 ( .A(P1_EAX_PTR25), .B(_02044__PTR25), .S(_02006_), .Z(_02096__PTR89) );
  MUX2_X1 U6895 ( .A(P1_EAX_PTR26), .B(_02044__PTR26), .S(_02006_), .Z(_02096__PTR90) );
  MUX2_X1 U6896 ( .A(P1_EAX_PTR27), .B(_02044__PTR27), .S(_02006_), .Z(_02096__PTR91) );
  MUX2_X1 U6897 ( .A(P1_EAX_PTR28), .B(_02044__PTR28), .S(_02006_), .Z(_02096__PTR92) );
  MUX2_X1 U6898 ( .A(P1_EAX_PTR29), .B(_02044__PTR29), .S(_02006_), .Z(_02096__PTR93) );
  MUX2_X1 U6899 ( .A(P1_EAX_PTR30), .B(_02044__PTR30), .S(_02006_), .Z(_02096__PTR94) );
  MUX2_X1 U6900 ( .A(P1_EAX_PTR31), .B(_02044__PTR31), .S(_02006_), .Z(_02096__PTR95) );
  MUX2_X1 U6901 ( .A(P1_EAX_PTR0), .B(_02016__PTR0), .S(_02006_), .Z(_02096__PTR96) );
  MUX2_X1 U6902 ( .A(P1_EAX_PTR1), .B(_02016__PTR1), .S(_02006_), .Z(_02096__PTR97) );
  MUX2_X1 U6903 ( .A(P1_EAX_PTR2), .B(_02016__PTR2), .S(_02006_), .Z(_02096__PTR98) );
  MUX2_X1 U6904 ( .A(P1_EAX_PTR3), .B(_02016__PTR3), .S(_02006_), .Z(_02096__PTR99) );
  MUX2_X1 U6905 ( .A(P1_EAX_PTR4), .B(_02016__PTR4), .S(_02006_), .Z(_02096__PTR100) );
  MUX2_X1 U6906 ( .A(P1_EAX_PTR5), .B(_02016__PTR5), .S(_02006_), .Z(_02096__PTR101) );
  MUX2_X1 U6907 ( .A(P1_EAX_PTR6), .B(_02016__PTR6), .S(_02006_), .Z(_02096__PTR102) );
  MUX2_X1 U6908 ( .A(P1_EAX_PTR7), .B(_02016__PTR7), .S(_02006_), .Z(_02096__PTR103) );
  MUX2_X1 U6909 ( .A(P1_EAX_PTR8), .B(_02016__PTR8), .S(_02006_), .Z(_02096__PTR104) );
  MUX2_X1 U6910 ( .A(P1_EAX_PTR9), .B(_02016__PTR9), .S(_02006_), .Z(_02096__PTR105) );
  MUX2_X1 U6911 ( .A(P1_EAX_PTR10), .B(_02016__PTR10), .S(_02006_), .Z(_02096__PTR106) );
  MUX2_X1 U6912 ( .A(P1_EAX_PTR11), .B(_02016__PTR11), .S(_02006_), .Z(_02096__PTR107) );
  MUX2_X1 U6913 ( .A(P1_EAX_PTR12), .B(_02016__PTR12), .S(_02006_), .Z(_02096__PTR108) );
  MUX2_X1 U6914 ( .A(P1_EAX_PTR13), .B(_02016__PTR13), .S(_02006_), .Z(_02096__PTR109) );
  MUX2_X1 U6915 ( .A(P1_EAX_PTR14), .B(_02016__PTR14), .S(_02006_), .Z(_02096__PTR110) );
  MUX2_X1 U6916 ( .A(P1_EAX_PTR15), .B(_02016__PTR15), .S(_02006_), .Z(_02096__PTR111) );
  MUX2_X1 U6917 ( .A(P1_EAX_PTR16), .B(_02016__PTR16), .S(_02006_), .Z(_02096__PTR112) );
  MUX2_X1 U6918 ( .A(P1_EAX_PTR17), .B(_02016__PTR17), .S(_02006_), .Z(_02096__PTR113) );
  MUX2_X1 U6919 ( .A(P1_EAX_PTR18), .B(_02016__PTR18), .S(_02006_), .Z(_02096__PTR114) );
  MUX2_X1 U6920 ( .A(P1_EAX_PTR19), .B(_02016__PTR19), .S(_02006_), .Z(_02096__PTR115) );
  MUX2_X1 U6921 ( .A(P1_EAX_PTR20), .B(_02016__PTR20), .S(_02006_), .Z(_02096__PTR116) );
  MUX2_X1 U6922 ( .A(P1_EAX_PTR21), .B(_02016__PTR21), .S(_02006_), .Z(_02096__PTR117) );
  MUX2_X1 U6923 ( .A(P1_EAX_PTR22), .B(_02016__PTR22), .S(_02006_), .Z(_02096__PTR118) );
  MUX2_X1 U6924 ( .A(P1_EAX_PTR23), .B(_02016__PTR23), .S(_02006_), .Z(_02096__PTR119) );
  MUX2_X1 U6925 ( .A(P1_EAX_PTR24), .B(_02016__PTR24), .S(_02006_), .Z(_02096__PTR120) );
  MUX2_X1 U6926 ( .A(P1_EAX_PTR25), .B(_02016__PTR25), .S(_02006_), .Z(_02096__PTR121) );
  MUX2_X1 U6927 ( .A(P1_EAX_PTR26), .B(_02016__PTR26), .S(_02006_), .Z(_02096__PTR122) );
  MUX2_X1 U6928 ( .A(P1_EAX_PTR27), .B(_02016__PTR27), .S(_02006_), .Z(_02096__PTR123) );
  MUX2_X1 U6929 ( .A(P1_EAX_PTR28), .B(_02016__PTR28), .S(_02006_), .Z(_02096__PTR124) );
  MUX2_X1 U6930 ( .A(P1_EAX_PTR29), .B(_02016__PTR29), .S(_02006_), .Z(_02096__PTR125) );
  MUX2_X1 U6931 ( .A(P1_EAX_PTR30), .B(_02016__PTR30), .S(_02006_), .Z(_02096__PTR126) );
  MUX2_X1 U6932 ( .A(P1_EAX_PTR31), .B(_02016__PTR31), .S(_02006_), .Z(_02096__PTR127) );
  INV_X1 U6933 ( .A(_01876__PTR21), .ZN(_01876__PTR20) );
  MUX2_X1 U6934 ( .A(_01939__PTR2), .B(1'b0), .S(_01876__PTR21), .Z(_01876__PTR22) );
  INV_X1 U6935 ( .A(_02011_), .ZN(_01939__PTR2) );
  MUX2_X1 U6936 ( .A(_02083__PTR1), .B(1'b0), .S(_02049_), .Z(_01876__PTR16) );
  MUX2_X1 U6937 ( .A(_02083__PTR1), .B(1'b1), .S(_02049_), .Z(_01876__PTR17) );
  MUX2_X1 U6938 ( .A(_02083__PTR2), .B(1'b1), .S(_02049_), .Z(_01876__PTR18) );
  MUX2_X1 U6939 ( .A(na), .B(1'b1), .S(_02060_), .Z(_02083__PTR1) );
  MUX2_X1 U6940 ( .A(_02003_), .B(1'b1), .S(_02060_), .Z(_02083__PTR2) );
  MUX2_X1 U6941 ( .A(_02043__PTR0), .B(1'b0), .S(_01769__PTR4), .Z(_01876__PTR12) );
  MUX2_X1 U6942 ( .A(_02043__PTR1), .B(1'b1), .S(_01769__PTR4), .Z(_01876__PTR13) );
  MUX2_X1 U6943 ( .A(_02043__PTR2), .B(1'b0), .S(_01769__PTR4), .Z(_01876__PTR14) );
  MUX2_X1 U6944 ( .A(_02042__PTR0), .B(1'b0), .S(_02001_), .Z(_02043__PTR0) );
  MUX2_X1 U6945 ( .A(_02042__PTR1), .B(1'b0), .S(_02001_), .Z(_02043__PTR1) );
  MUX2_X1 U6946 ( .A(_02042__PTR2), .B(1'b0), .S(_02001_), .Z(_02043__PTR2) );
  MUX2_X1 U6947 ( .A(_02041__PTR0), .B(1'b1), .S(_02005_), .Z(_02042__PTR0) );
  MUX2_X1 U6948 ( .A(_02041__PTR1), .B(1'b1), .S(_02005_), .Z(_02042__PTR1) );
  MUX2_X1 U6949 ( .A(_02041__PTR2), .B(1'b1), .S(_02005_), .Z(_02042__PTR2) );
  INV_X1 U6950 ( .A(_02008_), .ZN(_02041__PTR0) );
  MUX2_X1 U6951 ( .A(_02040__PTR1), .B(1'b1), .S(_02008_), .Z(_02041__PTR1) );
  MUX2_X1 U6952 ( .A(_02040__PTR2), .B(1'b1), .S(_02008_), .Z(_02041__PTR2) );
  MUX2_X1 U6953 ( .A(_02039__PTR1), .B(1'b0), .S(_02012_), .Z(_02040__PTR1) );
  MUX2_X1 U6954 ( .A(_02021_), .B(1'b0), .S(_02012_), .Z(_02040__PTR2) );
  INV_X1 U6955 ( .A(_02021_), .ZN(_02039__PTR1) );
  INV_X1 U6956 ( .A(P1_CodeFetch), .ZN(_01842__PTR6) );
  INV_X1 U6957 ( .A(P1_ReadRequest), .ZN(_01846__PTR6) );
  INV_X1 U6958 ( .A(P1_RequestPending), .ZN(_01876__PTR4) );
  MUX2_X1 U6959 ( .A(hold), .B(1'b0), .S(P1_RequestPending), .Z(_01876__PTR6) );
  MUX2_X1 U6960 ( .A(1'b0), .B(_02129__PTR0), .S(_01768__PTR2), .Z(_02222__PTR64) );
  MUX2_X1 U6961 ( .A(1'b0), .B(_02129__PTR1), .S(_01768__PTR2), .Z(_02222__PTR65) );
  MUX2_X1 U6962 ( .A(1'b0), .B(_02129__PTR2), .S(_01768__PTR2), .Z(_02222__PTR66) );
  MUX2_X1 U6963 ( .A(1'b0), .B(_02129__PTR3), .S(_01768__PTR2), .Z(_02222__PTR67) );
  MUX2_X1 U6964 ( .A(1'b0), .B(1'b0), .S(_01768__PTR2), .Z(_02222__PTR68) );
  MUX2_X1 U6965 ( .A(1'b0), .B(_02176__PTR3), .S(_01768__PTR2), .Z(_02224__PTR64) );
  MUX2_X1 U6966 ( .A(1'b0), .B(_02176__PTR4), .S(_01768__PTR2), .Z(_02224__PTR65) );
  MUX2_X1 U6967 ( .A(1'b0), .B(_02176__PTR5), .S(_01768__PTR2), .Z(_02224__PTR66) );
  MUX2_X1 U6968 ( .A(1'b0), .B(_02176__PTR6), .S(_01768__PTR2), .Z(_02224__PTR67) );
  MUX2_X1 U6969 ( .A(1'b0), .B(_02371__PTR0), .S(_01768__PTR2), .Z(_02220__PTR64) );
  MUX2_X1 U6970 ( .A(1'b0), .B(_02371__PTR1), .S(_01768__PTR2), .Z(_02220__PTR65) );
  MUX2_X1 U6971 ( .A(1'b0), .B(_02371__PTR2), .S(_01768__PTR2), .Z(_02220__PTR66) );
  MUX2_X1 U6972 ( .A(1'b0), .B(_02371__PTR3), .S(_01768__PTR2), .Z(_02220__PTR67) );
  MUX2_X1 U6973 ( .A(1'b0), .B(_02371__PTR4), .S(_01768__PTR2), .Z(_02220__PTR68) );
  MUX2_X1 U6974 ( .A(1'b0), .B(_02371__PTR5), .S(_01768__PTR2), .Z(_02220__PTR69) );
  MUX2_X1 U6975 ( .A(1'b0), .B(_02371__PTR6), .S(_01768__PTR2), .Z(_02220__PTR70) );
  MUX2_X1 U6976 ( .A(1'b0), .B(_02371__PTR7), .S(_01768__PTR2), .Z(_02220__PTR71) );
  MUX2_X1 U6977 ( .A(1'b0), .B(_02370__PTR0), .S(_01768__PTR2), .Z(_02218__PTR64) );
  MUX2_X1 U6978 ( .A(1'b0), .B(_02370__PTR1), .S(_01768__PTR2), .Z(_02218__PTR65) );
  MUX2_X1 U6979 ( .A(1'b0), .B(_02370__PTR2), .S(_01768__PTR2), .Z(_02218__PTR66) );
  MUX2_X1 U6980 ( .A(1'b0), .B(_02370__PTR3), .S(_01768__PTR2), .Z(_02218__PTR67) );
  MUX2_X1 U6981 ( .A(1'b0), .B(_02370__PTR4), .S(_01768__PTR2), .Z(_02218__PTR68) );
  MUX2_X1 U6982 ( .A(1'b0), .B(_02370__PTR5), .S(_01768__PTR2), .Z(_02218__PTR69) );
  MUX2_X1 U6983 ( .A(1'b0), .B(_02370__PTR6), .S(_01768__PTR2), .Z(_02218__PTR70) );
  MUX2_X1 U6984 ( .A(1'b0), .B(_02370__PTR7), .S(_01768__PTR2), .Z(_02218__PTR71) );
  MUX2_X1 U6985 ( .A(1'b0), .B(_02369__PTR0), .S(_01768__PTR2), .Z(_02216__PTR64) );
  MUX2_X1 U6986 ( .A(1'b0), .B(_02369__PTR1), .S(_01768__PTR2), .Z(_02216__PTR65) );
  MUX2_X1 U6987 ( .A(1'b0), .B(_02369__PTR2), .S(_01768__PTR2), .Z(_02216__PTR66) );
  MUX2_X1 U6988 ( .A(1'b0), .B(_02369__PTR3), .S(_01768__PTR2), .Z(_02216__PTR67) );
  MUX2_X1 U6989 ( .A(1'b0), .B(_02369__PTR4), .S(_01768__PTR2), .Z(_02216__PTR68) );
  MUX2_X1 U6990 ( .A(1'b0), .B(_02369__PTR5), .S(_01768__PTR2), .Z(_02216__PTR69) );
  MUX2_X1 U6991 ( .A(1'b0), .B(_02369__PTR6), .S(_01768__PTR2), .Z(_02216__PTR70) );
  MUX2_X1 U6992 ( .A(1'b0), .B(_02369__PTR7), .S(_01768__PTR2), .Z(_02216__PTR71) );
  MUX2_X1 U6993 ( .A(1'b0), .B(_02368__PTR0), .S(_01768__PTR2), .Z(_02214__PTR64) );
  MUX2_X1 U6994 ( .A(1'b0), .B(_02368__PTR1), .S(_01768__PTR2), .Z(_02214__PTR65) );
  MUX2_X1 U6995 ( .A(1'b0), .B(_02368__PTR2), .S(_01768__PTR2), .Z(_02214__PTR66) );
  MUX2_X1 U6996 ( .A(1'b0), .B(_02368__PTR3), .S(_01768__PTR2), .Z(_02214__PTR67) );
  MUX2_X1 U6997 ( .A(1'b0), .B(_02368__PTR4), .S(_01768__PTR2), .Z(_02214__PTR68) );
  MUX2_X1 U6998 ( .A(1'b0), .B(_02368__PTR5), .S(_01768__PTR2), .Z(_02214__PTR69) );
  MUX2_X1 U6999 ( .A(1'b0), .B(_02368__PTR6), .S(_01768__PTR2), .Z(_02214__PTR70) );
  MUX2_X1 U7000 ( .A(1'b0), .B(_02368__PTR7), .S(_01768__PTR2), .Z(_02214__PTR71) );
  MUX2_X1 U7001 ( .A(1'b0), .B(_02367__PTR0), .S(_01768__PTR2), .Z(_02212__PTR64) );
  MUX2_X1 U7002 ( .A(1'b0), .B(_02367__PTR1), .S(_01768__PTR2), .Z(_02212__PTR65) );
  MUX2_X1 U7003 ( .A(1'b0), .B(_02367__PTR2), .S(_01768__PTR2), .Z(_02212__PTR66) );
  MUX2_X1 U7004 ( .A(1'b0), .B(_02367__PTR3), .S(_01768__PTR2), .Z(_02212__PTR67) );
  MUX2_X1 U7005 ( .A(1'b0), .B(_02367__PTR4), .S(_01768__PTR2), .Z(_02212__PTR68) );
  MUX2_X1 U7006 ( .A(1'b0), .B(_02367__PTR5), .S(_01768__PTR2), .Z(_02212__PTR69) );
  MUX2_X1 U7007 ( .A(1'b0), .B(_02367__PTR6), .S(_01768__PTR2), .Z(_02212__PTR70) );
  MUX2_X1 U7008 ( .A(1'b0), .B(_02367__PTR7), .S(_01768__PTR2), .Z(_02212__PTR71) );
  MUX2_X1 U7009 ( .A(1'b0), .B(_02366__PTR0), .S(_01768__PTR2), .Z(_02210__PTR64) );
  MUX2_X1 U7010 ( .A(1'b0), .B(_02366__PTR1), .S(_01768__PTR2), .Z(_02210__PTR65) );
  MUX2_X1 U7011 ( .A(1'b0), .B(_02366__PTR2), .S(_01768__PTR2), .Z(_02210__PTR66) );
  MUX2_X1 U7012 ( .A(1'b0), .B(_02366__PTR3), .S(_01768__PTR2), .Z(_02210__PTR67) );
  MUX2_X1 U7013 ( .A(1'b0), .B(_02366__PTR4), .S(_01768__PTR2), .Z(_02210__PTR68) );
  MUX2_X1 U7014 ( .A(1'b0), .B(_02366__PTR5), .S(_01768__PTR2), .Z(_02210__PTR69) );
  MUX2_X1 U7015 ( .A(1'b0), .B(_02366__PTR6), .S(_01768__PTR2), .Z(_02210__PTR70) );
  MUX2_X1 U7016 ( .A(1'b0), .B(_02366__PTR7), .S(_01768__PTR2), .Z(_02210__PTR71) );
  MUX2_X1 U7017 ( .A(1'b0), .B(_02365__PTR0), .S(_01768__PTR2), .Z(_02208__PTR64) );
  MUX2_X1 U7018 ( .A(1'b0), .B(_02365__PTR1), .S(_01768__PTR2), .Z(_02208__PTR65) );
  MUX2_X1 U7019 ( .A(1'b0), .B(_02365__PTR2), .S(_01768__PTR2), .Z(_02208__PTR66) );
  MUX2_X1 U7020 ( .A(1'b0), .B(_02365__PTR3), .S(_01768__PTR2), .Z(_02208__PTR67) );
  MUX2_X1 U7021 ( .A(1'b0), .B(_02365__PTR4), .S(_01768__PTR2), .Z(_02208__PTR68) );
  MUX2_X1 U7022 ( .A(1'b0), .B(_02365__PTR5), .S(_01768__PTR2), .Z(_02208__PTR69) );
  MUX2_X1 U7023 ( .A(1'b0), .B(_02365__PTR6), .S(_01768__PTR2), .Z(_02208__PTR70) );
  MUX2_X1 U7024 ( .A(1'b0), .B(_02365__PTR7), .S(_01768__PTR2), .Z(_02208__PTR71) );
  MUX2_X1 U7025 ( .A(1'b0), .B(_02364__PTR0), .S(_01768__PTR2), .Z(_02206__PTR64) );
  MUX2_X1 U7026 ( .A(1'b0), .B(_02364__PTR1), .S(_01768__PTR2), .Z(_02206__PTR65) );
  MUX2_X1 U7027 ( .A(1'b0), .B(_02364__PTR2), .S(_01768__PTR2), .Z(_02206__PTR66) );
  MUX2_X1 U7028 ( .A(1'b0), .B(_02364__PTR3), .S(_01768__PTR2), .Z(_02206__PTR67) );
  MUX2_X1 U7029 ( .A(1'b0), .B(_02364__PTR4), .S(_01768__PTR2), .Z(_02206__PTR68) );
  MUX2_X1 U7030 ( .A(1'b0), .B(_02364__PTR5), .S(_01768__PTR2), .Z(_02206__PTR69) );
  MUX2_X1 U7031 ( .A(1'b0), .B(_02364__PTR6), .S(_01768__PTR2), .Z(_02206__PTR70) );
  MUX2_X1 U7032 ( .A(1'b0), .B(_02364__PTR7), .S(_01768__PTR2), .Z(_02206__PTR71) );
  MUX2_X1 U7033 ( .A(1'b0), .B(_02363__PTR0), .S(_01768__PTR2), .Z(_02204__PTR64) );
  MUX2_X1 U7034 ( .A(1'b0), .B(_02363__PTR1), .S(_01768__PTR2), .Z(_02204__PTR65) );
  MUX2_X1 U7035 ( .A(1'b0), .B(_02363__PTR2), .S(_01768__PTR2), .Z(_02204__PTR66) );
  MUX2_X1 U7036 ( .A(1'b0), .B(_02363__PTR3), .S(_01768__PTR2), .Z(_02204__PTR67) );
  MUX2_X1 U7037 ( .A(1'b0), .B(_02363__PTR4), .S(_01768__PTR2), .Z(_02204__PTR68) );
  MUX2_X1 U7038 ( .A(1'b0), .B(_02363__PTR5), .S(_01768__PTR2), .Z(_02204__PTR69) );
  MUX2_X1 U7039 ( .A(1'b0), .B(_02363__PTR6), .S(_01768__PTR2), .Z(_02204__PTR70) );
  MUX2_X1 U7040 ( .A(1'b0), .B(_02363__PTR7), .S(_01768__PTR2), .Z(_02204__PTR71) );
  MUX2_X1 U7041 ( .A(1'b0), .B(_02362__PTR0), .S(_01768__PTR2), .Z(_02202__PTR64) );
  MUX2_X1 U7042 ( .A(1'b0), .B(_02362__PTR1), .S(_01768__PTR2), .Z(_02202__PTR65) );
  MUX2_X1 U7043 ( .A(1'b0), .B(_02362__PTR2), .S(_01768__PTR2), .Z(_02202__PTR66) );
  MUX2_X1 U7044 ( .A(1'b0), .B(_02362__PTR3), .S(_01768__PTR2), .Z(_02202__PTR67) );
  MUX2_X1 U7045 ( .A(1'b0), .B(_02362__PTR4), .S(_01768__PTR2), .Z(_02202__PTR68) );
  MUX2_X1 U7046 ( .A(1'b0), .B(_02362__PTR5), .S(_01768__PTR2), .Z(_02202__PTR69) );
  MUX2_X1 U7047 ( .A(1'b0), .B(_02362__PTR6), .S(_01768__PTR2), .Z(_02202__PTR70) );
  MUX2_X1 U7048 ( .A(1'b0), .B(_02362__PTR7), .S(_01768__PTR2), .Z(_02202__PTR71) );
  MUX2_X1 U7049 ( .A(1'b0), .B(_02361__PTR0), .S(_01768__PTR2), .Z(_02200__PTR64) );
  MUX2_X1 U7050 ( .A(1'b0), .B(_02361__PTR1), .S(_01768__PTR2), .Z(_02200__PTR65) );
  MUX2_X1 U7051 ( .A(1'b0), .B(_02361__PTR2), .S(_01768__PTR2), .Z(_02200__PTR66) );
  MUX2_X1 U7052 ( .A(1'b0), .B(_02361__PTR3), .S(_01768__PTR2), .Z(_02200__PTR67) );
  MUX2_X1 U7053 ( .A(1'b0), .B(_02361__PTR4), .S(_01768__PTR2), .Z(_02200__PTR68) );
  MUX2_X1 U7054 ( .A(1'b0), .B(_02361__PTR5), .S(_01768__PTR2), .Z(_02200__PTR69) );
  MUX2_X1 U7055 ( .A(1'b0), .B(_02361__PTR6), .S(_01768__PTR2), .Z(_02200__PTR70) );
  MUX2_X1 U7056 ( .A(1'b0), .B(_02361__PTR7), .S(_01768__PTR2), .Z(_02200__PTR71) );
  MUX2_X1 U7057 ( .A(1'b0), .B(_02360__PTR0), .S(_01768__PTR2), .Z(_02198__PTR64) );
  MUX2_X1 U7058 ( .A(1'b0), .B(_02360__PTR1), .S(_01768__PTR2), .Z(_02198__PTR65) );
  MUX2_X1 U7059 ( .A(1'b0), .B(_02360__PTR2), .S(_01768__PTR2), .Z(_02198__PTR66) );
  MUX2_X1 U7060 ( .A(1'b0), .B(_02360__PTR3), .S(_01768__PTR2), .Z(_02198__PTR67) );
  MUX2_X1 U7061 ( .A(1'b0), .B(_02360__PTR4), .S(_01768__PTR2), .Z(_02198__PTR68) );
  MUX2_X1 U7062 ( .A(1'b0), .B(_02360__PTR5), .S(_01768__PTR2), .Z(_02198__PTR69) );
  MUX2_X1 U7063 ( .A(1'b0), .B(_02360__PTR6), .S(_01768__PTR2), .Z(_02198__PTR70) );
  MUX2_X1 U7064 ( .A(1'b0), .B(_02360__PTR7), .S(_01768__PTR2), .Z(_02198__PTR71) );
  MUX2_X1 U7065 ( .A(1'b0), .B(_02359__PTR0), .S(_01768__PTR2), .Z(_02196__PTR64) );
  MUX2_X1 U7066 ( .A(1'b0), .B(_02359__PTR1), .S(_01768__PTR2), .Z(_02196__PTR65) );
  MUX2_X1 U7067 ( .A(1'b0), .B(_02359__PTR2), .S(_01768__PTR2), .Z(_02196__PTR66) );
  MUX2_X1 U7068 ( .A(1'b0), .B(_02359__PTR3), .S(_01768__PTR2), .Z(_02196__PTR67) );
  MUX2_X1 U7069 ( .A(1'b0), .B(_02359__PTR4), .S(_01768__PTR2), .Z(_02196__PTR68) );
  MUX2_X1 U7070 ( .A(1'b0), .B(_02359__PTR5), .S(_01768__PTR2), .Z(_02196__PTR69) );
  MUX2_X1 U7071 ( .A(1'b0), .B(_02359__PTR6), .S(_01768__PTR2), .Z(_02196__PTR70) );
  MUX2_X1 U7072 ( .A(1'b0), .B(_02359__PTR7), .S(_01768__PTR2), .Z(_02196__PTR71) );
  MUX2_X1 U7073 ( .A(1'b0), .B(_02358__PTR0), .S(_01768__PTR2), .Z(_02194__PTR64) );
  MUX2_X1 U7074 ( .A(1'b0), .B(_02358__PTR1), .S(_01768__PTR2), .Z(_02194__PTR65) );
  MUX2_X1 U7075 ( .A(1'b0), .B(_02358__PTR2), .S(_01768__PTR2), .Z(_02194__PTR66) );
  MUX2_X1 U7076 ( .A(1'b0), .B(_02358__PTR3), .S(_01768__PTR2), .Z(_02194__PTR67) );
  MUX2_X1 U7077 ( .A(1'b0), .B(_02358__PTR4), .S(_01768__PTR2), .Z(_02194__PTR68) );
  MUX2_X1 U7078 ( .A(1'b0), .B(_02358__PTR5), .S(_01768__PTR2), .Z(_02194__PTR69) );
  MUX2_X1 U7079 ( .A(1'b0), .B(_02358__PTR6), .S(_01768__PTR2), .Z(_02194__PTR70) );
  MUX2_X1 U7080 ( .A(1'b0), .B(_02358__PTR7), .S(_01768__PTR2), .Z(_02194__PTR71) );
  MUX2_X1 U7081 ( .A(1'b0), .B(_02357__PTR0), .S(_01768__PTR2), .Z(_02192__PTR64) );
  MUX2_X1 U7082 ( .A(1'b0), .B(_02357__PTR1), .S(_01768__PTR2), .Z(_02192__PTR65) );
  MUX2_X1 U7083 ( .A(1'b0), .B(_02357__PTR2), .S(_01768__PTR2), .Z(_02192__PTR66) );
  MUX2_X1 U7084 ( .A(1'b0), .B(_02357__PTR3), .S(_01768__PTR2), .Z(_02192__PTR67) );
  MUX2_X1 U7085 ( .A(1'b0), .B(_02357__PTR4), .S(_01768__PTR2), .Z(_02192__PTR68) );
  MUX2_X1 U7086 ( .A(1'b0), .B(_02357__PTR5), .S(_01768__PTR2), .Z(_02192__PTR69) );
  MUX2_X1 U7087 ( .A(1'b0), .B(_02357__PTR6), .S(_01768__PTR2), .Z(_02192__PTR70) );
  MUX2_X1 U7088 ( .A(1'b0), .B(_02357__PTR7), .S(_01768__PTR2), .Z(_02192__PTR71) );
  MUX2_X1 U7089 ( .A(1'b0), .B(_02356__PTR0), .S(_01768__PTR2), .Z(_02190__PTR64) );
  MUX2_X1 U7090 ( .A(1'b0), .B(_02356__PTR1), .S(_01768__PTR2), .Z(_02190__PTR65) );
  MUX2_X1 U7091 ( .A(1'b0), .B(_02356__PTR2), .S(_01768__PTR2), .Z(_02190__PTR66) );
  MUX2_X1 U7092 ( .A(1'b0), .B(_02356__PTR3), .S(_01768__PTR2), .Z(_02190__PTR67) );
  MUX2_X1 U7093 ( .A(1'b0), .B(_02356__PTR4), .S(_01768__PTR2), .Z(_02190__PTR68) );
  MUX2_X1 U7094 ( .A(1'b0), .B(_02356__PTR5), .S(_01768__PTR2), .Z(_02190__PTR69) );
  MUX2_X1 U7095 ( .A(1'b0), .B(_02356__PTR6), .S(_01768__PTR2), .Z(_02190__PTR70) );
  MUX2_X1 U7096 ( .A(1'b0), .B(_02356__PTR7), .S(_01768__PTR2), .Z(_02190__PTR71) );
  MUX2_X1 U7097 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR0), .Z(_02371__PTR0) );
  MUX2_X1 U7098 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR0), .Z(_02371__PTR1) );
  MUX2_X1 U7099 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR0), .Z(_02371__PTR2) );
  MUX2_X1 U7100 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR0), .Z(_02371__PTR3) );
  MUX2_X1 U7101 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR0), .Z(_02371__PTR4) );
  MUX2_X1 U7102 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR0), .Z(_02371__PTR5) );
  MUX2_X1 U7103 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR0), .Z(_02371__PTR6) );
  MUX2_X1 U7104 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR0), .Z(_02371__PTR7) );
  MUX2_X1 U7105 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR1), .Z(_02370__PTR0) );
  MUX2_X1 U7106 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR1), .Z(_02370__PTR1) );
  MUX2_X1 U7107 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR1), .Z(_02370__PTR2) );
  MUX2_X1 U7108 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR1), .Z(_02370__PTR3) );
  MUX2_X1 U7109 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR1), .Z(_02370__PTR4) );
  MUX2_X1 U7110 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR1), .Z(_02370__PTR5) );
  MUX2_X1 U7111 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR1), .Z(_02370__PTR6) );
  MUX2_X1 U7112 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR1), .Z(_02370__PTR7) );
  MUX2_X1 U7113 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR2), .Z(_02369__PTR0) );
  MUX2_X1 U7114 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR2), .Z(_02369__PTR1) );
  MUX2_X1 U7115 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR2), .Z(_02369__PTR2) );
  MUX2_X1 U7116 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR2), .Z(_02369__PTR3) );
  MUX2_X1 U7117 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR2), .Z(_02369__PTR4) );
  MUX2_X1 U7118 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR2), .Z(_02369__PTR5) );
  MUX2_X1 U7119 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR2), .Z(_02369__PTR6) );
  MUX2_X1 U7120 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR2), .Z(_02369__PTR7) );
  MUX2_X1 U7121 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR3), .Z(_02368__PTR0) );
  MUX2_X1 U7122 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR3), .Z(_02368__PTR1) );
  MUX2_X1 U7123 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR3), .Z(_02368__PTR2) );
  MUX2_X1 U7124 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR3), .Z(_02368__PTR3) );
  MUX2_X1 U7125 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR3), .Z(_02368__PTR4) );
  MUX2_X1 U7126 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR3), .Z(_02368__PTR5) );
  MUX2_X1 U7127 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR3), .Z(_02368__PTR6) );
  MUX2_X1 U7128 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR3), .Z(_02368__PTR7) );
  MUX2_X1 U7129 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR4), .Z(_02367__PTR0) );
  MUX2_X1 U7130 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR4), .Z(_02367__PTR1) );
  MUX2_X1 U7131 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR4), .Z(_02367__PTR2) );
  MUX2_X1 U7132 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR4), .Z(_02367__PTR3) );
  MUX2_X1 U7133 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR4), .Z(_02367__PTR4) );
  MUX2_X1 U7134 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR4), .Z(_02367__PTR5) );
  MUX2_X1 U7135 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR4), .Z(_02367__PTR6) );
  MUX2_X1 U7136 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR4), .Z(_02367__PTR7) );
  MUX2_X1 U7137 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR5), .Z(_02366__PTR0) );
  MUX2_X1 U7138 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR5), .Z(_02366__PTR1) );
  MUX2_X1 U7139 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR5), .Z(_02366__PTR2) );
  MUX2_X1 U7140 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR5), .Z(_02366__PTR3) );
  MUX2_X1 U7141 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR5), .Z(_02366__PTR4) );
  MUX2_X1 U7142 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR5), .Z(_02366__PTR5) );
  MUX2_X1 U7143 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR5), .Z(_02366__PTR6) );
  MUX2_X1 U7144 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR5), .Z(_02366__PTR7) );
  MUX2_X1 U7145 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR6), .Z(_02365__PTR0) );
  MUX2_X1 U7146 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR6), .Z(_02365__PTR1) );
  MUX2_X1 U7147 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR6), .Z(_02365__PTR2) );
  MUX2_X1 U7148 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR6), .Z(_02365__PTR3) );
  MUX2_X1 U7149 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR6), .Z(_02365__PTR4) );
  MUX2_X1 U7150 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR6), .Z(_02365__PTR5) );
  MUX2_X1 U7151 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR6), .Z(_02365__PTR6) );
  MUX2_X1 U7152 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR6), .Z(_02365__PTR7) );
  MUX2_X1 U7153 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR7), .Z(_02364__PTR0) );
  MUX2_X1 U7154 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR7), .Z(_02364__PTR1) );
  MUX2_X1 U7155 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR7), .Z(_02364__PTR2) );
  MUX2_X1 U7156 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR7), .Z(_02364__PTR3) );
  MUX2_X1 U7157 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR7), .Z(_02364__PTR4) );
  MUX2_X1 U7158 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR7), .Z(_02364__PTR5) );
  MUX2_X1 U7159 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR7), .Z(_02364__PTR6) );
  MUX2_X1 U7160 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR7), .Z(_02364__PTR7) );
  MUX2_X1 U7161 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR8), .Z(_02363__PTR0) );
  MUX2_X1 U7162 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR8), .Z(_02363__PTR1) );
  MUX2_X1 U7163 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR8), .Z(_02363__PTR2) );
  MUX2_X1 U7164 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR8), .Z(_02363__PTR3) );
  MUX2_X1 U7165 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR8), .Z(_02363__PTR4) );
  MUX2_X1 U7166 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR8), .Z(_02363__PTR5) );
  MUX2_X1 U7167 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR8), .Z(_02363__PTR6) );
  MUX2_X1 U7168 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR8), .Z(_02363__PTR7) );
  MUX2_X1 U7169 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR9), .Z(_02362__PTR0) );
  MUX2_X1 U7170 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR9), .Z(_02362__PTR1) );
  MUX2_X1 U7171 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR9), .Z(_02362__PTR2) );
  MUX2_X1 U7172 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR9), .Z(_02362__PTR3) );
  MUX2_X1 U7173 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR9), .Z(_02362__PTR4) );
  MUX2_X1 U7174 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR9), .Z(_02362__PTR5) );
  MUX2_X1 U7175 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR9), .Z(_02362__PTR6) );
  MUX2_X1 U7176 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR9), .Z(_02362__PTR7) );
  MUX2_X1 U7177 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR10), .Z(_02361__PTR0) );
  MUX2_X1 U7178 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR10), .Z(_02361__PTR1) );
  MUX2_X1 U7179 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR10), .Z(_02361__PTR2) );
  MUX2_X1 U7180 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR10), .Z(_02361__PTR3) );
  MUX2_X1 U7181 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR10), .Z(_02361__PTR4) );
  MUX2_X1 U7182 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR10), .Z(_02361__PTR5) );
  MUX2_X1 U7183 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR10), .Z(_02361__PTR6) );
  MUX2_X1 U7184 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR10), .Z(_02361__PTR7) );
  MUX2_X1 U7185 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR11), .Z(_02360__PTR0) );
  MUX2_X1 U7186 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR11), .Z(_02360__PTR1) );
  MUX2_X1 U7187 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR11), .Z(_02360__PTR2) );
  MUX2_X1 U7188 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR11), .Z(_02360__PTR3) );
  MUX2_X1 U7189 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR11), .Z(_02360__PTR4) );
  MUX2_X1 U7190 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR11), .Z(_02360__PTR5) );
  MUX2_X1 U7191 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR11), .Z(_02360__PTR6) );
  MUX2_X1 U7192 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR11), .Z(_02360__PTR7) );
  MUX2_X1 U7193 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR12), .Z(_02359__PTR0) );
  MUX2_X1 U7194 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR12), .Z(_02359__PTR1) );
  MUX2_X1 U7195 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR12), .Z(_02359__PTR2) );
  MUX2_X1 U7196 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR12), .Z(_02359__PTR3) );
  MUX2_X1 U7197 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR12), .Z(_02359__PTR4) );
  MUX2_X1 U7198 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR12), .Z(_02359__PTR5) );
  MUX2_X1 U7199 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR12), .Z(_02359__PTR6) );
  MUX2_X1 U7200 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR12), .Z(_02359__PTR7) );
  MUX2_X1 U7201 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR13), .Z(_02358__PTR0) );
  MUX2_X1 U7202 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR13), .Z(_02358__PTR1) );
  MUX2_X1 U7203 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR13), .Z(_02358__PTR2) );
  MUX2_X1 U7204 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR13), .Z(_02358__PTR3) );
  MUX2_X1 U7205 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR13), .Z(_02358__PTR4) );
  MUX2_X1 U7206 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR13), .Z(_02358__PTR5) );
  MUX2_X1 U7207 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR13), .Z(_02358__PTR6) );
  MUX2_X1 U7208 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR13), .Z(_02358__PTR7) );
  MUX2_X1 U7209 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR14), .Z(_02357__PTR0) );
  MUX2_X1 U7210 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR14), .Z(_02357__PTR1) );
  MUX2_X1 U7211 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR14), .Z(_02357__PTR2) );
  MUX2_X1 U7212 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR14), .Z(_02357__PTR3) );
  MUX2_X1 U7213 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR14), .Z(_02357__PTR4) );
  MUX2_X1 U7214 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR14), .Z(_02357__PTR5) );
  MUX2_X1 U7215 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR14), .Z(_02357__PTR6) );
  MUX2_X1 U7216 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR14), .Z(_02357__PTR7) );
  MUX2_X1 U7217 ( .A(1'b0), .B(_02175__PTR0), .S(_02128__PTR15), .Z(_02356__PTR0) );
  MUX2_X1 U7218 ( .A(1'b0), .B(_02175__PTR1), .S(_02128__PTR15), .Z(_02356__PTR1) );
  MUX2_X1 U7219 ( .A(1'b0), .B(_02175__PTR2), .S(_02128__PTR15), .Z(_02356__PTR2) );
  MUX2_X1 U7220 ( .A(1'b0), .B(_02175__PTR3), .S(_02128__PTR15), .Z(_02356__PTR3) );
  MUX2_X1 U7221 ( .A(1'b0), .B(_02175__PTR4), .S(_02128__PTR15), .Z(_02356__PTR4) );
  MUX2_X1 U7222 ( .A(1'b0), .B(_02175__PTR5), .S(_02128__PTR15), .Z(_02356__PTR5) );
  MUX2_X1 U7223 ( .A(1'b0), .B(_02175__PTR6), .S(_02128__PTR15), .Z(_02356__PTR6) );
  MUX2_X1 U7224 ( .A(1'b0), .B(_02175__PTR7), .S(_02128__PTR15), .Z(_02356__PTR7) );
  MUX2_X1 U7225 ( .A(1'b0), .B(_02355__PTR0), .S(_02186__PTR28), .Z(_02222__PTR56) );
  MUX2_X1 U7226 ( .A(1'b0), .B(_02355__PTR4), .S(_02186__PTR28), .Z(_02222__PTR60) );
  MUX2_X1 U7227 ( .A(1'b0), .B(1'b1), .S(P2_P1_Flush), .Z(_02355__PTR0) );
  MUX2_X1 U7228 ( .A(1'b0), .B(1'b0), .S(P2_P1_Flush), .Z(_02355__PTR4) );
  MUX2_X1 U7229 ( .A(P2_P1_InstQueueRd_Addr_PTR0), .B(_02354__PTR0), .S(P2_P1_Flush), .Z(_02224__PTR56) );
  MUX2_X1 U7230 ( .A(P2_P1_InstQueueRd_Addr_PTR1), .B(_02354__PTR1), .S(P2_P1_Flush), .Z(_02224__PTR57) );
  MUX2_X1 U7231 ( .A(P2_P1_InstQueueRd_Addr_PTR2), .B(_02354__PTR2), .S(P2_P1_Flush), .Z(_02224__PTR58) );
  MUX2_X1 U7232 ( .A(P2_P1_InstQueueRd_Addr_PTR3), .B(1'b0), .S(P2_P1_Flush), .Z(_02224__PTR59) );
  MUX2_X1 U7233 ( .A(P2_P1_InstQueueRd_Addr_PTR4), .B(1'b0), .S(P2_P1_Flush), .Z(_02224__PTR60) );
  MUX2_X1 U7234 ( .A(1'b1), .B(_02373__PTR0), .S(P2_P1_InstAddrPointer_PTR0), .Z(_02354__PTR0) );
  MUX2_X1 U7235 ( .A(1'b0), .B(_03076__PTR1), .S(P2_P1_InstAddrPointer_PTR0), .Z(_02354__PTR1) );
  MUX2_X1 U7236 ( .A(1'b0), .B(_03075__PTR1), .S(P2_P1_InstAddrPointer_PTR0), .Z(_02354__PTR2) );
  MUX2_X1 U7237 ( .A(_03194__PTR1), .B(P2_P1_InstAddrPointer_PTR1), .S(_02989__PTR31), .Z(_03074__PTR1) );
  MUX2_X1 U7238 ( .A(1'b1), .B(1'b0), .S(P2_READY_n), .Z(_02186__PTR26) );
  MUX2_X1 U7239 ( .A(1'b0), .B(1'b0), .S(P2_READY_n), .Z(_02142__PTR6) );
  MUX2_X1 U7240 ( .A(_02410__PTR0), .B(1'b1), .S(_02353_), .Z(_02186__PTR20) );
  MUX2_X1 U7241 ( .A(_02410__PTR1), .B(1'b1), .S(_02353_), .Z(_02186__PTR21) );
  MUX2_X1 U7242 ( .A(_02410__PTR2), .B(1'b1), .S(_02353_), .Z(_02186__PTR22) );
  MUX2_X1 U7243 ( .A(_02410__PTR3), .B(1'b0), .S(_02353_), .Z(_02186__PTR23) );
  MUX2_X1 U7244 ( .A(P2_Datao_PTR16), .B(_02336__PTR16), .S(_02296_), .Z(_02403__PTR48) );
  MUX2_X1 U7245 ( .A(P2_Datao_PTR17), .B(_02336__PTR17), .S(_02296_), .Z(_02403__PTR49) );
  MUX2_X1 U7246 ( .A(P2_Datao_PTR18), .B(_02336__PTR18), .S(_02296_), .Z(_02403__PTR50) );
  MUX2_X1 U7247 ( .A(P2_Datao_PTR19), .B(_02336__PTR19), .S(_02296_), .Z(_02403__PTR51) );
  MUX2_X1 U7248 ( .A(P2_Datao_PTR20), .B(_02336__PTR20), .S(_02296_), .Z(_02403__PTR52) );
  MUX2_X1 U7249 ( .A(P2_Datao_PTR21), .B(_02336__PTR21), .S(_02296_), .Z(_02403__PTR53) );
  MUX2_X1 U7250 ( .A(P2_Datao_PTR22), .B(_02336__PTR22), .S(_02296_), .Z(_02403__PTR54) );
  MUX2_X1 U7251 ( .A(P2_Datao_PTR23), .B(_02336__PTR23), .S(_02296_), .Z(_02403__PTR55) );
  MUX2_X1 U7252 ( .A(P2_Datao_PTR24), .B(_02336__PTR24), .S(_02296_), .Z(_02403__PTR56) );
  MUX2_X1 U7253 ( .A(P2_Datao_PTR25), .B(_02336__PTR25), .S(_02296_), .Z(_02403__PTR57) );
  MUX2_X1 U7254 ( .A(P2_Datao_PTR26), .B(_02336__PTR26), .S(_02296_), .Z(_02403__PTR58) );
  MUX2_X1 U7255 ( .A(P2_Datao_PTR27), .B(_02336__PTR27), .S(_02296_), .Z(_02403__PTR59) );
  MUX2_X1 U7256 ( .A(P2_Datao_PTR28), .B(_02336__PTR28), .S(_02296_), .Z(_02403__PTR60) );
  MUX2_X1 U7257 ( .A(P2_Datao_PTR29), .B(_02336__PTR29), .S(_02296_), .Z(_02403__PTR61) );
  MUX2_X1 U7258 ( .A(P2_Datao_PTR30), .B(_02336__PTR30), .S(_02296_), .Z(_02403__PTR62) );
  MUX2_X1 U7259 ( .A(P2_Datao_PTR31), .B(_02321__PTR31), .S(_02296_), .Z(_02403__PTR95) );
  MUX2_X1 U7260 ( .A(P2_Datao_PTR0), .B(_02321__PTR0), .S(_02296_), .Z(_02403__PTR64) );
  MUX2_X1 U7261 ( .A(P2_Datao_PTR1), .B(_02321__PTR1), .S(_02296_), .Z(_02403__PTR65) );
  MUX2_X1 U7262 ( .A(P2_Datao_PTR2), .B(_02321__PTR2), .S(_02296_), .Z(_02403__PTR66) );
  MUX2_X1 U7263 ( .A(P2_Datao_PTR3), .B(_02321__PTR3), .S(_02296_), .Z(_02403__PTR67) );
  MUX2_X1 U7264 ( .A(P2_Datao_PTR4), .B(_02321__PTR4), .S(_02296_), .Z(_02403__PTR68) );
  MUX2_X1 U7265 ( .A(P2_Datao_PTR5), .B(_02321__PTR5), .S(_02296_), .Z(_02403__PTR69) );
  MUX2_X1 U7266 ( .A(P2_Datao_PTR6), .B(_02321__PTR6), .S(_02296_), .Z(_02403__PTR70) );
  MUX2_X1 U7267 ( .A(P2_Datao_PTR7), .B(_02321__PTR7), .S(_02296_), .Z(_02403__PTR71) );
  MUX2_X1 U7268 ( .A(P2_Datao_PTR8), .B(_02321__PTR8), .S(_02296_), .Z(_02403__PTR72) );
  MUX2_X1 U7269 ( .A(P2_Datao_PTR9), .B(_02321__PTR9), .S(_02296_), .Z(_02403__PTR73) );
  MUX2_X1 U7270 ( .A(P2_Datao_PTR10), .B(_02321__PTR10), .S(_02296_), .Z(_02403__PTR74) );
  MUX2_X1 U7271 ( .A(P2_Datao_PTR11), .B(_02321__PTR11), .S(_02296_), .Z(_02403__PTR75) );
  MUX2_X1 U7272 ( .A(P2_Datao_PTR12), .B(_02321__PTR12), .S(_02296_), .Z(_02403__PTR76) );
  MUX2_X1 U7273 ( .A(P2_Datao_PTR13), .B(_02321__PTR13), .S(_02296_), .Z(_02403__PTR77) );
  MUX2_X1 U7274 ( .A(P2_Datao_PTR14), .B(_02321__PTR14), .S(_02296_), .Z(_02403__PTR78) );
  MUX2_X1 U7275 ( .A(P2_Datao_PTR15), .B(_02321__PTR15), .S(_02296_), .Z(_02403__PTR79) );
  MUX2_X1 U7276 ( .A(P2_Datao_PTR16), .B(_02321__PTR16), .S(_02296_), .Z(_02403__PTR80) );
  MUX2_X1 U7277 ( .A(P2_Datao_PTR17), .B(_02321__PTR17), .S(_02296_), .Z(_02403__PTR81) );
  MUX2_X1 U7278 ( .A(P2_Datao_PTR18), .B(_02321__PTR18), .S(_02296_), .Z(_02403__PTR82) );
  MUX2_X1 U7279 ( .A(P2_Datao_PTR19), .B(_02321__PTR19), .S(_02296_), .Z(_02403__PTR83) );
  MUX2_X1 U7280 ( .A(P2_Datao_PTR20), .B(_02321__PTR20), .S(_02296_), .Z(_02403__PTR84) );
  MUX2_X1 U7281 ( .A(P2_Datao_PTR21), .B(_02321__PTR21), .S(_02296_), .Z(_02403__PTR85) );
  MUX2_X1 U7282 ( .A(P2_Datao_PTR22), .B(_02321__PTR22), .S(_02296_), .Z(_02403__PTR86) );
  MUX2_X1 U7283 ( .A(P2_Datao_PTR23), .B(_02321__PTR23), .S(_02296_), .Z(_02403__PTR87) );
  MUX2_X1 U7284 ( .A(P2_Datao_PTR24), .B(_02321__PTR24), .S(_02296_), .Z(_02403__PTR88) );
  MUX2_X1 U7285 ( .A(P2_Datao_PTR25), .B(_02321__PTR25), .S(_02296_), .Z(_02403__PTR89) );
  MUX2_X1 U7286 ( .A(P2_Datao_PTR26), .B(_02321__PTR26), .S(_02296_), .Z(_02403__PTR90) );
  MUX2_X1 U7287 ( .A(P2_Datao_PTR27), .B(_02321__PTR27), .S(_02296_), .Z(_02403__PTR91) );
  MUX2_X1 U7288 ( .A(P2_Datao_PTR28), .B(_02321__PTR28), .S(_02296_), .Z(_02403__PTR92) );
  MUX2_X1 U7289 ( .A(P2_Datao_PTR29), .B(_02321__PTR29), .S(_02296_), .Z(_02403__PTR93) );
  MUX2_X1 U7290 ( .A(P2_Datao_PTR30), .B(_02321__PTR30), .S(_02296_), .Z(_02403__PTR94) );
  MUX2_X1 U7291 ( .A(P2_RequestPending), .B(_02337_), .S(_02296_), .Z(_02154__PTR0) );
  MUX2_X1 U7292 ( .A(1'b1), .B(P2_READY_n), .S(_02315_), .Z(_02337_) );
  MUX2_X1 U7293 ( .A(P2_MemoryFetch), .B(1'b0), .S(_02296_), .Z(_02161__PTR0) );
  MUX2_X1 U7294 ( .A(1'b0), .B(_02326_), .S(_02296_), .Z(_02146__PTR0) );
  MUX2_X1 U7295 ( .A(1'b1), .B(_02325_), .S(_02296_), .Z(_02150__PTR0) );
  MUX2_X1 U7296 ( .A(P2_P1_State2_PTR0), .B(_02324__PTR0), .S(_02296_), .Z(_02407__PTR4) );
  MUX2_X1 U7297 ( .A(P2_P1_State2_PTR1), .B(_02324__PTR1), .S(_02296_), .Z(_02407__PTR5) );
  MUX2_X1 U7298 ( .A(P2_P1_State2_PTR2), .B(_02324__PTR2), .S(_02296_), .Z(_02407__PTR6) );
  MUX2_X1 U7299 ( .A(P2_P1_State2_PTR3), .B(_02324__PTR3), .S(_02296_), .Z(_02407__PTR7) );
  MUX2_X1 U7300 ( .A(P2_Datao_PTR16), .B(1'b0), .S(_02315_), .Z(_02336__PTR16) );
  MUX2_X1 U7301 ( .A(P2_Datao_PTR17), .B(1'b0), .S(_02315_), .Z(_02336__PTR17) );
  MUX2_X1 U7302 ( .A(P2_Datao_PTR18), .B(1'b0), .S(_02315_), .Z(_02336__PTR18) );
  MUX2_X1 U7303 ( .A(P2_Datao_PTR19), .B(1'b0), .S(_02315_), .Z(_02336__PTR19) );
  MUX2_X1 U7304 ( .A(P2_Datao_PTR20), .B(1'b0), .S(_02315_), .Z(_02336__PTR20) );
  MUX2_X1 U7305 ( .A(P2_Datao_PTR21), .B(1'b0), .S(_02315_), .Z(_02336__PTR21) );
  MUX2_X1 U7306 ( .A(P2_Datao_PTR22), .B(1'b0), .S(_02315_), .Z(_02336__PTR22) );
  MUX2_X1 U7307 ( .A(P2_Datao_PTR23), .B(1'b0), .S(_02315_), .Z(_02336__PTR23) );
  MUX2_X1 U7308 ( .A(P2_Datao_PTR24), .B(1'b0), .S(_02315_), .Z(_02336__PTR24) );
  MUX2_X1 U7309 ( .A(P2_Datao_PTR25), .B(1'b0), .S(_02315_), .Z(_02336__PTR25) );
  MUX2_X1 U7310 ( .A(P2_Datao_PTR26), .B(1'b0), .S(_02315_), .Z(_02336__PTR26) );
  MUX2_X1 U7311 ( .A(P2_Datao_PTR27), .B(1'b0), .S(_02315_), .Z(_02336__PTR27) );
  MUX2_X1 U7312 ( .A(P2_Datao_PTR28), .B(1'b0), .S(_02315_), .Z(_02336__PTR28) );
  MUX2_X1 U7313 ( .A(P2_Datao_PTR29), .B(1'b0), .S(_02315_), .Z(_02336__PTR29) );
  MUX2_X1 U7314 ( .A(P2_Datao_PTR30), .B(1'b0), .S(_02315_), .Z(_02336__PTR30) );
  MUX2_X1 U7315 ( .A(P2_Datao_PTR31), .B(1'b0), .S(_02315_), .Z(_02321__PTR31) );
  MUX2_X1 U7316 ( .A(P2_Datao_PTR0), .B(P2_EAX_PTR0), .S(_02315_), .Z(_02321__PTR0) );
  MUX2_X1 U7317 ( .A(P2_Datao_PTR1), .B(P2_EAX_PTR1), .S(_02315_), .Z(_02321__PTR1) );
  MUX2_X1 U7318 ( .A(P2_Datao_PTR2), .B(P2_EAX_PTR2), .S(_02315_), .Z(_02321__PTR2) );
  MUX2_X1 U7319 ( .A(P2_Datao_PTR3), .B(P2_EAX_PTR3), .S(_02315_), .Z(_02321__PTR3) );
  MUX2_X1 U7320 ( .A(P2_Datao_PTR4), .B(P2_EAX_PTR4), .S(_02315_), .Z(_02321__PTR4) );
  MUX2_X1 U7321 ( .A(P2_Datao_PTR5), .B(P2_EAX_PTR5), .S(_02315_), .Z(_02321__PTR5) );
  MUX2_X1 U7322 ( .A(P2_Datao_PTR6), .B(P2_EAX_PTR6), .S(_02315_), .Z(_02321__PTR6) );
  MUX2_X1 U7323 ( .A(P2_Datao_PTR7), .B(P2_EAX_PTR7), .S(_02315_), .Z(_02321__PTR7) );
  MUX2_X1 U7324 ( .A(P2_Datao_PTR8), .B(P2_EAX_PTR8), .S(_02315_), .Z(_02321__PTR8) );
  MUX2_X1 U7325 ( .A(P2_Datao_PTR9), .B(P2_EAX_PTR9), .S(_02315_), .Z(_02321__PTR9) );
  MUX2_X1 U7326 ( .A(P2_Datao_PTR10), .B(P2_EAX_PTR10), .S(_02315_), .Z(_02321__PTR10) );
  MUX2_X1 U7327 ( .A(P2_Datao_PTR11), .B(P2_EAX_PTR11), .S(_02315_), .Z(_02321__PTR11) );
  MUX2_X1 U7328 ( .A(P2_Datao_PTR12), .B(P2_EAX_PTR12), .S(_02315_), .Z(_02321__PTR12) );
  MUX2_X1 U7329 ( .A(P2_Datao_PTR13), .B(P2_EAX_PTR13), .S(_02315_), .Z(_02321__PTR13) );
  MUX2_X1 U7330 ( .A(P2_Datao_PTR14), .B(P2_EAX_PTR14), .S(_02315_), .Z(_02321__PTR14) );
  MUX2_X1 U7331 ( .A(P2_Datao_PTR15), .B(P2_EAX_PTR15), .S(_02315_), .Z(_02321__PTR15) );
  MUX2_X1 U7332 ( .A(P2_Datao_PTR16), .B(_03070__PTR0), .S(_02315_), .Z(_02321__PTR16) );
  MUX2_X1 U7333 ( .A(P2_Datao_PTR17), .B(_03071__PTR1), .S(_02315_), .Z(_02321__PTR17) );
  MUX2_X1 U7334 ( .A(P2_Datao_PTR18), .B(_03071__PTR2), .S(_02315_), .Z(_02321__PTR18) );
  MUX2_X1 U7335 ( .A(P2_Datao_PTR19), .B(_03071__PTR3), .S(_02315_), .Z(_02321__PTR19) );
  MUX2_X1 U7336 ( .A(P2_Datao_PTR20), .B(_03071__PTR4), .S(_02315_), .Z(_02321__PTR20) );
  MUX2_X1 U7337 ( .A(P2_Datao_PTR21), .B(_03071__PTR5), .S(_02315_), .Z(_02321__PTR21) );
  MUX2_X1 U7338 ( .A(P2_Datao_PTR22), .B(_03071__PTR6), .S(_02315_), .Z(_02321__PTR22) );
  MUX2_X1 U7339 ( .A(P2_Datao_PTR23), .B(_03071__PTR7), .S(_02315_), .Z(_02321__PTR23) );
  MUX2_X1 U7340 ( .A(P2_Datao_PTR24), .B(_03071__PTR8), .S(_02315_), .Z(_02321__PTR24) );
  MUX2_X1 U7341 ( .A(P2_Datao_PTR25), .B(_03071__PTR9), .S(_02315_), .Z(_02321__PTR25) );
  MUX2_X1 U7342 ( .A(P2_Datao_PTR26), .B(_03071__PTR10), .S(_02315_), .Z(_02321__PTR26) );
  MUX2_X1 U7343 ( .A(P2_Datao_PTR27), .B(_03071__PTR11), .S(_02315_), .Z(_02321__PTR27) );
  MUX2_X1 U7344 ( .A(P2_Datao_PTR28), .B(_03071__PTR12), .S(_02315_), .Z(_02321__PTR28) );
  MUX2_X1 U7345 ( .A(P2_Datao_PTR29), .B(_03071__PTR13), .S(_02315_), .Z(_02321__PTR29) );
  MUX2_X1 U7346 ( .A(P2_Datao_PTR30), .B(_03071__PTR14), .S(_02315_), .Z(_02321__PTR30) );
  MUX2_X1 U7347 ( .A(P2_ReadRequest), .B(1'b0), .S(_02296_), .Z(_02158__PTR0) );
  MUX2_X1 U7348 ( .A(P2_RequestPending), .B(_02322_), .S(_02296_), .Z(_02154__PTR2) );
  MUX2_X1 U7349 ( .A(P2_P1_InstQueueRd_Addr_PTR1), .B(_02310__PTR1), .S(_02315_), .Z(_02328__PTR1) );
  MUX2_X1 U7350 ( .A(P2_P1_InstQueueRd_Addr_PTR2), .B(_02310__PTR2), .S(_02315_), .Z(_02328__PTR2) );
  MUX2_X1 U7351 ( .A(P2_P1_InstQueueRd_Addr_PTR3), .B(_02310__PTR3), .S(_02315_), .Z(_02328__PTR3) );
  MUX2_X1 U7352 ( .A(P2_P1_InstQueueRd_Addr_PTR4), .B(_02310__PTR4), .S(_02315_), .Z(_02328__PTR4) );
  MUX2_X1 U7353 ( .A(P2_P1_InstAddrPointer_PTR1), .B(_02309__PTR1), .S(_02315_), .Z(_02327__PTR1) );
  MUX2_X1 U7354 ( .A(P2_P1_InstAddrPointer_PTR2), .B(_02309__PTR2), .S(_02315_), .Z(_02327__PTR2) );
  MUX2_X1 U7355 ( .A(P2_P1_InstAddrPointer_PTR3), .B(_02309__PTR3), .S(_02315_), .Z(_02327__PTR3) );
  MUX2_X1 U7356 ( .A(P2_P1_InstAddrPointer_PTR4), .B(_02309__PTR4), .S(_02315_), .Z(_02327__PTR4) );
  MUX2_X1 U7357 ( .A(P2_P1_InstAddrPointer_PTR5), .B(_02309__PTR5), .S(_02315_), .Z(_02327__PTR5) );
  MUX2_X1 U7358 ( .A(P2_P1_InstAddrPointer_PTR6), .B(_02309__PTR6), .S(_02315_), .Z(_02327__PTR6) );
  MUX2_X1 U7359 ( .A(P2_P1_InstAddrPointer_PTR7), .B(_02309__PTR7), .S(_02315_), .Z(_02327__PTR7) );
  MUX2_X1 U7360 ( .A(P2_P1_InstAddrPointer_PTR8), .B(_02309__PTR8), .S(_02315_), .Z(_02327__PTR8) );
  MUX2_X1 U7361 ( .A(P2_P1_InstAddrPointer_PTR9), .B(_02309__PTR9), .S(_02315_), .Z(_02327__PTR9) );
  MUX2_X1 U7362 ( .A(P2_P1_InstAddrPointer_PTR10), .B(_02309__PTR10), .S(_02315_), .Z(_02327__PTR10) );
  MUX2_X1 U7363 ( .A(P2_P1_InstAddrPointer_PTR11), .B(_02309__PTR11), .S(_02315_), .Z(_02327__PTR11) );
  MUX2_X1 U7364 ( .A(P2_P1_InstAddrPointer_PTR12), .B(_02309__PTR12), .S(_02315_), .Z(_02327__PTR12) );
  MUX2_X1 U7365 ( .A(P2_P1_InstAddrPointer_PTR13), .B(_02309__PTR13), .S(_02315_), .Z(_02327__PTR13) );
  MUX2_X1 U7366 ( .A(P2_P1_InstAddrPointer_PTR14), .B(_02309__PTR14), .S(_02315_), .Z(_02327__PTR14) );
  MUX2_X1 U7367 ( .A(P2_P1_InstAddrPointer_PTR15), .B(_02309__PTR15), .S(_02315_), .Z(_02327__PTR15) );
  MUX2_X1 U7368 ( .A(P2_P1_InstAddrPointer_PTR16), .B(_02309__PTR16), .S(_02315_), .Z(_02327__PTR16) );
  MUX2_X1 U7369 ( .A(P2_P1_InstAddrPointer_PTR17), .B(_02309__PTR17), .S(_02315_), .Z(_02327__PTR17) );
  MUX2_X1 U7370 ( .A(P2_P1_InstAddrPointer_PTR18), .B(_02309__PTR18), .S(_02315_), .Z(_02327__PTR18) );
  MUX2_X1 U7371 ( .A(P2_P1_InstAddrPointer_PTR19), .B(_02309__PTR19), .S(_02315_), .Z(_02327__PTR19) );
  MUX2_X1 U7372 ( .A(P2_P1_InstAddrPointer_PTR20), .B(_02309__PTR20), .S(_02315_), .Z(_02327__PTR20) );
  MUX2_X1 U7373 ( .A(P2_P1_InstAddrPointer_PTR21), .B(_02309__PTR21), .S(_02315_), .Z(_02327__PTR21) );
  MUX2_X1 U7374 ( .A(P2_P1_InstAddrPointer_PTR22), .B(_02309__PTR22), .S(_02315_), .Z(_02327__PTR22) );
  MUX2_X1 U7375 ( .A(P2_P1_InstAddrPointer_PTR23), .B(_02309__PTR23), .S(_02315_), .Z(_02327__PTR23) );
  MUX2_X1 U7376 ( .A(P2_P1_InstAddrPointer_PTR24), .B(_02309__PTR24), .S(_02315_), .Z(_02327__PTR24) );
  MUX2_X1 U7377 ( .A(P2_P1_InstAddrPointer_PTR25), .B(_02309__PTR25), .S(_02315_), .Z(_02327__PTR25) );
  MUX2_X1 U7378 ( .A(P2_P1_InstAddrPointer_PTR26), .B(_02309__PTR26), .S(_02315_), .Z(_02327__PTR26) );
  MUX2_X1 U7379 ( .A(P2_P1_InstAddrPointer_PTR27), .B(_02309__PTR27), .S(_02315_), .Z(_02327__PTR27) );
  MUX2_X1 U7380 ( .A(P2_P1_InstAddrPointer_PTR28), .B(_02309__PTR28), .S(_02315_), .Z(_02327__PTR28) );
  MUX2_X1 U7381 ( .A(P2_P1_InstAddrPointer_PTR29), .B(_02309__PTR29), .S(_02315_), .Z(_02327__PTR29) );
  MUX2_X1 U7382 ( .A(P2_P1_InstAddrPointer_PTR30), .B(_02309__PTR30), .S(_02315_), .Z(_02327__PTR30) );
  MUX2_X1 U7383 ( .A(P2_P1_InstAddrPointer_PTR31), .B(_02309__PTR31), .S(_02315_), .Z(_02327__PTR31) );
  MUX2_X1 U7384 ( .A(P2_P1_Flush), .B(_02308_), .S(_02315_), .Z(_02326_) );
  MUX2_X1 U7385 ( .A(P2_P1_More), .B(_02307_), .S(_02315_), .Z(_02325_) );
  MUX2_X1 U7386 ( .A(P2_P1_State2_PTR0), .B(_02320__PTR0), .S(_02315_), .Z(_02324__PTR0) );
  MUX2_X1 U7387 ( .A(P2_P1_State2_PTR1), .B(_02320__PTR1), .S(_02315_), .Z(_02324__PTR1) );
  MUX2_X1 U7388 ( .A(P2_P1_State2_PTR2), .B(_02320__PTR2), .S(_02315_), .Z(_02324__PTR2) );
  MUX2_X1 U7389 ( .A(P2_P1_State2_PTR3), .B(_02320__PTR3), .S(_02315_), .Z(_02324__PTR3) );
  MUX2_X1 U7390 ( .A(P2_EBX_PTR0), .B(_02305__PTR0), .S(_02315_), .Z(_02323__PTR0) );
  MUX2_X1 U7391 ( .A(P2_EBX_PTR1), .B(_02319__PTR1), .S(_02315_), .Z(_02323__PTR1) );
  MUX2_X1 U7392 ( .A(P2_EBX_PTR2), .B(_02319__PTR2), .S(_02315_), .Z(_02323__PTR2) );
  MUX2_X1 U7393 ( .A(P2_EBX_PTR3), .B(_02319__PTR3), .S(_02315_), .Z(_02323__PTR3) );
  MUX2_X1 U7394 ( .A(P2_EBX_PTR4), .B(_02319__PTR4), .S(_02315_), .Z(_02323__PTR4) );
  MUX2_X1 U7395 ( .A(P2_EBX_PTR5), .B(_02319__PTR5), .S(_02315_), .Z(_02323__PTR5) );
  MUX2_X1 U7396 ( .A(P2_EBX_PTR6), .B(_02319__PTR6), .S(_02315_), .Z(_02323__PTR6) );
  MUX2_X1 U7397 ( .A(P2_EBX_PTR7), .B(_02319__PTR7), .S(_02315_), .Z(_02323__PTR7) );
  MUX2_X1 U7398 ( .A(P2_EBX_PTR8), .B(_02319__PTR8), .S(_02315_), .Z(_02323__PTR8) );
  MUX2_X1 U7399 ( .A(P2_EBX_PTR9), .B(_02319__PTR9), .S(_02315_), .Z(_02323__PTR9) );
  MUX2_X1 U7400 ( .A(P2_EBX_PTR10), .B(_02319__PTR10), .S(_02315_), .Z(_02323__PTR10) );
  MUX2_X1 U7401 ( .A(P2_EBX_PTR11), .B(_02319__PTR11), .S(_02315_), .Z(_02323__PTR11) );
  MUX2_X1 U7402 ( .A(P2_EBX_PTR12), .B(_02319__PTR12), .S(_02315_), .Z(_02323__PTR12) );
  MUX2_X1 U7403 ( .A(P2_EBX_PTR13), .B(_02319__PTR13), .S(_02315_), .Z(_02323__PTR13) );
  MUX2_X1 U7404 ( .A(P2_EBX_PTR14), .B(_02319__PTR14), .S(_02315_), .Z(_02323__PTR14) );
  MUX2_X1 U7405 ( .A(P2_EBX_PTR15), .B(_02319__PTR15), .S(_02315_), .Z(_02323__PTR15) );
  MUX2_X1 U7406 ( .A(P2_EBX_PTR16), .B(_02319__PTR16), .S(_02315_), .Z(_02323__PTR16) );
  MUX2_X1 U7407 ( .A(P2_EBX_PTR17), .B(_02319__PTR17), .S(_02315_), .Z(_02323__PTR17) );
  MUX2_X1 U7408 ( .A(P2_EBX_PTR18), .B(_02319__PTR18), .S(_02315_), .Z(_02323__PTR18) );
  MUX2_X1 U7409 ( .A(P2_EBX_PTR19), .B(_02319__PTR19), .S(_02315_), .Z(_02323__PTR19) );
  MUX2_X1 U7410 ( .A(P2_EBX_PTR20), .B(_02319__PTR20), .S(_02315_), .Z(_02323__PTR20) );
  MUX2_X1 U7411 ( .A(P2_EBX_PTR21), .B(_02319__PTR21), .S(_02315_), .Z(_02323__PTR21) );
  MUX2_X1 U7412 ( .A(P2_EBX_PTR22), .B(_02319__PTR22), .S(_02315_), .Z(_02323__PTR22) );
  MUX2_X1 U7413 ( .A(P2_EBX_PTR23), .B(_02319__PTR23), .S(_02315_), .Z(_02323__PTR23) );
  MUX2_X1 U7414 ( .A(P2_EBX_PTR24), .B(_02319__PTR24), .S(_02315_), .Z(_02323__PTR24) );
  MUX2_X1 U7415 ( .A(P2_EBX_PTR25), .B(_02319__PTR25), .S(_02315_), .Z(_02323__PTR25) );
  MUX2_X1 U7416 ( .A(P2_EBX_PTR26), .B(_02319__PTR26), .S(_02315_), .Z(_02323__PTR26) );
  MUX2_X1 U7417 ( .A(P2_EBX_PTR27), .B(_02319__PTR27), .S(_02315_), .Z(_02323__PTR27) );
  MUX2_X1 U7418 ( .A(P2_EBX_PTR28), .B(_02319__PTR28), .S(_02315_), .Z(_02323__PTR28) );
  MUX2_X1 U7419 ( .A(P2_EBX_PTR29), .B(_02319__PTR29), .S(_02315_), .Z(_02323__PTR29) );
  MUX2_X1 U7420 ( .A(P2_EBX_PTR30), .B(_02319__PTR30), .S(_02315_), .Z(_02323__PTR30) );
  MUX2_X1 U7421 ( .A(P2_EBX_PTR31), .B(_02319__PTR31), .S(_02315_), .Z(_02323__PTR31) );
  MUX2_X1 U7422 ( .A(1'b1), .B(_02318_), .S(_02315_), .Z(_02322_) );
  MUX2_X1 U7423 ( .A(_02317__PTR0), .B(P2_P1_State2_PTR0), .S(P2_READY_n), .Z(_02320__PTR0) );
  MUX2_X1 U7424 ( .A(_02317__PTR1), .B(P2_P1_State2_PTR1), .S(P2_READY_n), .Z(_02320__PTR1) );
  MUX2_X1 U7425 ( .A(_02317__PTR2), .B(P2_P1_State2_PTR2), .S(P2_READY_n), .Z(_02320__PTR2) );
  MUX2_X1 U7426 ( .A(_02317__PTR3), .B(P2_P1_State2_PTR3), .S(P2_READY_n), .Z(_02320__PTR3) );
  MUX2_X1 U7427 ( .A(_02316__PTR1), .B(P2_EBX_PTR1), .S(P2_READY_n), .Z(_02319__PTR1) );
  MUX2_X1 U7428 ( .A(_02316__PTR2), .B(P2_EBX_PTR2), .S(P2_READY_n), .Z(_02319__PTR2) );
  MUX2_X1 U7429 ( .A(_02316__PTR3), .B(P2_EBX_PTR3), .S(P2_READY_n), .Z(_02319__PTR3) );
  MUX2_X1 U7430 ( .A(_02316__PTR4), .B(P2_EBX_PTR4), .S(P2_READY_n), .Z(_02319__PTR4) );
  MUX2_X1 U7431 ( .A(_02316__PTR5), .B(P2_EBX_PTR5), .S(P2_READY_n), .Z(_02319__PTR5) );
  MUX2_X1 U7432 ( .A(_02316__PTR6), .B(P2_EBX_PTR6), .S(P2_READY_n), .Z(_02319__PTR6) );
  MUX2_X1 U7433 ( .A(_02316__PTR7), .B(P2_EBX_PTR7), .S(P2_READY_n), .Z(_02319__PTR7) );
  MUX2_X1 U7434 ( .A(_02316__PTR8), .B(P2_EBX_PTR8), .S(P2_READY_n), .Z(_02319__PTR8) );
  MUX2_X1 U7435 ( .A(_02316__PTR9), .B(P2_EBX_PTR9), .S(P2_READY_n), .Z(_02319__PTR9) );
  MUX2_X1 U7436 ( .A(_02316__PTR10), .B(P2_EBX_PTR10), .S(P2_READY_n), .Z(_02319__PTR10) );
  MUX2_X1 U7437 ( .A(_02316__PTR11), .B(P2_EBX_PTR11), .S(P2_READY_n), .Z(_02319__PTR11) );
  MUX2_X1 U7438 ( .A(_02316__PTR12), .B(P2_EBX_PTR12), .S(P2_READY_n), .Z(_02319__PTR12) );
  MUX2_X1 U7439 ( .A(_02316__PTR13), .B(P2_EBX_PTR13), .S(P2_READY_n), .Z(_02319__PTR13) );
  MUX2_X1 U7440 ( .A(_02316__PTR14), .B(P2_EBX_PTR14), .S(P2_READY_n), .Z(_02319__PTR14) );
  MUX2_X1 U7441 ( .A(_02316__PTR15), .B(P2_EBX_PTR15), .S(P2_READY_n), .Z(_02319__PTR15) );
  MUX2_X1 U7442 ( .A(_02316__PTR16), .B(P2_EBX_PTR16), .S(P2_READY_n), .Z(_02319__PTR16) );
  MUX2_X1 U7443 ( .A(_02316__PTR17), .B(P2_EBX_PTR17), .S(P2_READY_n), .Z(_02319__PTR17) );
  MUX2_X1 U7444 ( .A(_02316__PTR18), .B(P2_EBX_PTR18), .S(P2_READY_n), .Z(_02319__PTR18) );
  MUX2_X1 U7445 ( .A(_02316__PTR19), .B(P2_EBX_PTR19), .S(P2_READY_n), .Z(_02319__PTR19) );
  MUX2_X1 U7446 ( .A(_02316__PTR20), .B(P2_EBX_PTR20), .S(P2_READY_n), .Z(_02319__PTR20) );
  MUX2_X1 U7447 ( .A(_02316__PTR21), .B(P2_EBX_PTR21), .S(P2_READY_n), .Z(_02319__PTR21) );
  MUX2_X1 U7448 ( .A(_02316__PTR22), .B(P2_EBX_PTR22), .S(P2_READY_n), .Z(_02319__PTR22) );
  MUX2_X1 U7449 ( .A(_02316__PTR23), .B(P2_EBX_PTR23), .S(P2_READY_n), .Z(_02319__PTR23) );
  MUX2_X1 U7450 ( .A(_02316__PTR24), .B(P2_EBX_PTR24), .S(P2_READY_n), .Z(_02319__PTR24) );
  MUX2_X1 U7451 ( .A(_02316__PTR25), .B(P2_EBX_PTR25), .S(P2_READY_n), .Z(_02319__PTR25) );
  MUX2_X1 U7452 ( .A(_02316__PTR26), .B(P2_EBX_PTR26), .S(P2_READY_n), .Z(_02319__PTR26) );
  MUX2_X1 U7453 ( .A(_02316__PTR27), .B(P2_EBX_PTR27), .S(P2_READY_n), .Z(_02319__PTR27) );
  MUX2_X1 U7454 ( .A(_02316__PTR28), .B(P2_EBX_PTR28), .S(P2_READY_n), .Z(_02319__PTR28) );
  MUX2_X1 U7455 ( .A(_02316__PTR29), .B(P2_EBX_PTR29), .S(P2_READY_n), .Z(_02319__PTR29) );
  MUX2_X1 U7456 ( .A(_02316__PTR30), .B(P2_EBX_PTR30), .S(P2_READY_n), .Z(_02319__PTR30) );
  MUX2_X1 U7457 ( .A(_02316__PTR31), .B(P2_EBX_PTR31), .S(P2_READY_n), .Z(_02319__PTR31) );
  MUX2_X1 U7458 ( .A(_02186__PTR9), .B(1'b1), .S(P2_READY_n), .Z(_02318_) );
  MUX2_X1 U7459 ( .A(1'b0), .B(P2_P1_State2_PTR0), .S(P2_StateBS16), .Z(_02317__PTR0) );
  MUX2_X1 U7460 ( .A(1'b1), .B(P2_P1_State2_PTR1), .S(P2_StateBS16), .Z(_02317__PTR1) );
  MUX2_X1 U7461 ( .A(1'b1), .B(P2_P1_State2_PTR2), .S(P2_StateBS16), .Z(_02317__PTR2) );
  MUX2_X1 U7462 ( .A(1'b0), .B(P2_P1_State2_PTR3), .S(P2_StateBS16), .Z(_02317__PTR3) );
  MUX2_X1 U7463 ( .A(_02174__PTR7), .B(P2_EBX_PTR1), .S(P2_StateBS16), .Z(_02316__PTR1) );
  MUX2_X1 U7464 ( .A(_03067__PTR1), .B(P2_EBX_PTR2), .S(P2_StateBS16), .Z(_02316__PTR2) );
  MUX2_X1 U7465 ( .A(_03067__PTR2), .B(P2_EBX_PTR3), .S(P2_StateBS16), .Z(_02316__PTR3) );
  MUX2_X1 U7466 ( .A(_03067__PTR3), .B(P2_EBX_PTR4), .S(P2_StateBS16), .Z(_02316__PTR4) );
  MUX2_X1 U7467 ( .A(_03067__PTR4), .B(P2_EBX_PTR5), .S(P2_StateBS16), .Z(_02316__PTR5) );
  MUX2_X1 U7468 ( .A(_03067__PTR5), .B(P2_EBX_PTR6), .S(P2_StateBS16), .Z(_02316__PTR6) );
  MUX2_X1 U7469 ( .A(_03067__PTR6), .B(P2_EBX_PTR7), .S(P2_StateBS16), .Z(_02316__PTR7) );
  MUX2_X1 U7470 ( .A(_03067__PTR7), .B(P2_EBX_PTR8), .S(P2_StateBS16), .Z(_02316__PTR8) );
  MUX2_X1 U7471 ( .A(_03067__PTR8), .B(P2_EBX_PTR9), .S(P2_StateBS16), .Z(_02316__PTR9) );
  MUX2_X1 U7472 ( .A(_03067__PTR9), .B(P2_EBX_PTR10), .S(P2_StateBS16), .Z(_02316__PTR10) );
  MUX2_X1 U7473 ( .A(_03067__PTR10), .B(P2_EBX_PTR11), .S(P2_StateBS16), .Z(_02316__PTR11) );
  MUX2_X1 U7474 ( .A(_03067__PTR11), .B(P2_EBX_PTR12), .S(P2_StateBS16), .Z(_02316__PTR12) );
  MUX2_X1 U7475 ( .A(_03067__PTR12), .B(P2_EBX_PTR13), .S(P2_StateBS16), .Z(_02316__PTR13) );
  MUX2_X1 U7476 ( .A(_03067__PTR13), .B(P2_EBX_PTR14), .S(P2_StateBS16), .Z(_02316__PTR14) );
  MUX2_X1 U7477 ( .A(_03067__PTR14), .B(P2_EBX_PTR15), .S(P2_StateBS16), .Z(_02316__PTR15) );
  MUX2_X1 U7478 ( .A(_03067__PTR15), .B(P2_EBX_PTR16), .S(P2_StateBS16), .Z(_02316__PTR16) );
  MUX2_X1 U7479 ( .A(_03067__PTR16), .B(P2_EBX_PTR17), .S(P2_StateBS16), .Z(_02316__PTR17) );
  MUX2_X1 U7480 ( .A(_03067__PTR17), .B(P2_EBX_PTR18), .S(P2_StateBS16), .Z(_02316__PTR18) );
  MUX2_X1 U7481 ( .A(_03067__PTR18), .B(P2_EBX_PTR19), .S(P2_StateBS16), .Z(_02316__PTR19) );
  MUX2_X1 U7482 ( .A(_03067__PTR19), .B(P2_EBX_PTR20), .S(P2_StateBS16), .Z(_02316__PTR20) );
  MUX2_X1 U7483 ( .A(_03067__PTR20), .B(P2_EBX_PTR21), .S(P2_StateBS16), .Z(_02316__PTR21) );
  MUX2_X1 U7484 ( .A(_03067__PTR21), .B(P2_EBX_PTR22), .S(P2_StateBS16), .Z(_02316__PTR22) );
  MUX2_X1 U7485 ( .A(_03067__PTR22), .B(P2_EBX_PTR23), .S(P2_StateBS16), .Z(_02316__PTR23) );
  MUX2_X1 U7486 ( .A(_03067__PTR23), .B(P2_EBX_PTR24), .S(P2_StateBS16), .Z(_02316__PTR24) );
  MUX2_X1 U7487 ( .A(_03067__PTR24), .B(P2_EBX_PTR25), .S(P2_StateBS16), .Z(_02316__PTR25) );
  MUX2_X1 U7488 ( .A(_03067__PTR25), .B(P2_EBX_PTR26), .S(P2_StateBS16), .Z(_02316__PTR26) );
  MUX2_X1 U7489 ( .A(_03067__PTR26), .B(P2_EBX_PTR27), .S(P2_StateBS16), .Z(_02316__PTR27) );
  MUX2_X1 U7490 ( .A(_03067__PTR27), .B(P2_EBX_PTR28), .S(P2_StateBS16), .Z(_02316__PTR28) );
  MUX2_X1 U7491 ( .A(_03067__PTR28), .B(P2_EBX_PTR29), .S(P2_StateBS16), .Z(_02316__PTR29) );
  MUX2_X1 U7492 ( .A(_03067__PTR29), .B(P2_EBX_PTR30), .S(P2_StateBS16), .Z(_02316__PTR30) );
  MUX2_X1 U7493 ( .A(_03067__PTR30), .B(P2_EBX_PTR31), .S(P2_StateBS16), .Z(_02316__PTR31) );
  MUX2_X1 U7494 ( .A(_03063__PTR3), .B(P2_P1_InstQueueRd_Addr_PTR4), .S(P2_READY_n), .Z(_02335__PTR4) );
  MUX2_X1 U7495 ( .A(_02182__PTR4), .B(P2_P1_InstQueueRd_Addr_PTR1), .S(P2_READY_n), .Z(_02310__PTR1) );
  MUX2_X1 U7496 ( .A(_02182__PTR5), .B(P2_P1_InstQueueRd_Addr_PTR2), .S(P2_READY_n), .Z(_02310__PTR2) );
  MUX2_X1 U7497 ( .A(_02182__PTR6), .B(P2_P1_InstQueueRd_Addr_PTR3), .S(P2_READY_n), .Z(_02310__PTR3) );
  MUX2_X1 U7498 ( .A(1'b0), .B(P2_P1_InstQueueRd_Addr_PTR4), .S(P2_READY_n), .Z(_02310__PTR4) );
  MUX2_X1 U7499 ( .A(P2_P1_lWord_PTR0), .B(P2_EAX_PTR0), .S(_02296_), .Z(_02400__PTR16) );
  MUX2_X1 U7500 ( .A(P2_P1_lWord_PTR1), .B(P2_EAX_PTR1), .S(_02296_), .Z(_02400__PTR17) );
  MUX2_X1 U7501 ( .A(P2_P1_lWord_PTR2), .B(P2_EAX_PTR2), .S(_02296_), .Z(_02400__PTR18) );
  MUX2_X1 U7502 ( .A(P2_P1_lWord_PTR3), .B(P2_EAX_PTR3), .S(_02296_), .Z(_02400__PTR19) );
  MUX2_X1 U7503 ( .A(P2_P1_lWord_PTR4), .B(P2_EAX_PTR4), .S(_02296_), .Z(_02400__PTR20) );
  MUX2_X1 U7504 ( .A(P2_P1_lWord_PTR5), .B(P2_EAX_PTR5), .S(_02296_), .Z(_02400__PTR21) );
  MUX2_X1 U7505 ( .A(P2_P1_lWord_PTR6), .B(P2_EAX_PTR6), .S(_02296_), .Z(_02400__PTR22) );
  MUX2_X1 U7506 ( .A(P2_P1_lWord_PTR7), .B(P2_EAX_PTR7), .S(_02296_), .Z(_02400__PTR23) );
  MUX2_X1 U7507 ( .A(P2_P1_lWord_PTR8), .B(P2_EAX_PTR8), .S(_02296_), .Z(_02400__PTR24) );
  MUX2_X1 U7508 ( .A(P2_P1_lWord_PTR9), .B(P2_EAX_PTR9), .S(_02296_), .Z(_02400__PTR25) );
  MUX2_X1 U7509 ( .A(P2_P1_lWord_PTR10), .B(P2_EAX_PTR10), .S(_02296_), .Z(_02400__PTR26) );
  MUX2_X1 U7510 ( .A(P2_P1_lWord_PTR11), .B(P2_EAX_PTR11), .S(_02296_), .Z(_02400__PTR27) );
  MUX2_X1 U7511 ( .A(P2_P1_lWord_PTR12), .B(P2_EAX_PTR12), .S(_02296_), .Z(_02400__PTR28) );
  MUX2_X1 U7512 ( .A(P2_P1_lWord_PTR13), .B(P2_EAX_PTR13), .S(_02296_), .Z(_02400__PTR29) );
  MUX2_X1 U7513 ( .A(P2_P1_lWord_PTR14), .B(P2_EAX_PTR14), .S(_02296_), .Z(_02400__PTR30) );
  MUX2_X1 U7514 ( .A(P2_P1_lWord_PTR15), .B(P2_EAX_PTR15), .S(_02296_), .Z(_02400__PTR31) );
  MUX2_X1 U7515 ( .A(P2_P1_lWord_PTR0), .B(_02304__PTR0), .S(_02296_), .Z(_02400__PTR32) );
  MUX2_X1 U7516 ( .A(P2_P1_lWord_PTR1), .B(_02304__PTR1), .S(_02296_), .Z(_02400__PTR33) );
  MUX2_X1 U7517 ( .A(P2_P1_lWord_PTR2), .B(_02304__PTR2), .S(_02296_), .Z(_02400__PTR34) );
  MUX2_X1 U7518 ( .A(P2_P1_lWord_PTR3), .B(_02304__PTR3), .S(_02296_), .Z(_02400__PTR35) );
  MUX2_X1 U7519 ( .A(P2_P1_lWord_PTR4), .B(_02304__PTR4), .S(_02296_), .Z(_02400__PTR36) );
  MUX2_X1 U7520 ( .A(P2_P1_lWord_PTR5), .B(_02304__PTR5), .S(_02296_), .Z(_02400__PTR37) );
  MUX2_X1 U7521 ( .A(P2_P1_lWord_PTR6), .B(_02304__PTR6), .S(_02296_), .Z(_02400__PTR38) );
  MUX2_X1 U7522 ( .A(P2_P1_lWord_PTR7), .B(_02304__PTR7), .S(_02296_), .Z(_02400__PTR39) );
  MUX2_X1 U7523 ( .A(P2_P1_lWord_PTR8), .B(_02304__PTR8), .S(_02296_), .Z(_02400__PTR40) );
  MUX2_X1 U7524 ( .A(P2_P1_lWord_PTR9), .B(_02304__PTR9), .S(_02296_), .Z(_02400__PTR41) );
  MUX2_X1 U7525 ( .A(P2_P1_lWord_PTR10), .B(_02304__PTR10), .S(_02296_), .Z(_02400__PTR42) );
  MUX2_X1 U7526 ( .A(P2_P1_lWord_PTR11), .B(_02304__PTR11), .S(_02296_), .Z(_02400__PTR43) );
  MUX2_X1 U7527 ( .A(P2_P1_lWord_PTR12), .B(_02304__PTR12), .S(_02296_), .Z(_02400__PTR44) );
  MUX2_X1 U7528 ( .A(P2_P1_lWord_PTR13), .B(_02304__PTR13), .S(_02296_), .Z(_02400__PTR45) );
  MUX2_X1 U7529 ( .A(P2_P1_lWord_PTR14), .B(_02304__PTR14), .S(_02296_), .Z(_02400__PTR46) );
  MUX2_X1 U7530 ( .A(P2_P1_lWord_PTR15), .B(_02304__PTR15), .S(_02296_), .Z(_02400__PTR47) );
  MUX2_X1 U7531 ( .A(1'b0), .B(_02308_), .S(_02296_), .Z(_02146__PTR1) );
  MUX2_X1 U7532 ( .A(1'b1), .B(_02307_), .S(_02296_), .Z(_02150__PTR1) );
  MUX2_X1 U7533 ( .A(di2_PTR16), .B(P2_EAX_PTR16), .S(P2_READY_n), .Z(_02334__PTR16) );
  MUX2_X1 U7534 ( .A(di2_PTR17), .B(P2_EAX_PTR17), .S(P2_READY_n), .Z(_02334__PTR17) );
  MUX2_X1 U7535 ( .A(di2_PTR18), .B(P2_EAX_PTR18), .S(P2_READY_n), .Z(_02334__PTR18) );
  MUX2_X1 U7536 ( .A(di2_PTR19), .B(P2_EAX_PTR19), .S(P2_READY_n), .Z(_02334__PTR19) );
  MUX2_X1 U7537 ( .A(di2_PTR20), .B(P2_EAX_PTR20), .S(P2_READY_n), .Z(_02334__PTR20) );
  MUX2_X1 U7538 ( .A(di2_PTR21), .B(P2_EAX_PTR21), .S(P2_READY_n), .Z(_02334__PTR21) );
  MUX2_X1 U7539 ( .A(di2_PTR22), .B(P2_EAX_PTR22), .S(P2_READY_n), .Z(_02334__PTR22) );
  MUX2_X1 U7540 ( .A(di2_PTR23), .B(P2_EAX_PTR23), .S(P2_READY_n), .Z(_02334__PTR23) );
  MUX2_X1 U7541 ( .A(di2_PTR24), .B(P2_EAX_PTR24), .S(P2_READY_n), .Z(_02334__PTR24) );
  MUX2_X1 U7542 ( .A(di2_PTR25), .B(P2_EAX_PTR25), .S(P2_READY_n), .Z(_02334__PTR25) );
  MUX2_X1 U7543 ( .A(di2_PTR26), .B(P2_EAX_PTR26), .S(P2_READY_n), .Z(_02334__PTR26) );
  MUX2_X1 U7544 ( .A(di2_PTR27), .B(P2_EAX_PTR27), .S(P2_READY_n), .Z(_02334__PTR27) );
  MUX2_X1 U7545 ( .A(di2_PTR28), .B(P2_EAX_PTR28), .S(P2_READY_n), .Z(_02334__PTR28) );
  MUX2_X1 U7546 ( .A(di2_PTR29), .B(P2_EAX_PTR29), .S(P2_READY_n), .Z(_02334__PTR29) );
  MUX2_X1 U7547 ( .A(di2_PTR30), .B(P2_EAX_PTR30), .S(P2_READY_n), .Z(_02334__PTR30) );
  MUX2_X1 U7548 ( .A(P2_Datai_PTR31), .B(P2_EAX_PTR31), .S(P2_READY_n), .Z(_02334__PTR31) );
  MUX2_X1 U7549 ( .A(di2_PTR0), .B(P2_EAX_PTR0), .S(P2_READY_n), .Z(_02306__PTR0) );
  MUX2_X1 U7550 ( .A(di2_PTR1), .B(P2_EAX_PTR1), .S(P2_READY_n), .Z(_02306__PTR1) );
  MUX2_X1 U7551 ( .A(di2_PTR2), .B(P2_EAX_PTR2), .S(P2_READY_n), .Z(_02306__PTR2) );
  MUX2_X1 U7552 ( .A(di2_PTR3), .B(P2_EAX_PTR3), .S(P2_READY_n), .Z(_02306__PTR3) );
  MUX2_X1 U7553 ( .A(di2_PTR4), .B(P2_EAX_PTR4), .S(P2_READY_n), .Z(_02306__PTR4) );
  MUX2_X1 U7554 ( .A(di2_PTR5), .B(P2_EAX_PTR5), .S(P2_READY_n), .Z(_02306__PTR5) );
  MUX2_X1 U7555 ( .A(di2_PTR6), .B(P2_EAX_PTR6), .S(P2_READY_n), .Z(_02306__PTR6) );
  MUX2_X1 U7556 ( .A(di2_PTR7), .B(P2_EAX_PTR7), .S(P2_READY_n), .Z(_02306__PTR7) );
  MUX2_X1 U7557 ( .A(di2_PTR8), .B(P2_EAX_PTR8), .S(P2_READY_n), .Z(_02306__PTR8) );
  MUX2_X1 U7558 ( .A(di2_PTR9), .B(P2_EAX_PTR9), .S(P2_READY_n), .Z(_02306__PTR9) );
  MUX2_X1 U7559 ( .A(di2_PTR10), .B(P2_EAX_PTR10), .S(P2_READY_n), .Z(_02306__PTR10) );
  MUX2_X1 U7560 ( .A(di2_PTR11), .B(P2_EAX_PTR11), .S(P2_READY_n), .Z(_02306__PTR11) );
  MUX2_X1 U7561 ( .A(di2_PTR12), .B(P2_EAX_PTR12), .S(P2_READY_n), .Z(_02306__PTR12) );
  MUX2_X1 U7562 ( .A(di2_PTR13), .B(P2_EAX_PTR13), .S(P2_READY_n), .Z(_02306__PTR13) );
  MUX2_X1 U7563 ( .A(di2_PTR14), .B(P2_EAX_PTR14), .S(P2_READY_n), .Z(_02306__PTR14) );
  MUX2_X1 U7564 ( .A(di2_PTR15), .B(P2_EAX_PTR15), .S(P2_READY_n), .Z(_02306__PTR15) );
  MUX2_X1 U7565 ( .A(di2_PTR0), .B(P2_EAX_PTR16), .S(P2_READY_n), .Z(_02306__PTR16) );
  MUX2_X1 U7566 ( .A(di2_PTR1), .B(P2_EAX_PTR17), .S(P2_READY_n), .Z(_02306__PTR17) );
  MUX2_X1 U7567 ( .A(di2_PTR2), .B(P2_EAX_PTR18), .S(P2_READY_n), .Z(_02306__PTR18) );
  MUX2_X1 U7568 ( .A(di2_PTR3), .B(P2_EAX_PTR19), .S(P2_READY_n), .Z(_02306__PTR19) );
  MUX2_X1 U7569 ( .A(di2_PTR4), .B(P2_EAX_PTR20), .S(P2_READY_n), .Z(_02306__PTR20) );
  MUX2_X1 U7570 ( .A(di2_PTR5), .B(P2_EAX_PTR21), .S(P2_READY_n), .Z(_02306__PTR21) );
  MUX2_X1 U7571 ( .A(di2_PTR6), .B(P2_EAX_PTR22), .S(P2_READY_n), .Z(_02306__PTR22) );
  MUX2_X1 U7572 ( .A(di2_PTR7), .B(P2_EAX_PTR23), .S(P2_READY_n), .Z(_02306__PTR23) );
  MUX2_X1 U7573 ( .A(di2_PTR8), .B(P2_EAX_PTR24), .S(P2_READY_n), .Z(_02306__PTR24) );
  MUX2_X1 U7574 ( .A(di2_PTR9), .B(P2_EAX_PTR25), .S(P2_READY_n), .Z(_02306__PTR25) );
  MUX2_X1 U7575 ( .A(di2_PTR10), .B(P2_EAX_PTR26), .S(P2_READY_n), .Z(_02306__PTR26) );
  MUX2_X1 U7576 ( .A(di2_PTR11), .B(P2_EAX_PTR27), .S(P2_READY_n), .Z(_02306__PTR27) );
  MUX2_X1 U7577 ( .A(di2_PTR12), .B(P2_EAX_PTR28), .S(P2_READY_n), .Z(_02306__PTR28) );
  MUX2_X1 U7578 ( .A(di2_PTR13), .B(P2_EAX_PTR29), .S(P2_READY_n), .Z(_02306__PTR29) );
  MUX2_X1 U7579 ( .A(di2_PTR14), .B(P2_EAX_PTR30), .S(P2_READY_n), .Z(_02306__PTR30) );
  MUX2_X1 U7580 ( .A(1'b0), .B(P2_EAX_PTR31), .S(P2_READY_n), .Z(_02306__PTR31) );
  MUX2_X1 U7581 ( .A(P2_P1_uWord_PTR0), .B(_03070__PTR0), .S(_02296_), .Z(_02396__PTR15) );
  MUX2_X1 U7582 ( .A(P2_P1_uWord_PTR1), .B(_03071__PTR1), .S(_02296_), .Z(_02396__PTR16) );
  MUX2_X1 U7583 ( .A(P2_P1_uWord_PTR2), .B(_03071__PTR2), .S(_02296_), .Z(_02396__PTR17) );
  MUX2_X1 U7584 ( .A(P2_P1_uWord_PTR3), .B(_03071__PTR3), .S(_02296_), .Z(_02396__PTR18) );
  MUX2_X1 U7585 ( .A(P2_P1_uWord_PTR4), .B(_03071__PTR4), .S(_02296_), .Z(_02396__PTR19) );
  MUX2_X1 U7586 ( .A(P2_P1_uWord_PTR5), .B(_03071__PTR5), .S(_02296_), .Z(_02396__PTR20) );
  MUX2_X1 U7587 ( .A(P2_P1_uWord_PTR6), .B(_03071__PTR6), .S(_02296_), .Z(_02396__PTR21) );
  MUX2_X1 U7588 ( .A(P2_P1_uWord_PTR7), .B(_03071__PTR7), .S(_02296_), .Z(_02396__PTR22) );
  MUX2_X1 U7589 ( .A(P2_P1_uWord_PTR8), .B(_03071__PTR8), .S(_02296_), .Z(_02396__PTR23) );
  MUX2_X1 U7590 ( .A(P2_P1_uWord_PTR9), .B(_03071__PTR9), .S(_02296_), .Z(_02396__PTR24) );
  MUX2_X1 U7591 ( .A(P2_P1_uWord_PTR10), .B(_03071__PTR10), .S(_02296_), .Z(_02396__PTR25) );
  MUX2_X1 U7592 ( .A(P2_P1_uWord_PTR11), .B(_03071__PTR11), .S(_02296_), .Z(_02396__PTR26) );
  MUX2_X1 U7593 ( .A(P2_P1_uWord_PTR12), .B(_03071__PTR12), .S(_02296_), .Z(_02396__PTR27) );
  MUX2_X1 U7594 ( .A(P2_P1_uWord_PTR13), .B(_03071__PTR13), .S(_02296_), .Z(_02396__PTR28) );
  MUX2_X1 U7595 ( .A(P2_P1_uWord_PTR14), .B(_03071__PTR14), .S(_02296_), .Z(_02396__PTR29) );
  MUX2_X1 U7596 ( .A(P2_P1_uWord_PTR0), .B(_02303__PTR0), .S(_02296_), .Z(_02396__PTR30) );
  MUX2_X1 U7597 ( .A(P2_P1_uWord_PTR1), .B(_02303__PTR1), .S(_02296_), .Z(_02396__PTR31) );
  MUX2_X1 U7598 ( .A(P2_P1_uWord_PTR2), .B(_02303__PTR2), .S(_02296_), .Z(_02396__PTR32) );
  MUX2_X1 U7599 ( .A(P2_P1_uWord_PTR3), .B(_02303__PTR3), .S(_02296_), .Z(_02396__PTR33) );
  MUX2_X1 U7600 ( .A(P2_P1_uWord_PTR4), .B(_02303__PTR4), .S(_02296_), .Z(_02396__PTR34) );
  MUX2_X1 U7601 ( .A(P2_P1_uWord_PTR5), .B(_02303__PTR5), .S(_02296_), .Z(_02396__PTR35) );
  MUX2_X1 U7602 ( .A(P2_P1_uWord_PTR6), .B(_02303__PTR6), .S(_02296_), .Z(_02396__PTR36) );
  MUX2_X1 U7603 ( .A(P2_P1_uWord_PTR7), .B(_02303__PTR7), .S(_02296_), .Z(_02396__PTR37) );
  MUX2_X1 U7604 ( .A(P2_P1_uWord_PTR8), .B(_02303__PTR8), .S(_02296_), .Z(_02396__PTR38) );
  MUX2_X1 U7605 ( .A(P2_P1_uWord_PTR9), .B(_02303__PTR9), .S(_02296_), .Z(_02396__PTR39) );
  MUX2_X1 U7606 ( .A(P2_P1_uWord_PTR10), .B(_02303__PTR10), .S(_02296_), .Z(_02396__PTR40) );
  MUX2_X1 U7607 ( .A(P2_P1_uWord_PTR11), .B(_02303__PTR11), .S(_02296_), .Z(_02396__PTR41) );
  MUX2_X1 U7608 ( .A(P2_P1_uWord_PTR12), .B(_02303__PTR12), .S(_02296_), .Z(_02396__PTR42) );
  MUX2_X1 U7609 ( .A(P2_P1_uWord_PTR13), .B(_02303__PTR13), .S(_02296_), .Z(_02396__PTR43) );
  MUX2_X1 U7610 ( .A(P2_P1_uWord_PTR14), .B(_02303__PTR14), .S(_02296_), .Z(_02396__PTR44) );
  MUX2_X1 U7611 ( .A(P2_CodeFetch), .B(1'b0), .S(_02296_), .Z(_02165__PTR0) );
  MUX2_X1 U7612 ( .A(P2_MemoryFetch), .B(1'b1), .S(_02296_), .Z(_02161__PTR1) );
  MUX2_X1 U7613 ( .A(P2_ReadRequest), .B(1'b1), .S(_02296_), .Z(_02158__PTR1) );
  MUX2_X1 U7614 ( .A(P2_RequestPending), .B(P2_READY_n), .S(_02296_), .Z(_02154__PTR1) );
  MUX2_X1 U7615 ( .A(P2_P1_InstQueueRd_Addr_PTR4), .B(_02335__PTR4), .S(_02296_), .Z(_02377__PTR19) );
  MUX2_X1 U7616 ( .A(P2_P1_InstQueueRd_Addr_PTR1), .B(_02328__PTR1), .S(_02296_), .Z(_02377__PTR11) );
  MUX2_X1 U7617 ( .A(P2_P1_InstQueueRd_Addr_PTR2), .B(_02328__PTR2), .S(_02296_), .Z(_02377__PTR12) );
  MUX2_X1 U7618 ( .A(P2_P1_InstQueueRd_Addr_PTR3), .B(_02328__PTR3), .S(_02296_), .Z(_02377__PTR13) );
  MUX2_X1 U7619 ( .A(P2_P1_InstQueueRd_Addr_PTR4), .B(_02328__PTR4), .S(_02296_), .Z(_02377__PTR14) );
  MUX2_X1 U7620 ( .A(P2_P1_InstQueueRd_Addr_PTR1), .B(_02310__PTR1), .S(_02296_), .Z(_02377__PTR21) );
  MUX2_X1 U7621 ( .A(P2_P1_InstQueueRd_Addr_PTR2), .B(_02310__PTR2), .S(_02296_), .Z(_02377__PTR22) );
  MUX2_X1 U7622 ( .A(P2_P1_InstQueueRd_Addr_PTR3), .B(_02310__PTR3), .S(_02296_), .Z(_02377__PTR23) );
  MUX2_X1 U7623 ( .A(P2_P1_InstQueueRd_Addr_PTR4), .B(_02310__PTR4), .S(_02296_), .Z(_02377__PTR24) );
  MUX2_X1 U7624 ( .A(_02373__PTR33), .B(P2_P1_InstAddrPointer_PTR1), .S(P2_READY_n), .Z(_02309__PTR1) );
  MUX2_X1 U7625 ( .A(_02373__PTR34), .B(P2_P1_InstAddrPointer_PTR2), .S(P2_READY_n), .Z(_02309__PTR2) );
  MUX2_X1 U7626 ( .A(_02373__PTR35), .B(P2_P1_InstAddrPointer_PTR3), .S(P2_READY_n), .Z(_02309__PTR3) );
  MUX2_X1 U7627 ( .A(_02373__PTR36), .B(P2_P1_InstAddrPointer_PTR4), .S(P2_READY_n), .Z(_02309__PTR4) );
  MUX2_X1 U7628 ( .A(_02373__PTR37), .B(P2_P1_InstAddrPointer_PTR5), .S(P2_READY_n), .Z(_02309__PTR5) );
  MUX2_X1 U7629 ( .A(_02373__PTR38), .B(P2_P1_InstAddrPointer_PTR6), .S(P2_READY_n), .Z(_02309__PTR6) );
  MUX2_X1 U7630 ( .A(_02373__PTR39), .B(P2_P1_InstAddrPointer_PTR7), .S(P2_READY_n), .Z(_02309__PTR7) );
  MUX2_X1 U7631 ( .A(_02373__PTR40), .B(P2_P1_InstAddrPointer_PTR8), .S(P2_READY_n), .Z(_02309__PTR8) );
  MUX2_X1 U7632 ( .A(_02373__PTR41), .B(P2_P1_InstAddrPointer_PTR9), .S(P2_READY_n), .Z(_02309__PTR9) );
  MUX2_X1 U7633 ( .A(_02373__PTR42), .B(P2_P1_InstAddrPointer_PTR10), .S(P2_READY_n), .Z(_02309__PTR10) );
  MUX2_X1 U7634 ( .A(_02373__PTR43), .B(P2_P1_InstAddrPointer_PTR11), .S(P2_READY_n), .Z(_02309__PTR11) );
  MUX2_X1 U7635 ( .A(_02373__PTR44), .B(P2_P1_InstAddrPointer_PTR12), .S(P2_READY_n), .Z(_02309__PTR12) );
  MUX2_X1 U7636 ( .A(_02373__PTR45), .B(P2_P1_InstAddrPointer_PTR13), .S(P2_READY_n), .Z(_02309__PTR13) );
  MUX2_X1 U7637 ( .A(_02373__PTR46), .B(P2_P1_InstAddrPointer_PTR14), .S(P2_READY_n), .Z(_02309__PTR14) );
  MUX2_X1 U7638 ( .A(_02373__PTR47), .B(P2_P1_InstAddrPointer_PTR15), .S(P2_READY_n), .Z(_02309__PTR15) );
  MUX2_X1 U7639 ( .A(_02373__PTR48), .B(P2_P1_InstAddrPointer_PTR16), .S(P2_READY_n), .Z(_02309__PTR16) );
  MUX2_X1 U7640 ( .A(_02373__PTR49), .B(P2_P1_InstAddrPointer_PTR17), .S(P2_READY_n), .Z(_02309__PTR17) );
  MUX2_X1 U7641 ( .A(_02373__PTR50), .B(P2_P1_InstAddrPointer_PTR18), .S(P2_READY_n), .Z(_02309__PTR18) );
  MUX2_X1 U7642 ( .A(_02373__PTR51), .B(P2_P1_InstAddrPointer_PTR19), .S(P2_READY_n), .Z(_02309__PTR19) );
  MUX2_X1 U7643 ( .A(_02373__PTR52), .B(P2_P1_InstAddrPointer_PTR20), .S(P2_READY_n), .Z(_02309__PTR20) );
  MUX2_X1 U7644 ( .A(_02373__PTR53), .B(P2_P1_InstAddrPointer_PTR21), .S(P2_READY_n), .Z(_02309__PTR21) );
  MUX2_X1 U7645 ( .A(_02373__PTR54), .B(P2_P1_InstAddrPointer_PTR22), .S(P2_READY_n), .Z(_02309__PTR22) );
  MUX2_X1 U7646 ( .A(_02373__PTR55), .B(P2_P1_InstAddrPointer_PTR23), .S(P2_READY_n), .Z(_02309__PTR23) );
  MUX2_X1 U7647 ( .A(_02373__PTR56), .B(P2_P1_InstAddrPointer_PTR24), .S(P2_READY_n), .Z(_02309__PTR24) );
  MUX2_X1 U7648 ( .A(_02373__PTR57), .B(P2_P1_InstAddrPointer_PTR25), .S(P2_READY_n), .Z(_02309__PTR25) );
  MUX2_X1 U7649 ( .A(_02373__PTR58), .B(P2_P1_InstAddrPointer_PTR26), .S(P2_READY_n), .Z(_02309__PTR26) );
  MUX2_X1 U7650 ( .A(_02373__PTR59), .B(P2_P1_InstAddrPointer_PTR27), .S(P2_READY_n), .Z(_02309__PTR27) );
  MUX2_X1 U7651 ( .A(_02373__PTR60), .B(P2_P1_InstAddrPointer_PTR28), .S(P2_READY_n), .Z(_02309__PTR28) );
  MUX2_X1 U7652 ( .A(_02373__PTR61), .B(P2_P1_InstAddrPointer_PTR29), .S(P2_READY_n), .Z(_02309__PTR29) );
  MUX2_X1 U7653 ( .A(_02373__PTR62), .B(P2_P1_InstAddrPointer_PTR30), .S(P2_READY_n), .Z(_02309__PTR30) );
  MUX2_X1 U7654 ( .A(_02373__PTR63), .B(P2_P1_InstAddrPointer_PTR31), .S(P2_READY_n), .Z(_02309__PTR31) );
  MUX2_X1 U7655 ( .A(1'b0), .B(P2_P1_Flush), .S(P2_READY_n), .Z(_02308_) );
  MUX2_X1 U7656 ( .A(1'b0), .B(P2_P1_More), .S(P2_READY_n), .Z(_02307_) );
  MUX2_X1 U7657 ( .A(_02300__PTR0), .B(P2_EBX_PTR0), .S(P2_READY_n), .Z(_02305__PTR0) );
  MUX2_X1 U7658 ( .A(_02300__PTR1), .B(_02299__PTR1), .S(P2_READY_n), .Z(_02305__PTR1) );
  MUX2_X1 U7659 ( .A(_02300__PTR2), .B(_02299__PTR2), .S(P2_READY_n), .Z(_02305__PTR2) );
  MUX2_X1 U7660 ( .A(_02300__PTR3), .B(_02299__PTR3), .S(P2_READY_n), .Z(_02305__PTR3) );
  MUX2_X1 U7661 ( .A(_02300__PTR4), .B(_02299__PTR4), .S(P2_READY_n), .Z(_02305__PTR4) );
  MUX2_X1 U7662 ( .A(_02300__PTR5), .B(_02299__PTR5), .S(P2_READY_n), .Z(_02305__PTR5) );
  MUX2_X1 U7663 ( .A(_02300__PTR6), .B(_02299__PTR6), .S(P2_READY_n), .Z(_02305__PTR6) );
  MUX2_X1 U7664 ( .A(_02300__PTR7), .B(_02299__PTR7), .S(P2_READY_n), .Z(_02305__PTR7) );
  MUX2_X1 U7665 ( .A(_02300__PTR8), .B(_02299__PTR8), .S(P2_READY_n), .Z(_02305__PTR8) );
  MUX2_X1 U7666 ( .A(_02300__PTR9), .B(_02299__PTR9), .S(P2_READY_n), .Z(_02305__PTR9) );
  MUX2_X1 U7667 ( .A(_02300__PTR10), .B(_02299__PTR10), .S(P2_READY_n), .Z(_02305__PTR10) );
  MUX2_X1 U7668 ( .A(_02300__PTR11), .B(_02299__PTR11), .S(P2_READY_n), .Z(_02305__PTR11) );
  MUX2_X1 U7669 ( .A(_02300__PTR12), .B(_02299__PTR12), .S(P2_READY_n), .Z(_02305__PTR12) );
  MUX2_X1 U7670 ( .A(_02300__PTR13), .B(_02299__PTR13), .S(P2_READY_n), .Z(_02305__PTR13) );
  MUX2_X1 U7671 ( .A(_02300__PTR14), .B(_02299__PTR14), .S(P2_READY_n), .Z(_02305__PTR14) );
  MUX2_X1 U7672 ( .A(_02300__PTR15), .B(_02299__PTR15), .S(P2_READY_n), .Z(_02305__PTR15) );
  MUX2_X1 U7673 ( .A(_02300__PTR16), .B(_02299__PTR16), .S(P2_READY_n), .Z(_02305__PTR16) );
  MUX2_X1 U7674 ( .A(_02300__PTR17), .B(_02299__PTR17), .S(P2_READY_n), .Z(_02305__PTR17) );
  MUX2_X1 U7675 ( .A(_02300__PTR18), .B(_02299__PTR18), .S(P2_READY_n), .Z(_02305__PTR18) );
  MUX2_X1 U7676 ( .A(_02300__PTR19), .B(_02299__PTR19), .S(P2_READY_n), .Z(_02305__PTR19) );
  MUX2_X1 U7677 ( .A(_02300__PTR20), .B(_02299__PTR20), .S(P2_READY_n), .Z(_02305__PTR20) );
  MUX2_X1 U7678 ( .A(_02300__PTR21), .B(_02299__PTR21), .S(P2_READY_n), .Z(_02305__PTR21) );
  MUX2_X1 U7679 ( .A(_02300__PTR22), .B(_02299__PTR22), .S(P2_READY_n), .Z(_02305__PTR22) );
  MUX2_X1 U7680 ( .A(_02300__PTR23), .B(_02299__PTR23), .S(P2_READY_n), .Z(_02305__PTR23) );
  MUX2_X1 U7681 ( .A(_02300__PTR24), .B(_02299__PTR24), .S(P2_READY_n), .Z(_02305__PTR24) );
  MUX2_X1 U7682 ( .A(_02300__PTR25), .B(_02299__PTR25), .S(P2_READY_n), .Z(_02305__PTR25) );
  MUX2_X1 U7683 ( .A(_02300__PTR26), .B(_02299__PTR26), .S(P2_READY_n), .Z(_02305__PTR26) );
  MUX2_X1 U7684 ( .A(_02300__PTR27), .B(_02299__PTR27), .S(P2_READY_n), .Z(_02305__PTR27) );
  MUX2_X1 U7685 ( .A(_02300__PTR28), .B(_02299__PTR28), .S(P2_READY_n), .Z(_02305__PTR28) );
  MUX2_X1 U7686 ( .A(_02300__PTR29), .B(_02299__PTR29), .S(P2_READY_n), .Z(_02305__PTR29) );
  MUX2_X1 U7687 ( .A(_02300__PTR30), .B(_02299__PTR30), .S(P2_READY_n), .Z(_02305__PTR30) );
  MUX2_X1 U7688 ( .A(_02300__PTR31), .B(_02299__PTR31), .S(P2_READY_n), .Z(_02305__PTR31) );
  MUX2_X1 U7689 ( .A(di2_PTR0), .B(P2_P1_lWord_PTR0), .S(P2_READY_n), .Z(_02304__PTR0) );
  MUX2_X1 U7690 ( .A(di2_PTR1), .B(P2_P1_lWord_PTR1), .S(P2_READY_n), .Z(_02304__PTR1) );
  MUX2_X1 U7691 ( .A(di2_PTR2), .B(P2_P1_lWord_PTR2), .S(P2_READY_n), .Z(_02304__PTR2) );
  MUX2_X1 U7692 ( .A(di2_PTR3), .B(P2_P1_lWord_PTR3), .S(P2_READY_n), .Z(_02304__PTR3) );
  MUX2_X1 U7693 ( .A(di2_PTR4), .B(P2_P1_lWord_PTR4), .S(P2_READY_n), .Z(_02304__PTR4) );
  MUX2_X1 U7694 ( .A(di2_PTR5), .B(P2_P1_lWord_PTR5), .S(P2_READY_n), .Z(_02304__PTR5) );
  MUX2_X1 U7695 ( .A(di2_PTR6), .B(P2_P1_lWord_PTR6), .S(P2_READY_n), .Z(_02304__PTR6) );
  MUX2_X1 U7696 ( .A(di2_PTR7), .B(P2_P1_lWord_PTR7), .S(P2_READY_n), .Z(_02304__PTR7) );
  MUX2_X1 U7697 ( .A(di2_PTR8), .B(P2_P1_lWord_PTR8), .S(P2_READY_n), .Z(_02304__PTR8) );
  MUX2_X1 U7698 ( .A(di2_PTR9), .B(P2_P1_lWord_PTR9), .S(P2_READY_n), .Z(_02304__PTR9) );
  MUX2_X1 U7699 ( .A(di2_PTR10), .B(P2_P1_lWord_PTR10), .S(P2_READY_n), .Z(_02304__PTR10) );
  MUX2_X1 U7700 ( .A(di2_PTR11), .B(P2_P1_lWord_PTR11), .S(P2_READY_n), .Z(_02304__PTR11) );
  MUX2_X1 U7701 ( .A(di2_PTR12), .B(P2_P1_lWord_PTR12), .S(P2_READY_n), .Z(_02304__PTR12) );
  MUX2_X1 U7702 ( .A(di2_PTR13), .B(P2_P1_lWord_PTR13), .S(P2_READY_n), .Z(_02304__PTR13) );
  MUX2_X1 U7703 ( .A(di2_PTR14), .B(P2_P1_lWord_PTR14), .S(P2_READY_n), .Z(_02304__PTR14) );
  MUX2_X1 U7704 ( .A(di2_PTR15), .B(P2_P1_lWord_PTR15), .S(P2_READY_n), .Z(_02304__PTR15) );
  MUX2_X1 U7705 ( .A(di2_PTR0), .B(P2_P1_uWord_PTR0), .S(P2_READY_n), .Z(_02303__PTR0) );
  MUX2_X1 U7706 ( .A(di2_PTR1), .B(P2_P1_uWord_PTR1), .S(P2_READY_n), .Z(_02303__PTR1) );
  MUX2_X1 U7707 ( .A(di2_PTR2), .B(P2_P1_uWord_PTR2), .S(P2_READY_n), .Z(_02303__PTR2) );
  MUX2_X1 U7708 ( .A(di2_PTR3), .B(P2_P1_uWord_PTR3), .S(P2_READY_n), .Z(_02303__PTR3) );
  MUX2_X1 U7709 ( .A(di2_PTR4), .B(P2_P1_uWord_PTR4), .S(P2_READY_n), .Z(_02303__PTR4) );
  MUX2_X1 U7710 ( .A(di2_PTR5), .B(P2_P1_uWord_PTR5), .S(P2_READY_n), .Z(_02303__PTR5) );
  MUX2_X1 U7711 ( .A(di2_PTR6), .B(P2_P1_uWord_PTR6), .S(P2_READY_n), .Z(_02303__PTR6) );
  MUX2_X1 U7712 ( .A(di2_PTR7), .B(P2_P1_uWord_PTR7), .S(P2_READY_n), .Z(_02303__PTR7) );
  MUX2_X1 U7713 ( .A(di2_PTR8), .B(P2_P1_uWord_PTR8), .S(P2_READY_n), .Z(_02303__PTR8) );
  MUX2_X1 U7714 ( .A(di2_PTR9), .B(P2_P1_uWord_PTR9), .S(P2_READY_n), .Z(_02303__PTR9) );
  MUX2_X1 U7715 ( .A(di2_PTR10), .B(P2_P1_uWord_PTR10), .S(P2_READY_n), .Z(_02303__PTR10) );
  MUX2_X1 U7716 ( .A(di2_PTR11), .B(P2_P1_uWord_PTR11), .S(P2_READY_n), .Z(_02303__PTR11) );
  MUX2_X1 U7717 ( .A(di2_PTR12), .B(P2_P1_uWord_PTR12), .S(P2_READY_n), .Z(_02303__PTR12) );
  MUX2_X1 U7718 ( .A(di2_PTR13), .B(P2_P1_uWord_PTR13), .S(P2_READY_n), .Z(_02303__PTR13) );
  MUX2_X1 U7719 ( .A(di2_PTR14), .B(P2_P1_uWord_PTR14), .S(P2_READY_n), .Z(_02303__PTR14) );
  MUX2_X1 U7720 ( .A(P2_P1_InstAddrPointer_PTR0), .B(_02373__PTR0), .S(_02146__PTR2), .Z(_02373__PTR128) );
  MUX2_X1 U7721 ( .A(P2_P1_InstAddrPointer_PTR1), .B(_02373__PTR1), .S(_02146__PTR2), .Z(_02373__PTR129) );
  MUX2_X1 U7722 ( .A(P2_P1_InstAddrPointer_PTR2), .B(_03052__PTR2), .S(_02146__PTR2), .Z(_02373__PTR130) );
  MUX2_X1 U7723 ( .A(P2_P1_InstAddrPointer_PTR3), .B(_03052__PTR3), .S(_02146__PTR2), .Z(_02373__PTR131) );
  MUX2_X1 U7724 ( .A(P2_P1_InstAddrPointer_PTR4), .B(_03052__PTR4), .S(_02146__PTR2), .Z(_02373__PTR132) );
  MUX2_X1 U7725 ( .A(P2_P1_InstAddrPointer_PTR5), .B(_03052__PTR5), .S(_02146__PTR2), .Z(_02373__PTR133) );
  MUX2_X1 U7726 ( .A(P2_P1_InstAddrPointer_PTR6), .B(_03052__PTR6), .S(_02146__PTR2), .Z(_02373__PTR134) );
  MUX2_X1 U7727 ( .A(P2_P1_InstAddrPointer_PTR7), .B(_03052__PTR7), .S(_02146__PTR2), .Z(_02373__PTR135) );
  MUX2_X1 U7728 ( .A(P2_P1_InstAddrPointer_PTR8), .B(_03052__PTR8), .S(_02146__PTR2), .Z(_02373__PTR136) );
  MUX2_X1 U7729 ( .A(P2_P1_InstAddrPointer_PTR9), .B(_03052__PTR9), .S(_02146__PTR2), .Z(_02373__PTR137) );
  MUX2_X1 U7730 ( .A(P2_P1_InstAddrPointer_PTR10), .B(_03052__PTR10), .S(_02146__PTR2), .Z(_02373__PTR138) );
  MUX2_X1 U7731 ( .A(P2_P1_InstAddrPointer_PTR11), .B(_03052__PTR11), .S(_02146__PTR2), .Z(_02373__PTR139) );
  MUX2_X1 U7732 ( .A(P2_P1_InstAddrPointer_PTR12), .B(_03052__PTR12), .S(_02146__PTR2), .Z(_02373__PTR140) );
  MUX2_X1 U7733 ( .A(P2_P1_InstAddrPointer_PTR13), .B(_03052__PTR13), .S(_02146__PTR2), .Z(_02373__PTR141) );
  MUX2_X1 U7734 ( .A(P2_P1_InstAddrPointer_PTR14), .B(_03052__PTR14), .S(_02146__PTR2), .Z(_02373__PTR142) );
  MUX2_X1 U7735 ( .A(P2_P1_InstAddrPointer_PTR15), .B(_03052__PTR15), .S(_02146__PTR2), .Z(_02373__PTR143) );
  MUX2_X1 U7736 ( .A(P2_P1_InstAddrPointer_PTR16), .B(_03052__PTR16), .S(_02146__PTR2), .Z(_02373__PTR144) );
  MUX2_X1 U7737 ( .A(P2_P1_InstAddrPointer_PTR17), .B(_03052__PTR17), .S(_02146__PTR2), .Z(_02373__PTR145) );
  MUX2_X1 U7738 ( .A(P2_P1_InstAddrPointer_PTR18), .B(_03052__PTR18), .S(_02146__PTR2), .Z(_02373__PTR146) );
  MUX2_X1 U7739 ( .A(P2_P1_InstAddrPointer_PTR19), .B(_03052__PTR19), .S(_02146__PTR2), .Z(_02373__PTR147) );
  MUX2_X1 U7740 ( .A(P2_P1_InstAddrPointer_PTR20), .B(_03052__PTR20), .S(_02146__PTR2), .Z(_02373__PTR148) );
  MUX2_X1 U7741 ( .A(P2_P1_InstAddrPointer_PTR21), .B(_03052__PTR21), .S(_02146__PTR2), .Z(_02373__PTR149) );
  MUX2_X1 U7742 ( .A(P2_P1_InstAddrPointer_PTR22), .B(_03052__PTR22), .S(_02146__PTR2), .Z(_02373__PTR150) );
  MUX2_X1 U7743 ( .A(P2_P1_InstAddrPointer_PTR23), .B(_03052__PTR23), .S(_02146__PTR2), .Z(_02373__PTR151) );
  MUX2_X1 U7744 ( .A(P2_P1_InstAddrPointer_PTR24), .B(_03052__PTR24), .S(_02146__PTR2), .Z(_02373__PTR152) );
  MUX2_X1 U7745 ( .A(P2_P1_InstAddrPointer_PTR25), .B(_03052__PTR25), .S(_02146__PTR2), .Z(_02373__PTR153) );
  MUX2_X1 U7746 ( .A(P2_P1_InstAddrPointer_PTR26), .B(_03052__PTR26), .S(_02146__PTR2), .Z(_02373__PTR154) );
  MUX2_X1 U7747 ( .A(P2_P1_InstAddrPointer_PTR27), .B(_03052__PTR27), .S(_02146__PTR2), .Z(_02373__PTR155) );
  MUX2_X1 U7748 ( .A(P2_P1_InstAddrPointer_PTR28), .B(_03052__PTR28), .S(_02146__PTR2), .Z(_02373__PTR156) );
  MUX2_X1 U7749 ( .A(P2_P1_InstAddrPointer_PTR29), .B(_03052__PTR29), .S(_02146__PTR2), .Z(_02373__PTR157) );
  MUX2_X1 U7750 ( .A(P2_P1_InstAddrPointer_PTR30), .B(_03052__PTR30), .S(_02146__PTR2), .Z(_02373__PTR158) );
  MUX2_X1 U7751 ( .A(P2_P1_InstAddrPointer_PTR31), .B(_03052__PTR31), .S(_02146__PTR2), .Z(_02373__PTR159) );
  MUX2_X1 U7752 ( .A(P2_P1_InstAddrPointer_PTR0), .B(_03054__PTR0), .S(_02146__PTR2), .Z(_02373__PTR160) );
  MUX2_X1 U7753 ( .A(P2_P1_InstAddrPointer_PTR1), .B(_03055__PTR1), .S(_02146__PTR2), .Z(_02373__PTR161) );
  MUX2_X1 U7754 ( .A(P2_P1_InstAddrPointer_PTR2), .B(_03055__PTR2), .S(_02146__PTR2), .Z(_02373__PTR162) );
  MUX2_X1 U7755 ( .A(P2_P1_InstAddrPointer_PTR3), .B(_03055__PTR3), .S(_02146__PTR2), .Z(_02373__PTR163) );
  MUX2_X1 U7756 ( .A(P2_P1_InstAddrPointer_PTR4), .B(_03055__PTR4), .S(_02146__PTR2), .Z(_02373__PTR164) );
  MUX2_X1 U7757 ( .A(P2_P1_InstAddrPointer_PTR5), .B(_03055__PTR5), .S(_02146__PTR2), .Z(_02373__PTR165) );
  MUX2_X1 U7758 ( .A(P2_P1_InstAddrPointer_PTR6), .B(_03055__PTR6), .S(_02146__PTR2), .Z(_02373__PTR166) );
  MUX2_X1 U7759 ( .A(P2_P1_InstAddrPointer_PTR7), .B(_03055__PTR7), .S(_02146__PTR2), .Z(_02373__PTR167) );
  MUX2_X1 U7760 ( .A(P2_P1_InstAddrPointer_PTR8), .B(_03055__PTR8), .S(_02146__PTR2), .Z(_02373__PTR168) );
  MUX2_X1 U7761 ( .A(P2_P1_InstAddrPointer_PTR9), .B(_03055__PTR9), .S(_02146__PTR2), .Z(_02373__PTR169) );
  MUX2_X1 U7762 ( .A(P2_P1_InstAddrPointer_PTR10), .B(_03055__PTR10), .S(_02146__PTR2), .Z(_02373__PTR170) );
  MUX2_X1 U7763 ( .A(P2_P1_InstAddrPointer_PTR11), .B(_03055__PTR11), .S(_02146__PTR2), .Z(_02373__PTR171) );
  MUX2_X1 U7764 ( .A(P2_P1_InstAddrPointer_PTR12), .B(_03055__PTR12), .S(_02146__PTR2), .Z(_02373__PTR172) );
  MUX2_X1 U7765 ( .A(P2_P1_InstAddrPointer_PTR13), .B(_03055__PTR13), .S(_02146__PTR2), .Z(_02373__PTR173) );
  MUX2_X1 U7766 ( .A(P2_P1_InstAddrPointer_PTR14), .B(_03055__PTR14), .S(_02146__PTR2), .Z(_02373__PTR174) );
  MUX2_X1 U7767 ( .A(P2_P1_InstAddrPointer_PTR15), .B(_03055__PTR15), .S(_02146__PTR2), .Z(_02373__PTR175) );
  MUX2_X1 U7768 ( .A(P2_P1_InstAddrPointer_PTR16), .B(_03055__PTR16), .S(_02146__PTR2), .Z(_02373__PTR176) );
  MUX2_X1 U7769 ( .A(P2_P1_InstAddrPointer_PTR17), .B(_03055__PTR17), .S(_02146__PTR2), .Z(_02373__PTR177) );
  MUX2_X1 U7770 ( .A(P2_P1_InstAddrPointer_PTR18), .B(_03055__PTR18), .S(_02146__PTR2), .Z(_02373__PTR178) );
  MUX2_X1 U7771 ( .A(P2_P1_InstAddrPointer_PTR19), .B(_03055__PTR19), .S(_02146__PTR2), .Z(_02373__PTR179) );
  MUX2_X1 U7772 ( .A(P2_P1_InstAddrPointer_PTR20), .B(_03055__PTR20), .S(_02146__PTR2), .Z(_02373__PTR180) );
  MUX2_X1 U7773 ( .A(P2_P1_InstAddrPointer_PTR21), .B(_03055__PTR21), .S(_02146__PTR2), .Z(_02373__PTR181) );
  MUX2_X1 U7774 ( .A(P2_P1_InstAddrPointer_PTR22), .B(_03055__PTR22), .S(_02146__PTR2), .Z(_02373__PTR182) );
  MUX2_X1 U7775 ( .A(P2_P1_InstAddrPointer_PTR23), .B(_03055__PTR23), .S(_02146__PTR2), .Z(_02373__PTR183) );
  MUX2_X1 U7776 ( .A(P2_P1_InstAddrPointer_PTR24), .B(_03055__PTR24), .S(_02146__PTR2), .Z(_02373__PTR184) );
  MUX2_X1 U7777 ( .A(P2_P1_InstAddrPointer_PTR25), .B(_03055__PTR25), .S(_02146__PTR2), .Z(_02373__PTR185) );
  MUX2_X1 U7778 ( .A(P2_P1_InstAddrPointer_PTR26), .B(_03055__PTR26), .S(_02146__PTR2), .Z(_02373__PTR186) );
  MUX2_X1 U7779 ( .A(P2_P1_InstAddrPointer_PTR27), .B(_03055__PTR27), .S(_02146__PTR2), .Z(_02373__PTR187) );
  MUX2_X1 U7780 ( .A(P2_P1_InstAddrPointer_PTR28), .B(_03055__PTR28), .S(_02146__PTR2), .Z(_02373__PTR188) );
  MUX2_X1 U7781 ( .A(P2_P1_InstAddrPointer_PTR29), .B(_03055__PTR29), .S(_02146__PTR2), .Z(_02373__PTR189) );
  MUX2_X1 U7782 ( .A(P2_P1_InstAddrPointer_PTR30), .B(_03055__PTR30), .S(_02146__PTR2), .Z(_02373__PTR190) );
  MUX2_X1 U7783 ( .A(P2_P1_InstAddrPointer_PTR31), .B(_03055__PTR31), .S(_02146__PTR2), .Z(_02373__PTR191) );
  MUX2_X1 U7784 ( .A(P2_rEIP_PTR0), .B(_02176__PTR3), .S(_02296_), .Z(_02393__PTR32) );
  MUX2_X1 U7785 ( .A(P2_rEIP_PTR1), .B(_02176__PTR4), .S(_02296_), .Z(_02393__PTR33) );
  MUX2_X1 U7786 ( .A(P2_rEIP_PTR2), .B(_02176__PTR5), .S(_02296_), .Z(_02393__PTR34) );
  MUX2_X1 U7787 ( .A(P2_rEIP_PTR3), .B(_02176__PTR6), .S(_02296_), .Z(_02393__PTR35) );
  MUX2_X1 U7788 ( .A(P2_rEIP_PTR4), .B(_03045__PTR4), .S(_02296_), .Z(_02393__PTR36) );
  MUX2_X1 U7789 ( .A(P2_rEIP_PTR5), .B(_03044__PTR4), .S(_02296_), .Z(_02393__PTR37) );
  MUX2_X1 U7790 ( .A(P2_rEIP_PTR6), .B(1'b0), .S(_02296_), .Z(_02393__PTR38) );
  MUX2_X1 U7791 ( .A(P2_rEIP_PTR7), .B(1'b0), .S(_02296_), .Z(_02393__PTR39) );
  MUX2_X1 U7792 ( .A(P2_rEIP_PTR8), .B(1'b0), .S(_02296_), .Z(_02393__PTR40) );
  MUX2_X1 U7793 ( .A(P2_rEIP_PTR9), .B(1'b0), .S(_02296_), .Z(_02393__PTR41) );
  MUX2_X1 U7794 ( .A(P2_rEIP_PTR10), .B(1'b0), .S(_02296_), .Z(_02393__PTR42) );
  MUX2_X1 U7795 ( .A(P2_rEIP_PTR11), .B(1'b0), .S(_02296_), .Z(_02393__PTR43) );
  MUX2_X1 U7796 ( .A(P2_rEIP_PTR12), .B(1'b0), .S(_02296_), .Z(_02393__PTR44) );
  MUX2_X1 U7797 ( .A(P2_rEIP_PTR13), .B(1'b0), .S(_02296_), .Z(_02393__PTR45) );
  MUX2_X1 U7798 ( .A(P2_rEIP_PTR14), .B(1'b0), .S(_02296_), .Z(_02393__PTR46) );
  MUX2_X1 U7799 ( .A(P2_rEIP_PTR15), .B(1'b0), .S(_02296_), .Z(_02393__PTR47) );
  MUX2_X1 U7800 ( .A(P2_rEIP_PTR16), .B(1'b0), .S(_02296_), .Z(_02393__PTR48) );
  MUX2_X1 U7801 ( .A(P2_rEIP_PTR17), .B(1'b0), .S(_02296_), .Z(_02393__PTR49) );
  MUX2_X1 U7802 ( .A(P2_rEIP_PTR18), .B(1'b0), .S(_02296_), .Z(_02393__PTR50) );
  MUX2_X1 U7803 ( .A(P2_rEIP_PTR19), .B(1'b0), .S(_02296_), .Z(_02393__PTR51) );
  MUX2_X1 U7804 ( .A(P2_rEIP_PTR20), .B(1'b0), .S(_02296_), .Z(_02393__PTR52) );
  MUX2_X1 U7805 ( .A(P2_rEIP_PTR21), .B(1'b0), .S(_02296_), .Z(_02393__PTR53) );
  MUX2_X1 U7806 ( .A(P2_rEIP_PTR22), .B(1'b0), .S(_02296_), .Z(_02393__PTR54) );
  MUX2_X1 U7807 ( .A(P2_rEIP_PTR23), .B(1'b0), .S(_02296_), .Z(_02393__PTR55) );
  MUX2_X1 U7808 ( .A(P2_rEIP_PTR24), .B(1'b0), .S(_02296_), .Z(_02393__PTR56) );
  MUX2_X1 U7809 ( .A(P2_rEIP_PTR25), .B(1'b0), .S(_02296_), .Z(_02393__PTR57) );
  MUX2_X1 U7810 ( .A(P2_rEIP_PTR26), .B(1'b0), .S(_02296_), .Z(_02393__PTR58) );
  MUX2_X1 U7811 ( .A(P2_rEIP_PTR27), .B(1'b0), .S(_02296_), .Z(_02393__PTR59) );
  MUX2_X1 U7812 ( .A(P2_rEIP_PTR28), .B(1'b0), .S(_02296_), .Z(_02393__PTR60) );
  MUX2_X1 U7813 ( .A(P2_rEIP_PTR29), .B(1'b0), .S(_02296_), .Z(_02393__PTR61) );
  MUX2_X1 U7814 ( .A(P2_rEIP_PTR30), .B(1'b0), .S(_02296_), .Z(_02393__PTR62) );
  MUX2_X1 U7815 ( .A(P2_rEIP_PTR31), .B(1'b0), .S(_02296_), .Z(_02393__PTR63) );
  MUX2_X1 U7816 ( .A(P2_rEIP_PTR0), .B(_02323__PTR0), .S(_02296_), .Z(_02393__PTR64) );
  MUX2_X1 U7817 ( .A(P2_rEIP_PTR1), .B(_02323__PTR1), .S(_02296_), .Z(_02393__PTR65) );
  MUX2_X1 U7818 ( .A(P2_rEIP_PTR2), .B(_02323__PTR2), .S(_02296_), .Z(_02393__PTR66) );
  MUX2_X1 U7819 ( .A(P2_rEIP_PTR3), .B(_02323__PTR3), .S(_02296_), .Z(_02393__PTR67) );
  MUX2_X1 U7820 ( .A(P2_rEIP_PTR4), .B(_02323__PTR4), .S(_02296_), .Z(_02393__PTR68) );
  MUX2_X1 U7821 ( .A(P2_rEIP_PTR5), .B(_02323__PTR5), .S(_02296_), .Z(_02393__PTR69) );
  MUX2_X1 U7822 ( .A(P2_rEIP_PTR6), .B(_02323__PTR6), .S(_02296_), .Z(_02393__PTR70) );
  MUX2_X1 U7823 ( .A(P2_rEIP_PTR7), .B(_02323__PTR7), .S(_02296_), .Z(_02393__PTR71) );
  MUX2_X1 U7824 ( .A(P2_rEIP_PTR8), .B(_02323__PTR8), .S(_02296_), .Z(_02393__PTR72) );
  MUX2_X1 U7825 ( .A(P2_rEIP_PTR9), .B(_02323__PTR9), .S(_02296_), .Z(_02393__PTR73) );
  MUX2_X1 U7826 ( .A(P2_rEIP_PTR10), .B(_02323__PTR10), .S(_02296_), .Z(_02393__PTR74) );
  MUX2_X1 U7827 ( .A(P2_rEIP_PTR11), .B(_02323__PTR11), .S(_02296_), .Z(_02393__PTR75) );
  MUX2_X1 U7828 ( .A(P2_rEIP_PTR12), .B(_02323__PTR12), .S(_02296_), .Z(_02393__PTR76) );
  MUX2_X1 U7829 ( .A(P2_rEIP_PTR13), .B(_02323__PTR13), .S(_02296_), .Z(_02393__PTR77) );
  MUX2_X1 U7830 ( .A(P2_rEIP_PTR14), .B(_02323__PTR14), .S(_02296_), .Z(_02393__PTR78) );
  MUX2_X1 U7831 ( .A(P2_rEIP_PTR15), .B(_02323__PTR15), .S(_02296_), .Z(_02393__PTR79) );
  MUX2_X1 U7832 ( .A(P2_rEIP_PTR16), .B(_02323__PTR16), .S(_02296_), .Z(_02393__PTR80) );
  MUX2_X1 U7833 ( .A(P2_rEIP_PTR17), .B(_02323__PTR17), .S(_02296_), .Z(_02393__PTR81) );
  MUX2_X1 U7834 ( .A(P2_rEIP_PTR18), .B(_02323__PTR18), .S(_02296_), .Z(_02393__PTR82) );
  MUX2_X1 U7835 ( .A(P2_rEIP_PTR19), .B(_02323__PTR19), .S(_02296_), .Z(_02393__PTR83) );
  MUX2_X1 U7836 ( .A(P2_rEIP_PTR20), .B(_02323__PTR20), .S(_02296_), .Z(_02393__PTR84) );
  MUX2_X1 U7837 ( .A(P2_rEIP_PTR21), .B(_02323__PTR21), .S(_02296_), .Z(_02393__PTR85) );
  MUX2_X1 U7838 ( .A(P2_rEIP_PTR22), .B(_02323__PTR22), .S(_02296_), .Z(_02393__PTR86) );
  MUX2_X1 U7839 ( .A(P2_rEIP_PTR23), .B(_02323__PTR23), .S(_02296_), .Z(_02393__PTR87) );
  MUX2_X1 U7840 ( .A(P2_rEIP_PTR24), .B(_02323__PTR24), .S(_02296_), .Z(_02393__PTR88) );
  MUX2_X1 U7841 ( .A(P2_rEIP_PTR25), .B(_02323__PTR25), .S(_02296_), .Z(_02393__PTR89) );
  MUX2_X1 U7842 ( .A(P2_rEIP_PTR26), .B(_02323__PTR26), .S(_02296_), .Z(_02393__PTR90) );
  MUX2_X1 U7843 ( .A(P2_rEIP_PTR27), .B(_02323__PTR27), .S(_02296_), .Z(_02393__PTR91) );
  MUX2_X1 U7844 ( .A(P2_rEIP_PTR28), .B(_02323__PTR28), .S(_02296_), .Z(_02393__PTR92) );
  MUX2_X1 U7845 ( .A(P2_rEIP_PTR29), .B(_02323__PTR29), .S(_02296_), .Z(_02393__PTR93) );
  MUX2_X1 U7846 ( .A(P2_rEIP_PTR30), .B(_02323__PTR30), .S(_02296_), .Z(_02393__PTR94) );
  MUX2_X1 U7847 ( .A(P2_rEIP_PTR31), .B(_02323__PTR31), .S(_02296_), .Z(_02393__PTR95) );
  MUX2_X1 U7848 ( .A(P2_rEIP_PTR0), .B(_02305__PTR0), .S(_02296_), .Z(_02393__PTR96) );
  MUX2_X1 U7849 ( .A(P2_rEIP_PTR1), .B(_02305__PTR1), .S(_02296_), .Z(_02393__PTR97) );
  MUX2_X1 U7850 ( .A(P2_rEIP_PTR2), .B(_02305__PTR2), .S(_02296_), .Z(_02393__PTR98) );
  MUX2_X1 U7851 ( .A(P2_rEIP_PTR3), .B(_02305__PTR3), .S(_02296_), .Z(_02393__PTR99) );
  MUX2_X1 U7852 ( .A(P2_rEIP_PTR4), .B(_02305__PTR4), .S(_02296_), .Z(_02393__PTR100) );
  MUX2_X1 U7853 ( .A(P2_rEIP_PTR5), .B(_02305__PTR5), .S(_02296_), .Z(_02393__PTR101) );
  MUX2_X1 U7854 ( .A(P2_rEIP_PTR6), .B(_02305__PTR6), .S(_02296_), .Z(_02393__PTR102) );
  MUX2_X1 U7855 ( .A(P2_rEIP_PTR7), .B(_02305__PTR7), .S(_02296_), .Z(_02393__PTR103) );
  MUX2_X1 U7856 ( .A(P2_rEIP_PTR8), .B(_02305__PTR8), .S(_02296_), .Z(_02393__PTR104) );
  MUX2_X1 U7857 ( .A(P2_rEIP_PTR9), .B(_02305__PTR9), .S(_02296_), .Z(_02393__PTR105) );
  MUX2_X1 U7858 ( .A(P2_rEIP_PTR10), .B(_02305__PTR10), .S(_02296_), .Z(_02393__PTR106) );
  MUX2_X1 U7859 ( .A(P2_rEIP_PTR11), .B(_02305__PTR11), .S(_02296_), .Z(_02393__PTR107) );
  MUX2_X1 U7860 ( .A(P2_rEIP_PTR12), .B(_02305__PTR12), .S(_02296_), .Z(_02393__PTR108) );
  MUX2_X1 U7861 ( .A(P2_rEIP_PTR13), .B(_02305__PTR13), .S(_02296_), .Z(_02393__PTR109) );
  MUX2_X1 U7862 ( .A(P2_rEIP_PTR14), .B(_02305__PTR14), .S(_02296_), .Z(_02393__PTR110) );
  MUX2_X1 U7863 ( .A(P2_rEIP_PTR15), .B(_02305__PTR15), .S(_02296_), .Z(_02393__PTR111) );
  MUX2_X1 U7864 ( .A(P2_rEIP_PTR16), .B(_02305__PTR16), .S(_02296_), .Z(_02393__PTR112) );
  MUX2_X1 U7865 ( .A(P2_rEIP_PTR17), .B(_02305__PTR17), .S(_02296_), .Z(_02393__PTR113) );
  MUX2_X1 U7866 ( .A(P2_rEIP_PTR18), .B(_02305__PTR18), .S(_02296_), .Z(_02393__PTR114) );
  MUX2_X1 U7867 ( .A(P2_rEIP_PTR19), .B(_02305__PTR19), .S(_02296_), .Z(_02393__PTR115) );
  MUX2_X1 U7868 ( .A(P2_rEIP_PTR20), .B(_02305__PTR20), .S(_02296_), .Z(_02393__PTR116) );
  MUX2_X1 U7869 ( .A(P2_rEIP_PTR21), .B(_02305__PTR21), .S(_02296_), .Z(_02393__PTR117) );
  MUX2_X1 U7870 ( .A(P2_rEIP_PTR22), .B(_02305__PTR22), .S(_02296_), .Z(_02393__PTR118) );
  MUX2_X1 U7871 ( .A(P2_rEIP_PTR23), .B(_02305__PTR23), .S(_02296_), .Z(_02393__PTR119) );
  MUX2_X1 U7872 ( .A(P2_rEIP_PTR24), .B(_02305__PTR24), .S(_02296_), .Z(_02393__PTR120) );
  MUX2_X1 U7873 ( .A(P2_rEIP_PTR25), .B(_02305__PTR25), .S(_02296_), .Z(_02393__PTR121) );
  MUX2_X1 U7874 ( .A(P2_rEIP_PTR26), .B(_02305__PTR26), .S(_02296_), .Z(_02393__PTR122) );
  MUX2_X1 U7875 ( .A(P2_rEIP_PTR27), .B(_02305__PTR27), .S(_02296_), .Z(_02393__PTR123) );
  MUX2_X1 U7876 ( .A(P2_rEIP_PTR28), .B(_02305__PTR28), .S(_02296_), .Z(_02393__PTR124) );
  MUX2_X1 U7877 ( .A(P2_rEIP_PTR29), .B(_02305__PTR29), .S(_02296_), .Z(_02393__PTR125) );
  MUX2_X1 U7878 ( .A(P2_rEIP_PTR30), .B(_02305__PTR30), .S(_02296_), .Z(_02393__PTR126) );
  MUX2_X1 U7879 ( .A(P2_rEIP_PTR31), .B(_02305__PTR31), .S(_02296_), .Z(_02393__PTR127) );
  MUX2_X1 U7880 ( .A(P2_rEIP_PTR0), .B(P2_EBX_PTR0), .S(P2_StateBS16), .Z(_02300__PTR0) );
  MUX2_X1 U7881 ( .A(_02174__PTR7), .B(_02299__PTR1), .S(P2_StateBS16), .Z(_02300__PTR1) );
  MUX2_X1 U7882 ( .A(_03067__PTR1), .B(_02299__PTR2), .S(P2_StateBS16), .Z(_02300__PTR2) );
  MUX2_X1 U7883 ( .A(_03067__PTR2), .B(_02299__PTR3), .S(P2_StateBS16), .Z(_02300__PTR3) );
  MUX2_X1 U7884 ( .A(_03067__PTR3), .B(_02299__PTR4), .S(P2_StateBS16), .Z(_02300__PTR4) );
  MUX2_X1 U7885 ( .A(_03067__PTR4), .B(_02299__PTR5), .S(P2_StateBS16), .Z(_02300__PTR5) );
  MUX2_X1 U7886 ( .A(_03067__PTR5), .B(_02299__PTR6), .S(P2_StateBS16), .Z(_02300__PTR6) );
  MUX2_X1 U7887 ( .A(_03067__PTR6), .B(_02299__PTR7), .S(P2_StateBS16), .Z(_02300__PTR7) );
  MUX2_X1 U7888 ( .A(_03067__PTR7), .B(_02299__PTR8), .S(P2_StateBS16), .Z(_02300__PTR8) );
  MUX2_X1 U7889 ( .A(_03067__PTR8), .B(_02299__PTR9), .S(P2_StateBS16), .Z(_02300__PTR9) );
  MUX2_X1 U7890 ( .A(_03067__PTR9), .B(_02299__PTR10), .S(P2_StateBS16), .Z(_02300__PTR10) );
  MUX2_X1 U7891 ( .A(_03067__PTR10), .B(_02299__PTR11), .S(P2_StateBS16), .Z(_02300__PTR11) );
  MUX2_X1 U7892 ( .A(_03067__PTR11), .B(_02299__PTR12), .S(P2_StateBS16), .Z(_02300__PTR12) );
  MUX2_X1 U7893 ( .A(_03067__PTR12), .B(_02299__PTR13), .S(P2_StateBS16), .Z(_02300__PTR13) );
  MUX2_X1 U7894 ( .A(_03067__PTR13), .B(_02299__PTR14), .S(P2_StateBS16), .Z(_02300__PTR14) );
  MUX2_X1 U7895 ( .A(_03067__PTR14), .B(_02299__PTR15), .S(P2_StateBS16), .Z(_02300__PTR15) );
  MUX2_X1 U7896 ( .A(_03067__PTR15), .B(_02299__PTR16), .S(P2_StateBS16), .Z(_02300__PTR16) );
  MUX2_X1 U7897 ( .A(_03067__PTR16), .B(_02299__PTR17), .S(P2_StateBS16), .Z(_02300__PTR17) );
  MUX2_X1 U7898 ( .A(_03067__PTR17), .B(_02299__PTR18), .S(P2_StateBS16), .Z(_02300__PTR18) );
  MUX2_X1 U7899 ( .A(_03067__PTR18), .B(_02299__PTR19), .S(P2_StateBS16), .Z(_02300__PTR19) );
  MUX2_X1 U7900 ( .A(_03067__PTR19), .B(_02299__PTR20), .S(P2_StateBS16), .Z(_02300__PTR20) );
  MUX2_X1 U7901 ( .A(_03067__PTR20), .B(_02299__PTR21), .S(P2_StateBS16), .Z(_02300__PTR21) );
  MUX2_X1 U7902 ( .A(_03067__PTR21), .B(_02299__PTR22), .S(P2_StateBS16), .Z(_02300__PTR22) );
  MUX2_X1 U7903 ( .A(_03067__PTR22), .B(_02299__PTR23), .S(P2_StateBS16), .Z(_02300__PTR23) );
  MUX2_X1 U7904 ( .A(_03067__PTR23), .B(_02299__PTR24), .S(P2_StateBS16), .Z(_02300__PTR24) );
  MUX2_X1 U7905 ( .A(_03067__PTR24), .B(_02299__PTR25), .S(P2_StateBS16), .Z(_02300__PTR25) );
  MUX2_X1 U7906 ( .A(_03067__PTR25), .B(_02299__PTR26), .S(P2_StateBS16), .Z(_02300__PTR26) );
  MUX2_X1 U7907 ( .A(_03067__PTR26), .B(_02299__PTR27), .S(P2_StateBS16), .Z(_02300__PTR27) );
  MUX2_X1 U7908 ( .A(_03067__PTR27), .B(_02299__PTR28), .S(P2_StateBS16), .Z(_02300__PTR28) );
  MUX2_X1 U7909 ( .A(_03067__PTR28), .B(_02299__PTR29), .S(P2_StateBS16), .Z(_02300__PTR29) );
  MUX2_X1 U7910 ( .A(_03067__PTR29), .B(_02299__PTR30), .S(P2_StateBS16), .Z(_02300__PTR30) );
  MUX2_X1 U7911 ( .A(_03067__PTR30), .B(_02299__PTR31), .S(P2_StateBS16), .Z(_02300__PTR31) );
  MUX2_X1 U7912 ( .A(_03193__PTR1), .B(P2_EBX_PTR1), .S(_02978__PTR31), .Z(_02299__PTR1) );
  MUX2_X1 U7913 ( .A(_03193__PTR2), .B(P2_EBX_PTR2), .S(_02978__PTR31), .Z(_02299__PTR2) );
  MUX2_X1 U7914 ( .A(_03193__PTR3), .B(P2_EBX_PTR3), .S(_02978__PTR31), .Z(_02299__PTR3) );
  MUX2_X1 U7915 ( .A(_03193__PTR4), .B(P2_EBX_PTR4), .S(_02978__PTR31), .Z(_02299__PTR4) );
  MUX2_X1 U7916 ( .A(_03193__PTR5), .B(P2_EBX_PTR5), .S(_02978__PTR31), .Z(_02299__PTR5) );
  MUX2_X1 U7917 ( .A(_03193__PTR6), .B(P2_EBX_PTR6), .S(_02978__PTR31), .Z(_02299__PTR6) );
  MUX2_X1 U7918 ( .A(_03193__PTR7), .B(P2_EBX_PTR7), .S(_02978__PTR31), .Z(_02299__PTR7) );
  MUX2_X1 U7919 ( .A(_03193__PTR8), .B(P2_EBX_PTR8), .S(_02978__PTR31), .Z(_02299__PTR8) );
  MUX2_X1 U7920 ( .A(_03193__PTR9), .B(P2_EBX_PTR9), .S(_02978__PTR31), .Z(_02299__PTR9) );
  MUX2_X1 U7921 ( .A(_03193__PTR10), .B(P2_EBX_PTR10), .S(_02978__PTR31), .Z(_02299__PTR10) );
  MUX2_X1 U7922 ( .A(_03193__PTR11), .B(P2_EBX_PTR11), .S(_02978__PTR31), .Z(_02299__PTR11) );
  MUX2_X1 U7923 ( .A(_03193__PTR12), .B(P2_EBX_PTR12), .S(_02978__PTR31), .Z(_02299__PTR12) );
  MUX2_X1 U7924 ( .A(_03193__PTR13), .B(P2_EBX_PTR13), .S(_02978__PTR31), .Z(_02299__PTR13) );
  MUX2_X1 U7925 ( .A(_03193__PTR14), .B(P2_EBX_PTR14), .S(_02978__PTR31), .Z(_02299__PTR14) );
  MUX2_X1 U7926 ( .A(_03193__PTR15), .B(P2_EBX_PTR15), .S(_02978__PTR31), .Z(_02299__PTR15) );
  MUX2_X1 U7927 ( .A(_03193__PTR16), .B(P2_EBX_PTR16), .S(_02978__PTR31), .Z(_02299__PTR16) );
  MUX2_X1 U7928 ( .A(_03193__PTR17), .B(P2_EBX_PTR17), .S(_02978__PTR31), .Z(_02299__PTR17) );
  MUX2_X1 U7929 ( .A(_03193__PTR18), .B(P2_EBX_PTR18), .S(_02978__PTR31), .Z(_02299__PTR18) );
  MUX2_X1 U7930 ( .A(_03193__PTR19), .B(P2_EBX_PTR19), .S(_02978__PTR31), .Z(_02299__PTR19) );
  MUX2_X1 U7931 ( .A(_03193__PTR20), .B(P2_EBX_PTR20), .S(_02978__PTR31), .Z(_02299__PTR20) );
  MUX2_X1 U7932 ( .A(_03193__PTR21), .B(P2_EBX_PTR21), .S(_02978__PTR31), .Z(_02299__PTR21) );
  MUX2_X1 U7933 ( .A(_03193__PTR22), .B(P2_EBX_PTR22), .S(_02978__PTR31), .Z(_02299__PTR22) );
  MUX2_X1 U7934 ( .A(_03193__PTR23), .B(P2_EBX_PTR23), .S(_02978__PTR31), .Z(_02299__PTR23) );
  MUX2_X1 U7935 ( .A(_03193__PTR24), .B(P2_EBX_PTR24), .S(_02978__PTR31), .Z(_02299__PTR24) );
  MUX2_X1 U7936 ( .A(_03193__PTR25), .B(P2_EBX_PTR25), .S(_02978__PTR31), .Z(_02299__PTR25) );
  MUX2_X1 U7937 ( .A(_03193__PTR26), .B(P2_EBX_PTR26), .S(_02978__PTR31), .Z(_02299__PTR26) );
  MUX2_X1 U7938 ( .A(_03193__PTR27), .B(P2_EBX_PTR27), .S(_02978__PTR31), .Z(_02299__PTR27) );
  MUX2_X1 U7939 ( .A(_03193__PTR28), .B(P2_EBX_PTR28), .S(_02978__PTR31), .Z(_02299__PTR28) );
  MUX2_X1 U7940 ( .A(_03193__PTR29), .B(P2_EBX_PTR29), .S(_02978__PTR31), .Z(_02299__PTR29) );
  MUX2_X1 U7941 ( .A(_03193__PTR30), .B(P2_EBX_PTR30), .S(_02978__PTR31), .Z(_02299__PTR30) );
  MUX2_X1 U7942 ( .A(_03193__PTR31), .B(P2_EBX_PTR31), .S(_02978__PTR31), .Z(_02299__PTR31) );
  MUX2_X1 U7943 ( .A(P2_EBX_PTR0), .B(P2_P1_InstQueue_PTR0_PTR0), .S(_02146__PTR2), .Z(_02389__PTR64) );
  MUX2_X1 U7944 ( .A(P2_EBX_PTR1), .B(P2_P1_InstQueue_PTR0_PTR1), .S(_02146__PTR2), .Z(_02389__PTR65) );
  MUX2_X1 U7945 ( .A(P2_EBX_PTR2), .B(P2_P1_InstQueue_PTR0_PTR2), .S(_02146__PTR2), .Z(_02389__PTR66) );
  MUX2_X1 U7946 ( .A(P2_EBX_PTR3), .B(P2_P1_InstQueue_PTR0_PTR3), .S(_02146__PTR2), .Z(_02389__PTR67) );
  MUX2_X1 U7947 ( .A(P2_EBX_PTR4), .B(P2_P1_InstQueue_PTR0_PTR4), .S(_02146__PTR2), .Z(_02389__PTR68) );
  MUX2_X1 U7948 ( .A(P2_EBX_PTR5), .B(P2_P1_InstQueue_PTR0_PTR5), .S(_02146__PTR2), .Z(_02389__PTR69) );
  MUX2_X1 U7949 ( .A(P2_EBX_PTR6), .B(P2_P1_InstQueue_PTR0_PTR6), .S(_02146__PTR2), .Z(_02389__PTR70) );
  MUX2_X1 U7950 ( .A(P2_EBX_PTR7), .B(P2_P1_InstQueue_PTR0_PTR7), .S(_02146__PTR2), .Z(_02389__PTR71) );
  MUX2_X1 U7951 ( .A(P2_EBX_PTR8), .B(_02183__PTR0), .S(_02146__PTR2), .Z(_02389__PTR72) );
  MUX2_X1 U7952 ( .A(P2_EBX_PTR9), .B(_02183__PTR1), .S(_02146__PTR2), .Z(_02389__PTR73) );
  MUX2_X1 U7953 ( .A(P2_EBX_PTR10), .B(_02183__PTR2), .S(_02146__PTR2), .Z(_02389__PTR74) );
  MUX2_X1 U7954 ( .A(P2_EBX_PTR11), .B(_02183__PTR3), .S(_02146__PTR2), .Z(_02389__PTR75) );
  MUX2_X1 U7955 ( .A(P2_EBX_PTR12), .B(_02183__PTR4), .S(_02146__PTR2), .Z(_02389__PTR76) );
  MUX2_X1 U7956 ( .A(P2_EBX_PTR13), .B(_02183__PTR5), .S(_02146__PTR2), .Z(_02389__PTR77) );
  MUX2_X1 U7957 ( .A(P2_EBX_PTR14), .B(_02183__PTR6), .S(_02146__PTR2), .Z(_02389__PTR78) );
  MUX2_X1 U7958 ( .A(P2_EBX_PTR15), .B(_02183__PTR7), .S(_02146__PTR2), .Z(_02389__PTR79) );
  MUX2_X1 U7959 ( .A(P2_EBX_PTR16), .B(_02181__PTR0), .S(_02146__PTR2), .Z(_02389__PTR80) );
  MUX2_X1 U7960 ( .A(P2_EBX_PTR17), .B(_02181__PTR1), .S(_02146__PTR2), .Z(_02389__PTR81) );
  MUX2_X1 U7961 ( .A(P2_EBX_PTR18), .B(_02181__PTR2), .S(_02146__PTR2), .Z(_02389__PTR82) );
  MUX2_X1 U7962 ( .A(P2_EBX_PTR19), .B(_02181__PTR3), .S(_02146__PTR2), .Z(_02389__PTR83) );
  MUX2_X1 U7963 ( .A(P2_EBX_PTR20), .B(_02181__PTR4), .S(_02146__PTR2), .Z(_02389__PTR84) );
  MUX2_X1 U7964 ( .A(P2_EBX_PTR21), .B(_02181__PTR5), .S(_02146__PTR2), .Z(_02389__PTR85) );
  MUX2_X1 U7965 ( .A(P2_EBX_PTR22), .B(_02181__PTR6), .S(_02146__PTR2), .Z(_02389__PTR86) );
  MUX2_X1 U7966 ( .A(P2_EBX_PTR23), .B(_03060__PTR0), .S(_02146__PTR2), .Z(_02389__PTR87) );
  MUX2_X1 U7967 ( .A(P2_EBX_PTR24), .B(_03061__PTR1), .S(_02146__PTR2), .Z(_02389__PTR88) );
  MUX2_X1 U7968 ( .A(P2_EBX_PTR25), .B(_03061__PTR2), .S(_02146__PTR2), .Z(_02389__PTR89) );
  MUX2_X1 U7969 ( .A(P2_EBX_PTR26), .B(_03061__PTR3), .S(_02146__PTR2), .Z(_02389__PTR90) );
  MUX2_X1 U7970 ( .A(P2_EBX_PTR27), .B(_03061__PTR4), .S(_02146__PTR2), .Z(_02389__PTR91) );
  MUX2_X1 U7971 ( .A(P2_EBX_PTR28), .B(_03061__PTR5), .S(_02146__PTR2), .Z(_02389__PTR92) );
  MUX2_X1 U7972 ( .A(P2_EBX_PTR29), .B(_03061__PTR6), .S(_02146__PTR2), .Z(_02389__PTR93) );
  MUX2_X1 U7973 ( .A(P2_EBX_PTR30), .B(_03061__PTR7), .S(_02146__PTR2), .Z(_02389__PTR94) );
  MUX2_X1 U7974 ( .A(P2_EBX_PTR31), .B(_03059__PTR7), .S(_02146__PTR2), .Z(_02389__PTR95) );
  MUX2_X1 U7975 ( .A(P2_P1_InstQueueRd_Addr_PTR0), .B(_02176__PTR3), .S(_02146__PTR2), .Z(_02377__PTR25) );
  MUX2_X1 U7976 ( .A(P2_P1_InstQueueRd_Addr_PTR1), .B(_02176__PTR4), .S(_02146__PTR2), .Z(_02377__PTR26) );
  MUX2_X1 U7977 ( .A(P2_P1_InstQueueRd_Addr_PTR2), .B(_03065__PTR2), .S(_02146__PTR2), .Z(_02377__PTR27) );
  MUX2_X1 U7978 ( .A(P2_P1_InstQueueRd_Addr_PTR3), .B(_03065__PTR3), .S(_02146__PTR2), .Z(_02377__PTR28) );
  MUX2_X1 U7979 ( .A(P2_P1_InstQueueRd_Addr_PTR4), .B(1'b0), .S(_02146__PTR2), .Z(_02377__PTR29) );
  MUX2_X1 U7980 ( .A(P2_EAX_PTR0), .B(_02177__PTR0), .S(_02146__PTR2), .Z(_02385__PTR128) );
  MUX2_X1 U7981 ( .A(P2_EAX_PTR1), .B(_02177__PTR1), .S(_02146__PTR2), .Z(_02385__PTR129) );
  MUX2_X1 U7982 ( .A(P2_EAX_PTR2), .B(_02177__PTR2), .S(_02146__PTR2), .Z(_02385__PTR130) );
  MUX2_X1 U7983 ( .A(P2_EAX_PTR3), .B(_02177__PTR3), .S(_02146__PTR2), .Z(_02385__PTR131) );
  MUX2_X1 U7984 ( .A(P2_EAX_PTR4), .B(_02177__PTR4), .S(_02146__PTR2), .Z(_02385__PTR132) );
  MUX2_X1 U7985 ( .A(P2_EAX_PTR5), .B(_02177__PTR5), .S(_02146__PTR2), .Z(_02385__PTR133) );
  MUX2_X1 U7986 ( .A(P2_EAX_PTR6), .B(_02177__PTR6), .S(_02146__PTR2), .Z(_02385__PTR134) );
  MUX2_X1 U7987 ( .A(P2_EAX_PTR7), .B(_02177__PTR7), .S(_02146__PTR2), .Z(_02385__PTR135) );
  MUX2_X1 U7988 ( .A(P2_EAX_PTR8), .B(_02183__PTR0), .S(_02146__PTR2), .Z(_02385__PTR136) );
  MUX2_X1 U7989 ( .A(P2_EAX_PTR9), .B(_02183__PTR1), .S(_02146__PTR2), .Z(_02385__PTR137) );
  MUX2_X1 U7990 ( .A(P2_EAX_PTR10), .B(_02183__PTR2), .S(_02146__PTR2), .Z(_02385__PTR138) );
  MUX2_X1 U7991 ( .A(P2_EAX_PTR11), .B(_02183__PTR3), .S(_02146__PTR2), .Z(_02385__PTR139) );
  MUX2_X1 U7992 ( .A(P2_EAX_PTR12), .B(_02183__PTR4), .S(_02146__PTR2), .Z(_02385__PTR140) );
  MUX2_X1 U7993 ( .A(P2_EAX_PTR13), .B(_02183__PTR5), .S(_02146__PTR2), .Z(_02385__PTR141) );
  MUX2_X1 U7994 ( .A(P2_EAX_PTR14), .B(_02183__PTR6), .S(_02146__PTR2), .Z(_02385__PTR142) );
  MUX2_X1 U7995 ( .A(P2_EAX_PTR15), .B(_02183__PTR7), .S(_02146__PTR2), .Z(_02385__PTR143) );
  MUX2_X1 U7996 ( .A(P2_EAX_PTR16), .B(_02181__PTR0), .S(_02146__PTR2), .Z(_02385__PTR144) );
  MUX2_X1 U7997 ( .A(P2_EAX_PTR17), .B(_02181__PTR1), .S(_02146__PTR2), .Z(_02385__PTR145) );
  MUX2_X1 U7998 ( .A(P2_EAX_PTR18), .B(_02181__PTR2), .S(_02146__PTR2), .Z(_02385__PTR146) );
  MUX2_X1 U7999 ( .A(P2_EAX_PTR19), .B(_02181__PTR3), .S(_02146__PTR2), .Z(_02385__PTR147) );
  MUX2_X1 U8000 ( .A(P2_EAX_PTR20), .B(_02181__PTR4), .S(_02146__PTR2), .Z(_02385__PTR148) );
  MUX2_X1 U8001 ( .A(P2_EAX_PTR21), .B(_02181__PTR5), .S(_02146__PTR2), .Z(_02385__PTR149) );
  MUX2_X1 U8002 ( .A(P2_EAX_PTR22), .B(_02181__PTR6), .S(_02146__PTR2), .Z(_02385__PTR150) );
  MUX2_X1 U8003 ( .A(P2_EAX_PTR23), .B(_03060__PTR0), .S(_02146__PTR2), .Z(_02385__PTR151) );
  MUX2_X1 U8004 ( .A(P2_EAX_PTR24), .B(_03061__PTR1), .S(_02146__PTR2), .Z(_02385__PTR152) );
  MUX2_X1 U8005 ( .A(P2_EAX_PTR25), .B(_03061__PTR2), .S(_02146__PTR2), .Z(_02385__PTR153) );
  MUX2_X1 U8006 ( .A(P2_EAX_PTR26), .B(_03061__PTR3), .S(_02146__PTR2), .Z(_02385__PTR154) );
  MUX2_X1 U8007 ( .A(P2_EAX_PTR27), .B(_03061__PTR4), .S(_02146__PTR2), .Z(_02385__PTR155) );
  MUX2_X1 U8008 ( .A(P2_EAX_PTR28), .B(_03061__PTR5), .S(_02146__PTR2), .Z(_02385__PTR156) );
  MUX2_X1 U8009 ( .A(P2_EAX_PTR29), .B(_03061__PTR6), .S(_02146__PTR2), .Z(_02385__PTR157) );
  MUX2_X1 U8010 ( .A(P2_EAX_PTR30), .B(_03061__PTR7), .S(_02146__PTR2), .Z(_02385__PTR158) );
  MUX2_X1 U8011 ( .A(P2_EAX_PTR31), .B(_03059__PTR7), .S(_02146__PTR2), .Z(_02385__PTR159) );
  MUX2_X1 U8012 ( .A(P2_P1_PhyAddrPointer_PTR0), .B(_03054__PTR0), .S(_02146__PTR2), .Z(_02381__PTR32) );
  MUX2_X1 U8013 ( .A(P2_P1_PhyAddrPointer_PTR1), .B(_03055__PTR1), .S(_02146__PTR2), .Z(_02381__PTR33) );
  MUX2_X1 U8014 ( .A(P2_P1_PhyAddrPointer_PTR2), .B(_03055__PTR2), .S(_02146__PTR2), .Z(_02381__PTR34) );
  MUX2_X1 U8015 ( .A(P2_P1_PhyAddrPointer_PTR3), .B(_03055__PTR3), .S(_02146__PTR2), .Z(_02381__PTR35) );
  MUX2_X1 U8016 ( .A(P2_P1_PhyAddrPointer_PTR4), .B(_03055__PTR4), .S(_02146__PTR2), .Z(_02381__PTR36) );
  MUX2_X1 U8017 ( .A(P2_P1_PhyAddrPointer_PTR5), .B(_03055__PTR5), .S(_02146__PTR2), .Z(_02381__PTR37) );
  MUX2_X1 U8018 ( .A(P2_P1_PhyAddrPointer_PTR6), .B(_03055__PTR6), .S(_02146__PTR2), .Z(_02381__PTR38) );
  MUX2_X1 U8019 ( .A(P2_P1_PhyAddrPointer_PTR7), .B(_03055__PTR7), .S(_02146__PTR2), .Z(_02381__PTR39) );
  MUX2_X1 U8020 ( .A(P2_P1_PhyAddrPointer_PTR8), .B(_03055__PTR8), .S(_02146__PTR2), .Z(_02381__PTR40) );
  MUX2_X1 U8021 ( .A(P2_P1_PhyAddrPointer_PTR9), .B(_03055__PTR9), .S(_02146__PTR2), .Z(_02381__PTR41) );
  MUX2_X1 U8022 ( .A(P2_P1_PhyAddrPointer_PTR10), .B(_03055__PTR10), .S(_02146__PTR2), .Z(_02381__PTR42) );
  MUX2_X1 U8023 ( .A(P2_P1_PhyAddrPointer_PTR11), .B(_03055__PTR11), .S(_02146__PTR2), .Z(_02381__PTR43) );
  MUX2_X1 U8024 ( .A(P2_P1_PhyAddrPointer_PTR12), .B(_03055__PTR12), .S(_02146__PTR2), .Z(_02381__PTR44) );
  MUX2_X1 U8025 ( .A(P2_P1_PhyAddrPointer_PTR13), .B(_03055__PTR13), .S(_02146__PTR2), .Z(_02381__PTR45) );
  MUX2_X1 U8026 ( .A(P2_P1_PhyAddrPointer_PTR14), .B(_03055__PTR14), .S(_02146__PTR2), .Z(_02381__PTR46) );
  MUX2_X1 U8027 ( .A(P2_P1_PhyAddrPointer_PTR15), .B(_03055__PTR15), .S(_02146__PTR2), .Z(_02381__PTR47) );
  MUX2_X1 U8028 ( .A(P2_P1_PhyAddrPointer_PTR16), .B(_03055__PTR16), .S(_02146__PTR2), .Z(_02381__PTR48) );
  MUX2_X1 U8029 ( .A(P2_P1_PhyAddrPointer_PTR17), .B(_03055__PTR17), .S(_02146__PTR2), .Z(_02381__PTR49) );
  MUX2_X1 U8030 ( .A(P2_P1_PhyAddrPointer_PTR18), .B(_03055__PTR18), .S(_02146__PTR2), .Z(_02381__PTR50) );
  MUX2_X1 U8031 ( .A(P2_P1_PhyAddrPointer_PTR19), .B(_03055__PTR19), .S(_02146__PTR2), .Z(_02381__PTR51) );
  MUX2_X1 U8032 ( .A(P2_P1_PhyAddrPointer_PTR20), .B(_03055__PTR20), .S(_02146__PTR2), .Z(_02381__PTR52) );
  MUX2_X1 U8033 ( .A(P2_P1_PhyAddrPointer_PTR21), .B(_03055__PTR21), .S(_02146__PTR2), .Z(_02381__PTR53) );
  MUX2_X1 U8034 ( .A(P2_P1_PhyAddrPointer_PTR22), .B(_03055__PTR22), .S(_02146__PTR2), .Z(_02381__PTR54) );
  MUX2_X1 U8035 ( .A(P2_P1_PhyAddrPointer_PTR23), .B(_03055__PTR23), .S(_02146__PTR2), .Z(_02381__PTR55) );
  MUX2_X1 U8036 ( .A(P2_P1_PhyAddrPointer_PTR24), .B(_03055__PTR24), .S(_02146__PTR2), .Z(_02381__PTR56) );
  MUX2_X1 U8037 ( .A(P2_P1_PhyAddrPointer_PTR25), .B(_03055__PTR25), .S(_02146__PTR2), .Z(_02381__PTR57) );
  MUX2_X1 U8038 ( .A(P2_P1_PhyAddrPointer_PTR26), .B(_03055__PTR26), .S(_02146__PTR2), .Z(_02381__PTR58) );
  MUX2_X1 U8039 ( .A(P2_P1_PhyAddrPointer_PTR27), .B(_03055__PTR27), .S(_02146__PTR2), .Z(_02381__PTR59) );
  MUX2_X1 U8040 ( .A(P2_P1_PhyAddrPointer_PTR28), .B(_03055__PTR28), .S(_02146__PTR2), .Z(_02381__PTR60) );
  MUX2_X1 U8041 ( .A(P2_P1_PhyAddrPointer_PTR29), .B(_03055__PTR29), .S(_02146__PTR2), .Z(_02381__PTR61) );
  MUX2_X1 U8042 ( .A(P2_P1_PhyAddrPointer_PTR30), .B(_03055__PTR30), .S(_02146__PTR2), .Z(_02381__PTR62) );
  MUX2_X1 U8043 ( .A(P2_P1_PhyAddrPointer_PTR31), .B(_03055__PTR31), .S(_02146__PTR2), .Z(_02381__PTR63) );
  MUX2_X1 U8044 ( .A(P2_P1_InstAddrPointer_PTR1), .B(_02327__PTR1), .S(_02296_), .Z(_02373__PTR65) );
  MUX2_X1 U8045 ( .A(P2_P1_InstAddrPointer_PTR2), .B(_02327__PTR2), .S(_02296_), .Z(_02373__PTR66) );
  MUX2_X1 U8046 ( .A(P2_P1_InstAddrPointer_PTR3), .B(_02327__PTR3), .S(_02296_), .Z(_02373__PTR67) );
  MUX2_X1 U8047 ( .A(P2_P1_InstAddrPointer_PTR4), .B(_02327__PTR4), .S(_02296_), .Z(_02373__PTR68) );
  MUX2_X1 U8048 ( .A(P2_P1_InstAddrPointer_PTR5), .B(_02327__PTR5), .S(_02296_), .Z(_02373__PTR69) );
  MUX2_X1 U8049 ( .A(P2_P1_InstAddrPointer_PTR6), .B(_02327__PTR6), .S(_02296_), .Z(_02373__PTR70) );
  MUX2_X1 U8050 ( .A(P2_P1_InstAddrPointer_PTR7), .B(_02327__PTR7), .S(_02296_), .Z(_02373__PTR71) );
  MUX2_X1 U8051 ( .A(P2_P1_InstAddrPointer_PTR8), .B(_02327__PTR8), .S(_02296_), .Z(_02373__PTR72) );
  MUX2_X1 U8052 ( .A(P2_P1_InstAddrPointer_PTR9), .B(_02327__PTR9), .S(_02296_), .Z(_02373__PTR73) );
  MUX2_X1 U8053 ( .A(P2_P1_InstAddrPointer_PTR10), .B(_02327__PTR10), .S(_02296_), .Z(_02373__PTR74) );
  MUX2_X1 U8054 ( .A(P2_P1_InstAddrPointer_PTR11), .B(_02327__PTR11), .S(_02296_), .Z(_02373__PTR75) );
  MUX2_X1 U8055 ( .A(P2_P1_InstAddrPointer_PTR12), .B(_02327__PTR12), .S(_02296_), .Z(_02373__PTR76) );
  MUX2_X1 U8056 ( .A(P2_P1_InstAddrPointer_PTR13), .B(_02327__PTR13), .S(_02296_), .Z(_02373__PTR77) );
  MUX2_X1 U8057 ( .A(P2_P1_InstAddrPointer_PTR14), .B(_02327__PTR14), .S(_02296_), .Z(_02373__PTR78) );
  MUX2_X1 U8058 ( .A(P2_P1_InstAddrPointer_PTR15), .B(_02327__PTR15), .S(_02296_), .Z(_02373__PTR79) );
  MUX2_X1 U8059 ( .A(P2_P1_InstAddrPointer_PTR16), .B(_02327__PTR16), .S(_02296_), .Z(_02373__PTR80) );
  MUX2_X1 U8060 ( .A(P2_P1_InstAddrPointer_PTR17), .B(_02327__PTR17), .S(_02296_), .Z(_02373__PTR81) );
  MUX2_X1 U8061 ( .A(P2_P1_InstAddrPointer_PTR18), .B(_02327__PTR18), .S(_02296_), .Z(_02373__PTR82) );
  MUX2_X1 U8062 ( .A(P2_P1_InstAddrPointer_PTR19), .B(_02327__PTR19), .S(_02296_), .Z(_02373__PTR83) );
  MUX2_X1 U8063 ( .A(P2_P1_InstAddrPointer_PTR20), .B(_02327__PTR20), .S(_02296_), .Z(_02373__PTR84) );
  MUX2_X1 U8064 ( .A(P2_P1_InstAddrPointer_PTR21), .B(_02327__PTR21), .S(_02296_), .Z(_02373__PTR85) );
  MUX2_X1 U8065 ( .A(P2_P1_InstAddrPointer_PTR22), .B(_02327__PTR22), .S(_02296_), .Z(_02373__PTR86) );
  MUX2_X1 U8066 ( .A(P2_P1_InstAddrPointer_PTR23), .B(_02327__PTR23), .S(_02296_), .Z(_02373__PTR87) );
  MUX2_X1 U8067 ( .A(P2_P1_InstAddrPointer_PTR24), .B(_02327__PTR24), .S(_02296_), .Z(_02373__PTR88) );
  MUX2_X1 U8068 ( .A(P2_P1_InstAddrPointer_PTR25), .B(_02327__PTR25), .S(_02296_), .Z(_02373__PTR89) );
  MUX2_X1 U8069 ( .A(P2_P1_InstAddrPointer_PTR26), .B(_02327__PTR26), .S(_02296_), .Z(_02373__PTR90) );
  MUX2_X1 U8070 ( .A(P2_P1_InstAddrPointer_PTR27), .B(_02327__PTR27), .S(_02296_), .Z(_02373__PTR91) );
  MUX2_X1 U8071 ( .A(P2_P1_InstAddrPointer_PTR28), .B(_02327__PTR28), .S(_02296_), .Z(_02373__PTR92) );
  MUX2_X1 U8072 ( .A(P2_P1_InstAddrPointer_PTR29), .B(_02327__PTR29), .S(_02296_), .Z(_02373__PTR93) );
  MUX2_X1 U8073 ( .A(P2_P1_InstAddrPointer_PTR30), .B(_02327__PTR30), .S(_02296_), .Z(_02373__PTR94) );
  MUX2_X1 U8074 ( .A(P2_P1_InstAddrPointer_PTR31), .B(_02327__PTR31), .S(_02296_), .Z(_02373__PTR95) );
  MUX2_X1 U8075 ( .A(P2_P1_InstAddrPointer_PTR1), .B(_02309__PTR1), .S(_02296_), .Z(_02373__PTR97) );
  MUX2_X1 U8076 ( .A(P2_P1_InstAddrPointer_PTR2), .B(_02309__PTR2), .S(_02296_), .Z(_02373__PTR98) );
  MUX2_X1 U8077 ( .A(P2_P1_InstAddrPointer_PTR3), .B(_02309__PTR3), .S(_02296_), .Z(_02373__PTR99) );
  MUX2_X1 U8078 ( .A(P2_P1_InstAddrPointer_PTR4), .B(_02309__PTR4), .S(_02296_), .Z(_02373__PTR100) );
  MUX2_X1 U8079 ( .A(P2_P1_InstAddrPointer_PTR5), .B(_02309__PTR5), .S(_02296_), .Z(_02373__PTR101) );
  MUX2_X1 U8080 ( .A(P2_P1_InstAddrPointer_PTR6), .B(_02309__PTR6), .S(_02296_), .Z(_02373__PTR102) );
  MUX2_X1 U8081 ( .A(P2_P1_InstAddrPointer_PTR7), .B(_02309__PTR7), .S(_02296_), .Z(_02373__PTR103) );
  MUX2_X1 U8082 ( .A(P2_P1_InstAddrPointer_PTR8), .B(_02309__PTR8), .S(_02296_), .Z(_02373__PTR104) );
  MUX2_X1 U8083 ( .A(P2_P1_InstAddrPointer_PTR9), .B(_02309__PTR9), .S(_02296_), .Z(_02373__PTR105) );
  MUX2_X1 U8084 ( .A(P2_P1_InstAddrPointer_PTR10), .B(_02309__PTR10), .S(_02296_), .Z(_02373__PTR106) );
  MUX2_X1 U8085 ( .A(P2_P1_InstAddrPointer_PTR11), .B(_02309__PTR11), .S(_02296_), .Z(_02373__PTR107) );
  MUX2_X1 U8086 ( .A(P2_P1_InstAddrPointer_PTR12), .B(_02309__PTR12), .S(_02296_), .Z(_02373__PTR108) );
  MUX2_X1 U8087 ( .A(P2_P1_InstAddrPointer_PTR13), .B(_02309__PTR13), .S(_02296_), .Z(_02373__PTR109) );
  MUX2_X1 U8088 ( .A(P2_P1_InstAddrPointer_PTR14), .B(_02309__PTR14), .S(_02296_), .Z(_02373__PTR110) );
  MUX2_X1 U8089 ( .A(P2_P1_InstAddrPointer_PTR15), .B(_02309__PTR15), .S(_02296_), .Z(_02373__PTR111) );
  MUX2_X1 U8090 ( .A(P2_P1_InstAddrPointer_PTR16), .B(_02309__PTR16), .S(_02296_), .Z(_02373__PTR112) );
  MUX2_X1 U8091 ( .A(P2_P1_InstAddrPointer_PTR17), .B(_02309__PTR17), .S(_02296_), .Z(_02373__PTR113) );
  MUX2_X1 U8092 ( .A(P2_P1_InstAddrPointer_PTR18), .B(_02309__PTR18), .S(_02296_), .Z(_02373__PTR114) );
  MUX2_X1 U8093 ( .A(P2_P1_InstAddrPointer_PTR19), .B(_02309__PTR19), .S(_02296_), .Z(_02373__PTR115) );
  MUX2_X1 U8094 ( .A(P2_P1_InstAddrPointer_PTR20), .B(_02309__PTR20), .S(_02296_), .Z(_02373__PTR116) );
  MUX2_X1 U8095 ( .A(P2_P1_InstAddrPointer_PTR21), .B(_02309__PTR21), .S(_02296_), .Z(_02373__PTR117) );
  MUX2_X1 U8096 ( .A(P2_P1_InstAddrPointer_PTR22), .B(_02309__PTR22), .S(_02296_), .Z(_02373__PTR118) );
  MUX2_X1 U8097 ( .A(P2_P1_InstAddrPointer_PTR23), .B(_02309__PTR23), .S(_02296_), .Z(_02373__PTR119) );
  MUX2_X1 U8098 ( .A(P2_P1_InstAddrPointer_PTR24), .B(_02309__PTR24), .S(_02296_), .Z(_02373__PTR120) );
  MUX2_X1 U8099 ( .A(P2_P1_InstAddrPointer_PTR25), .B(_02309__PTR25), .S(_02296_), .Z(_02373__PTR121) );
  MUX2_X1 U8100 ( .A(P2_P1_InstAddrPointer_PTR26), .B(_02309__PTR26), .S(_02296_), .Z(_02373__PTR122) );
  MUX2_X1 U8101 ( .A(P2_P1_InstAddrPointer_PTR27), .B(_02309__PTR27), .S(_02296_), .Z(_02373__PTR123) );
  MUX2_X1 U8102 ( .A(P2_P1_InstAddrPointer_PTR28), .B(_02309__PTR28), .S(_02296_), .Z(_02373__PTR124) );
  MUX2_X1 U8103 ( .A(P2_P1_InstAddrPointer_PTR29), .B(_02309__PTR29), .S(_02296_), .Z(_02373__PTR125) );
  MUX2_X1 U8104 ( .A(P2_P1_InstAddrPointer_PTR30), .B(_02309__PTR30), .S(_02296_), .Z(_02373__PTR126) );
  MUX2_X1 U8105 ( .A(P2_P1_InstAddrPointer_PTR31), .B(_02309__PTR31), .S(_02296_), .Z(_02373__PTR127) );
  MUX2_X1 U8106 ( .A(P2_P1_InstAddrPointer_PTR0), .B(_02290__PTR0), .S(_02146__PTR3), .Z(_02373__PTR192) );
  MUX2_X1 U8107 ( .A(P2_P1_InstAddrPointer_PTR1), .B(_02290__PTR1), .S(_02146__PTR3), .Z(_02373__PTR193) );
  MUX2_X1 U8108 ( .A(P2_P1_InstAddrPointer_PTR2), .B(_02290__PTR2), .S(_02146__PTR3), .Z(_02373__PTR194) );
  MUX2_X1 U8109 ( .A(P2_P1_InstAddrPointer_PTR3), .B(_02290__PTR3), .S(_02146__PTR3), .Z(_02373__PTR195) );
  MUX2_X1 U8110 ( .A(P2_P1_InstAddrPointer_PTR4), .B(_02290__PTR4), .S(_02146__PTR3), .Z(_02373__PTR196) );
  MUX2_X1 U8111 ( .A(P2_P1_InstAddrPointer_PTR5), .B(_02290__PTR5), .S(_02146__PTR3), .Z(_02373__PTR197) );
  MUX2_X1 U8112 ( .A(P2_P1_InstAddrPointer_PTR6), .B(_02290__PTR6), .S(_02146__PTR3), .Z(_02373__PTR198) );
  MUX2_X1 U8113 ( .A(P2_P1_InstAddrPointer_PTR7), .B(_02290__PTR7), .S(_02146__PTR3), .Z(_02373__PTR199) );
  MUX2_X1 U8114 ( .A(P2_P1_InstAddrPointer_PTR8), .B(_02290__PTR8), .S(_02146__PTR3), .Z(_02373__PTR200) );
  MUX2_X1 U8115 ( .A(P2_P1_InstAddrPointer_PTR9), .B(_02290__PTR9), .S(_02146__PTR3), .Z(_02373__PTR201) );
  MUX2_X1 U8116 ( .A(P2_P1_InstAddrPointer_PTR10), .B(_02290__PTR10), .S(_02146__PTR3), .Z(_02373__PTR202) );
  MUX2_X1 U8117 ( .A(P2_P1_InstAddrPointer_PTR11), .B(_02290__PTR11), .S(_02146__PTR3), .Z(_02373__PTR203) );
  MUX2_X1 U8118 ( .A(P2_P1_InstAddrPointer_PTR12), .B(_02290__PTR12), .S(_02146__PTR3), .Z(_02373__PTR204) );
  MUX2_X1 U8119 ( .A(P2_P1_InstAddrPointer_PTR13), .B(_02290__PTR13), .S(_02146__PTR3), .Z(_02373__PTR205) );
  MUX2_X1 U8120 ( .A(P2_P1_InstAddrPointer_PTR14), .B(_02290__PTR14), .S(_02146__PTR3), .Z(_02373__PTR206) );
  MUX2_X1 U8121 ( .A(P2_P1_InstAddrPointer_PTR15), .B(_02290__PTR15), .S(_02146__PTR3), .Z(_02373__PTR207) );
  MUX2_X1 U8122 ( .A(P2_P1_InstAddrPointer_PTR16), .B(_02290__PTR16), .S(_02146__PTR3), .Z(_02373__PTR208) );
  MUX2_X1 U8123 ( .A(P2_P1_InstAddrPointer_PTR17), .B(_02290__PTR17), .S(_02146__PTR3), .Z(_02373__PTR209) );
  MUX2_X1 U8124 ( .A(P2_P1_InstAddrPointer_PTR18), .B(_02290__PTR18), .S(_02146__PTR3), .Z(_02373__PTR210) );
  MUX2_X1 U8125 ( .A(P2_P1_InstAddrPointer_PTR19), .B(_02290__PTR19), .S(_02146__PTR3), .Z(_02373__PTR211) );
  MUX2_X1 U8126 ( .A(P2_P1_InstAddrPointer_PTR20), .B(_02290__PTR20), .S(_02146__PTR3), .Z(_02373__PTR212) );
  MUX2_X1 U8127 ( .A(P2_P1_InstAddrPointer_PTR21), .B(_02290__PTR21), .S(_02146__PTR3), .Z(_02373__PTR213) );
  MUX2_X1 U8128 ( .A(P2_P1_InstAddrPointer_PTR22), .B(_02290__PTR22), .S(_02146__PTR3), .Z(_02373__PTR214) );
  MUX2_X1 U8129 ( .A(P2_P1_InstAddrPointer_PTR23), .B(_02290__PTR23), .S(_02146__PTR3), .Z(_02373__PTR215) );
  MUX2_X1 U8130 ( .A(P2_P1_InstAddrPointer_PTR24), .B(_02290__PTR24), .S(_02146__PTR3), .Z(_02373__PTR216) );
  MUX2_X1 U8131 ( .A(P2_P1_InstAddrPointer_PTR25), .B(_02290__PTR25), .S(_02146__PTR3), .Z(_02373__PTR217) );
  MUX2_X1 U8132 ( .A(P2_P1_InstAddrPointer_PTR26), .B(_02290__PTR26), .S(_02146__PTR3), .Z(_02373__PTR218) );
  MUX2_X1 U8133 ( .A(P2_P1_InstAddrPointer_PTR27), .B(_02290__PTR27), .S(_02146__PTR3), .Z(_02373__PTR219) );
  MUX2_X1 U8134 ( .A(P2_P1_InstAddrPointer_PTR28), .B(_02290__PTR28), .S(_02146__PTR3), .Z(_02373__PTR220) );
  MUX2_X1 U8135 ( .A(P2_P1_InstAddrPointer_PTR29), .B(_02290__PTR29), .S(_02146__PTR3), .Z(_02373__PTR221) );
  MUX2_X1 U8136 ( .A(P2_P1_InstAddrPointer_PTR30), .B(_02290__PTR30), .S(_02146__PTR3), .Z(_02373__PTR222) );
  MUX2_X1 U8137 ( .A(P2_P1_InstAddrPointer_PTR31), .B(_02290__PTR31), .S(_02146__PTR3), .Z(_02373__PTR223) );
  MUX2_X1 U8138 ( .A(P2_P1_PhyAddrPointer_PTR0), .B(_02290__PTR0), .S(_02146__PTR3), .Z(_02381__PTR64) );
  MUX2_X1 U8139 ( .A(P2_P1_PhyAddrPointer_PTR1), .B(_02290__PTR1), .S(_02146__PTR3), .Z(_02381__PTR65) );
  MUX2_X1 U8140 ( .A(P2_P1_PhyAddrPointer_PTR2), .B(_02290__PTR2), .S(_02146__PTR3), .Z(_02381__PTR66) );
  MUX2_X1 U8141 ( .A(P2_P1_PhyAddrPointer_PTR3), .B(_02290__PTR3), .S(_02146__PTR3), .Z(_02381__PTR67) );
  MUX2_X1 U8142 ( .A(P2_P1_PhyAddrPointer_PTR4), .B(_02290__PTR4), .S(_02146__PTR3), .Z(_02381__PTR68) );
  MUX2_X1 U8143 ( .A(P2_P1_PhyAddrPointer_PTR5), .B(_02290__PTR5), .S(_02146__PTR3), .Z(_02381__PTR69) );
  MUX2_X1 U8144 ( .A(P2_P1_PhyAddrPointer_PTR6), .B(_02290__PTR6), .S(_02146__PTR3), .Z(_02381__PTR70) );
  MUX2_X1 U8145 ( .A(P2_P1_PhyAddrPointer_PTR7), .B(_02290__PTR7), .S(_02146__PTR3), .Z(_02381__PTR71) );
  MUX2_X1 U8146 ( .A(P2_P1_PhyAddrPointer_PTR8), .B(_02290__PTR8), .S(_02146__PTR3), .Z(_02381__PTR72) );
  MUX2_X1 U8147 ( .A(P2_P1_PhyAddrPointer_PTR9), .B(_02290__PTR9), .S(_02146__PTR3), .Z(_02381__PTR73) );
  MUX2_X1 U8148 ( .A(P2_P1_PhyAddrPointer_PTR10), .B(_02290__PTR10), .S(_02146__PTR3), .Z(_02381__PTR74) );
  MUX2_X1 U8149 ( .A(P2_P1_PhyAddrPointer_PTR11), .B(_02290__PTR11), .S(_02146__PTR3), .Z(_02381__PTR75) );
  MUX2_X1 U8150 ( .A(P2_P1_PhyAddrPointer_PTR12), .B(_02290__PTR12), .S(_02146__PTR3), .Z(_02381__PTR76) );
  MUX2_X1 U8151 ( .A(P2_P1_PhyAddrPointer_PTR13), .B(_02290__PTR13), .S(_02146__PTR3), .Z(_02381__PTR77) );
  MUX2_X1 U8152 ( .A(P2_P1_PhyAddrPointer_PTR14), .B(_02290__PTR14), .S(_02146__PTR3), .Z(_02381__PTR78) );
  MUX2_X1 U8153 ( .A(P2_P1_PhyAddrPointer_PTR15), .B(_02290__PTR15), .S(_02146__PTR3), .Z(_02381__PTR79) );
  MUX2_X1 U8154 ( .A(P2_P1_PhyAddrPointer_PTR16), .B(_02290__PTR16), .S(_02146__PTR3), .Z(_02381__PTR80) );
  MUX2_X1 U8155 ( .A(P2_P1_PhyAddrPointer_PTR17), .B(_02290__PTR17), .S(_02146__PTR3), .Z(_02381__PTR81) );
  MUX2_X1 U8156 ( .A(P2_P1_PhyAddrPointer_PTR18), .B(_02290__PTR18), .S(_02146__PTR3), .Z(_02381__PTR82) );
  MUX2_X1 U8157 ( .A(P2_P1_PhyAddrPointer_PTR19), .B(_02290__PTR19), .S(_02146__PTR3), .Z(_02381__PTR83) );
  MUX2_X1 U8158 ( .A(P2_P1_PhyAddrPointer_PTR20), .B(_02290__PTR20), .S(_02146__PTR3), .Z(_02381__PTR84) );
  MUX2_X1 U8159 ( .A(P2_P1_PhyAddrPointer_PTR21), .B(_02290__PTR21), .S(_02146__PTR3), .Z(_02381__PTR85) );
  MUX2_X1 U8160 ( .A(P2_P1_PhyAddrPointer_PTR22), .B(_02290__PTR22), .S(_02146__PTR3), .Z(_02381__PTR86) );
  MUX2_X1 U8161 ( .A(P2_P1_PhyAddrPointer_PTR23), .B(_02290__PTR23), .S(_02146__PTR3), .Z(_02381__PTR87) );
  MUX2_X1 U8162 ( .A(P2_P1_PhyAddrPointer_PTR24), .B(_02290__PTR24), .S(_02146__PTR3), .Z(_02381__PTR88) );
  MUX2_X1 U8163 ( .A(P2_P1_PhyAddrPointer_PTR25), .B(_02290__PTR25), .S(_02146__PTR3), .Z(_02381__PTR89) );
  MUX2_X1 U8164 ( .A(P2_P1_PhyAddrPointer_PTR26), .B(_02290__PTR26), .S(_02146__PTR3), .Z(_02381__PTR90) );
  MUX2_X1 U8165 ( .A(P2_P1_PhyAddrPointer_PTR27), .B(_02290__PTR27), .S(_02146__PTR3), .Z(_02381__PTR91) );
  MUX2_X1 U8166 ( .A(P2_P1_PhyAddrPointer_PTR28), .B(_02290__PTR28), .S(_02146__PTR3), .Z(_02381__PTR92) );
  MUX2_X1 U8167 ( .A(P2_P1_PhyAddrPointer_PTR29), .B(_02290__PTR29), .S(_02146__PTR3), .Z(_02381__PTR93) );
  MUX2_X1 U8168 ( .A(P2_P1_PhyAddrPointer_PTR30), .B(_02290__PTR30), .S(_02146__PTR3), .Z(_02381__PTR94) );
  MUX2_X1 U8169 ( .A(P2_P1_PhyAddrPointer_PTR31), .B(_02290__PTR31), .S(_02146__PTR3), .Z(_02381__PTR95) );
  MUX2_X1 U8170 ( .A(_03184__PTR0), .B(_03048__PTR0), .S(_02969__PTR7), .Z(_02290__PTR0) );
  MUX2_X1 U8171 ( .A(_03184__PTR1), .B(_03049__PTR1), .S(_02969__PTR7), .Z(_02290__PTR1) );
  MUX2_X1 U8172 ( .A(_03184__PTR2), .B(_03049__PTR2), .S(_02969__PTR7), .Z(_02290__PTR2) );
  MUX2_X1 U8173 ( .A(_03184__PTR3), .B(_03049__PTR3), .S(_02969__PTR7), .Z(_02290__PTR3) );
  MUX2_X1 U8174 ( .A(_03184__PTR4), .B(_03049__PTR4), .S(_02969__PTR7), .Z(_02290__PTR4) );
  MUX2_X1 U8175 ( .A(_03184__PTR5), .B(_03049__PTR5), .S(_02969__PTR7), .Z(_02290__PTR5) );
  MUX2_X1 U8176 ( .A(_03184__PTR6), .B(_03049__PTR6), .S(_02969__PTR7), .Z(_02290__PTR6) );
  MUX2_X1 U8177 ( .A(_03184__PTR7), .B(_03049__PTR7), .S(_02969__PTR7), .Z(_02290__PTR7) );
  MUX2_X1 U8178 ( .A(_03184__PTR8), .B(_03049__PTR8), .S(_02969__PTR7), .Z(_02290__PTR8) );
  MUX2_X1 U8179 ( .A(_03184__PTR9), .B(_03049__PTR9), .S(_02969__PTR7), .Z(_02290__PTR9) );
  MUX2_X1 U8180 ( .A(_03184__PTR10), .B(_03049__PTR10), .S(_02969__PTR7), .Z(_02290__PTR10) );
  MUX2_X1 U8181 ( .A(_03184__PTR11), .B(_03049__PTR11), .S(_02969__PTR7), .Z(_02290__PTR11) );
  MUX2_X1 U8182 ( .A(_03184__PTR12), .B(_03049__PTR12), .S(_02969__PTR7), .Z(_02290__PTR12) );
  MUX2_X1 U8183 ( .A(_03184__PTR13), .B(_03049__PTR13), .S(_02969__PTR7), .Z(_02290__PTR13) );
  MUX2_X1 U8184 ( .A(_03184__PTR14), .B(_03049__PTR14), .S(_02969__PTR7), .Z(_02290__PTR14) );
  MUX2_X1 U8185 ( .A(_03184__PTR15), .B(_03049__PTR15), .S(_02969__PTR7), .Z(_02290__PTR15) );
  MUX2_X1 U8186 ( .A(_03184__PTR16), .B(_03049__PTR16), .S(_02969__PTR7), .Z(_02290__PTR16) );
  MUX2_X1 U8187 ( .A(_03184__PTR17), .B(_03049__PTR17), .S(_02969__PTR7), .Z(_02290__PTR17) );
  MUX2_X1 U8188 ( .A(_03184__PTR18), .B(_03049__PTR18), .S(_02969__PTR7), .Z(_02290__PTR18) );
  MUX2_X1 U8189 ( .A(_03184__PTR19), .B(_03049__PTR19), .S(_02969__PTR7), .Z(_02290__PTR19) );
  MUX2_X1 U8190 ( .A(_03184__PTR20), .B(_03049__PTR20), .S(_02969__PTR7), .Z(_02290__PTR20) );
  MUX2_X1 U8191 ( .A(_03184__PTR21), .B(_03049__PTR21), .S(_02969__PTR7), .Z(_02290__PTR21) );
  MUX2_X1 U8192 ( .A(_03184__PTR22), .B(_03049__PTR22), .S(_02969__PTR7), .Z(_02290__PTR22) );
  MUX2_X1 U8193 ( .A(_03184__PTR23), .B(_03049__PTR23), .S(_02969__PTR7), .Z(_02290__PTR23) );
  MUX2_X1 U8194 ( .A(_03184__PTR24), .B(_03049__PTR24), .S(_02969__PTR7), .Z(_02290__PTR24) );
  MUX2_X1 U8195 ( .A(_03184__PTR25), .B(_03049__PTR25), .S(_02969__PTR7), .Z(_02290__PTR25) );
  MUX2_X1 U8196 ( .A(_03184__PTR26), .B(_03049__PTR26), .S(_02969__PTR7), .Z(_02290__PTR26) );
  MUX2_X1 U8197 ( .A(_03184__PTR27), .B(_03049__PTR27), .S(_02969__PTR7), .Z(_02290__PTR27) );
  MUX2_X1 U8198 ( .A(_03184__PTR28), .B(_03049__PTR28), .S(_02969__PTR7), .Z(_02290__PTR28) );
  MUX2_X1 U8199 ( .A(_03184__PTR29), .B(_03049__PTR29), .S(_02969__PTR7), .Z(_02290__PTR29) );
  MUX2_X1 U8200 ( .A(_03184__PTR30), .B(_03049__PTR30), .S(_02969__PTR7), .Z(_02290__PTR30) );
  MUX2_X1 U8201 ( .A(_03184__PTR31), .B(_03049__PTR31), .S(_02969__PTR7), .Z(_02290__PTR31) );
  MUX2_X1 U8202 ( .A(P2_P1_PhyAddrPointer_PTR0), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR128) );
  MUX2_X1 U8203 ( .A(_02288__PTR1), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR129) );
  MUX2_X1 U8204 ( .A(_02288__PTR2), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR130) );
  MUX2_X1 U8205 ( .A(_02288__PTR3), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR131) );
  MUX2_X1 U8206 ( .A(_02288__PTR4), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR132) );
  MUX2_X1 U8207 ( .A(_02288__PTR5), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR133) );
  MUX2_X1 U8208 ( .A(_02288__PTR6), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR134) );
  MUX2_X1 U8209 ( .A(_02288__PTR7), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR135) );
  MUX2_X1 U8210 ( .A(_02288__PTR8), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR136) );
  MUX2_X1 U8211 ( .A(_02288__PTR9), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR137) );
  MUX2_X1 U8212 ( .A(_02288__PTR10), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR138) );
  MUX2_X1 U8213 ( .A(_02288__PTR11), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR139) );
  MUX2_X1 U8214 ( .A(_02288__PTR12), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR140) );
  MUX2_X1 U8215 ( .A(_02288__PTR13), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR141) );
  MUX2_X1 U8216 ( .A(_02288__PTR14), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR142) );
  MUX2_X1 U8217 ( .A(_02288__PTR15), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR143) );
  MUX2_X1 U8218 ( .A(_02288__PTR16), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR144) );
  MUX2_X1 U8219 ( .A(_02288__PTR17), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR145) );
  MUX2_X1 U8220 ( .A(_02288__PTR18), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR146) );
  MUX2_X1 U8221 ( .A(_02288__PTR19), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR147) );
  MUX2_X1 U8222 ( .A(_02288__PTR20), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR148) );
  MUX2_X1 U8223 ( .A(_02288__PTR21), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR149) );
  MUX2_X1 U8224 ( .A(_02288__PTR22), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR150) );
  MUX2_X1 U8225 ( .A(_02288__PTR23), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR151) );
  MUX2_X1 U8226 ( .A(_02288__PTR24), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR152) );
  MUX2_X1 U8227 ( .A(_02288__PTR25), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR153) );
  MUX2_X1 U8228 ( .A(_02288__PTR26), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR154) );
  MUX2_X1 U8229 ( .A(_02288__PTR27), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR155) );
  MUX2_X1 U8230 ( .A(_02288__PTR28), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR156) );
  MUX2_X1 U8231 ( .A(_02288__PTR29), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR157) );
  MUX2_X1 U8232 ( .A(_02288__PTR30), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR158) );
  MUX2_X1 U8233 ( .A(_02288__PTR31), .B(1'b0), .S(P2_StateBS16), .Z(_02188__PTR160) );
  MUX2_X1 U8234 ( .A(_02184__PTR129), .B(1'b0), .S(P2_StateBS16), .Z(_02184__PTR65) );
  MUX2_X1 U8235 ( .A(_02184__PTR130), .B(_03040__PTR0), .S(P2_StateBS16), .Z(_02184__PTR66) );
  MUX2_X1 U8236 ( .A(_02184__PTR131), .B(_03041__PTR1), .S(P2_StateBS16), .Z(_02184__PTR67) );
  MUX2_X1 U8237 ( .A(_02184__PTR132), .B(_03041__PTR2), .S(P2_StateBS16), .Z(_02184__PTR68) );
  MUX2_X1 U8238 ( .A(_02184__PTR133), .B(_03041__PTR3), .S(P2_StateBS16), .Z(_02184__PTR69) );
  MUX2_X1 U8239 ( .A(_02184__PTR134), .B(_03041__PTR4), .S(P2_StateBS16), .Z(_02184__PTR70) );
  MUX2_X1 U8240 ( .A(_02184__PTR135), .B(_03041__PTR5), .S(P2_StateBS16), .Z(_02184__PTR71) );
  MUX2_X1 U8241 ( .A(_02184__PTR136), .B(_03041__PTR6), .S(P2_StateBS16), .Z(_02184__PTR72) );
  MUX2_X1 U8242 ( .A(_02184__PTR137), .B(_03041__PTR7), .S(P2_StateBS16), .Z(_02184__PTR73) );
  MUX2_X1 U8243 ( .A(_02184__PTR138), .B(_03041__PTR8), .S(P2_StateBS16), .Z(_02184__PTR74) );
  MUX2_X1 U8244 ( .A(_02184__PTR139), .B(_03041__PTR9), .S(P2_StateBS16), .Z(_02184__PTR75) );
  MUX2_X1 U8245 ( .A(_02184__PTR140), .B(_03041__PTR10), .S(P2_StateBS16), .Z(_02184__PTR76) );
  MUX2_X1 U8246 ( .A(_02184__PTR141), .B(_03041__PTR11), .S(P2_StateBS16), .Z(_02184__PTR77) );
  MUX2_X1 U8247 ( .A(_02184__PTR142), .B(_03041__PTR12), .S(P2_StateBS16), .Z(_02184__PTR78) );
  MUX2_X1 U8248 ( .A(_02184__PTR143), .B(_03041__PTR13), .S(P2_StateBS16), .Z(_02184__PTR79) );
  MUX2_X1 U8249 ( .A(_02184__PTR144), .B(_03041__PTR14), .S(P2_StateBS16), .Z(_02184__PTR80) );
  MUX2_X1 U8250 ( .A(_02184__PTR145), .B(_03041__PTR15), .S(P2_StateBS16), .Z(_02184__PTR81) );
  MUX2_X1 U8251 ( .A(_02184__PTR146), .B(_03041__PTR16), .S(P2_StateBS16), .Z(_02184__PTR82) );
  MUX2_X1 U8252 ( .A(_02184__PTR147), .B(_03041__PTR17), .S(P2_StateBS16), .Z(_02184__PTR83) );
  MUX2_X1 U8253 ( .A(_02184__PTR148), .B(_03041__PTR18), .S(P2_StateBS16), .Z(_02184__PTR84) );
  MUX2_X1 U8254 ( .A(_02184__PTR149), .B(_03041__PTR19), .S(P2_StateBS16), .Z(_02184__PTR85) );
  MUX2_X1 U8255 ( .A(_02184__PTR150), .B(_03041__PTR20), .S(P2_StateBS16), .Z(_02184__PTR86) );
  MUX2_X1 U8256 ( .A(_02184__PTR151), .B(_03041__PTR21), .S(P2_StateBS16), .Z(_02184__PTR87) );
  MUX2_X1 U8257 ( .A(_02184__PTR152), .B(_03041__PTR22), .S(P2_StateBS16), .Z(_02184__PTR88) );
  MUX2_X1 U8258 ( .A(_02184__PTR153), .B(_03041__PTR23), .S(P2_StateBS16), .Z(_02184__PTR89) );
  MUX2_X1 U8259 ( .A(_02184__PTR154), .B(_03041__PTR24), .S(P2_StateBS16), .Z(_02184__PTR90) );
  MUX2_X1 U8260 ( .A(_02184__PTR155), .B(_03041__PTR25), .S(P2_StateBS16), .Z(_02184__PTR91) );
  MUX2_X1 U8261 ( .A(_02184__PTR156), .B(_03041__PTR26), .S(P2_StateBS16), .Z(_02184__PTR92) );
  MUX2_X1 U8262 ( .A(_02184__PTR157), .B(_03041__PTR27), .S(P2_StateBS16), .Z(_02184__PTR93) );
  MUX2_X1 U8263 ( .A(_02184__PTR158), .B(_03041__PTR28), .S(P2_StateBS16), .Z(_02184__PTR94) );
  MUX2_X1 U8264 ( .A(_02184__PTR159), .B(_03041__PTR29), .S(P2_StateBS16), .Z(_02184__PTR95) );
  MUX2_X1 U8265 ( .A(_02131__PTR1), .B(_03036__PTR1), .S(P2_StateBS16), .Z(_02222__PTR17) );
  MUX2_X1 U8266 ( .A(_02131__PTR2), .B(_03036__PTR2), .S(P2_StateBS16), .Z(_02222__PTR18) );
  MUX2_X1 U8267 ( .A(_02131__PTR3), .B(_03036__PTR3), .S(P2_StateBS16), .Z(_02222__PTR19) );
  MUX2_X1 U8268 ( .A(_02220__PTR32), .B(_02287__PTR0), .S(P2_StateBS16), .Z(_02220__PTR16) );
  MUX2_X1 U8269 ( .A(_02220__PTR33), .B(_02287__PTR1), .S(P2_StateBS16), .Z(_02220__PTR17) );
  MUX2_X1 U8270 ( .A(_02220__PTR34), .B(_02287__PTR2), .S(P2_StateBS16), .Z(_02220__PTR18) );
  MUX2_X1 U8271 ( .A(_02220__PTR35), .B(_02287__PTR3), .S(P2_StateBS16), .Z(_02220__PTR19) );
  MUX2_X1 U8272 ( .A(_02220__PTR36), .B(_02287__PTR4), .S(P2_StateBS16), .Z(_02220__PTR20) );
  MUX2_X1 U8273 ( .A(_02220__PTR37), .B(_02287__PTR5), .S(P2_StateBS16), .Z(_02220__PTR21) );
  MUX2_X1 U8274 ( .A(_02220__PTR38), .B(_02287__PTR6), .S(P2_StateBS16), .Z(_02220__PTR22) );
  MUX2_X1 U8275 ( .A(_02220__PTR39), .B(_02287__PTR7), .S(P2_StateBS16), .Z(_02220__PTR23) );
  MUX2_X1 U8276 ( .A(_02218__PTR32), .B(_02286__PTR0), .S(P2_StateBS16), .Z(_02218__PTR16) );
  MUX2_X1 U8277 ( .A(_02218__PTR33), .B(_02286__PTR1), .S(P2_StateBS16), .Z(_02218__PTR17) );
  MUX2_X1 U8278 ( .A(_02218__PTR34), .B(_02286__PTR2), .S(P2_StateBS16), .Z(_02218__PTR18) );
  MUX2_X1 U8279 ( .A(_02218__PTR35), .B(_02286__PTR3), .S(P2_StateBS16), .Z(_02218__PTR19) );
  MUX2_X1 U8280 ( .A(_02218__PTR36), .B(_02286__PTR4), .S(P2_StateBS16), .Z(_02218__PTR20) );
  MUX2_X1 U8281 ( .A(_02218__PTR37), .B(_02286__PTR5), .S(P2_StateBS16), .Z(_02218__PTR21) );
  MUX2_X1 U8282 ( .A(_02218__PTR38), .B(_02286__PTR6), .S(P2_StateBS16), .Z(_02218__PTR22) );
  MUX2_X1 U8283 ( .A(_02218__PTR39), .B(_02286__PTR7), .S(P2_StateBS16), .Z(_02218__PTR23) );
  MUX2_X1 U8284 ( .A(_02216__PTR32), .B(_02285__PTR0), .S(P2_StateBS16), .Z(_02216__PTR16) );
  MUX2_X1 U8285 ( .A(_02216__PTR33), .B(_02285__PTR1), .S(P2_StateBS16), .Z(_02216__PTR17) );
  MUX2_X1 U8286 ( .A(_02216__PTR34), .B(_02285__PTR2), .S(P2_StateBS16), .Z(_02216__PTR18) );
  MUX2_X1 U8287 ( .A(_02216__PTR35), .B(_02285__PTR3), .S(P2_StateBS16), .Z(_02216__PTR19) );
  MUX2_X1 U8288 ( .A(_02216__PTR36), .B(_02285__PTR4), .S(P2_StateBS16), .Z(_02216__PTR20) );
  MUX2_X1 U8289 ( .A(_02216__PTR37), .B(_02285__PTR5), .S(P2_StateBS16), .Z(_02216__PTR21) );
  MUX2_X1 U8290 ( .A(_02216__PTR38), .B(_02285__PTR6), .S(P2_StateBS16), .Z(_02216__PTR22) );
  MUX2_X1 U8291 ( .A(_02216__PTR39), .B(_02285__PTR7), .S(P2_StateBS16), .Z(_02216__PTR23) );
  MUX2_X1 U8292 ( .A(_02214__PTR32), .B(_02284__PTR0), .S(P2_StateBS16), .Z(_02214__PTR16) );
  MUX2_X1 U8293 ( .A(_02214__PTR33), .B(_02284__PTR1), .S(P2_StateBS16), .Z(_02214__PTR17) );
  MUX2_X1 U8294 ( .A(_02214__PTR34), .B(_02284__PTR2), .S(P2_StateBS16), .Z(_02214__PTR18) );
  MUX2_X1 U8295 ( .A(_02214__PTR35), .B(_02284__PTR3), .S(P2_StateBS16), .Z(_02214__PTR19) );
  MUX2_X1 U8296 ( .A(_02214__PTR36), .B(_02284__PTR4), .S(P2_StateBS16), .Z(_02214__PTR20) );
  MUX2_X1 U8297 ( .A(_02214__PTR37), .B(_02284__PTR5), .S(P2_StateBS16), .Z(_02214__PTR21) );
  MUX2_X1 U8298 ( .A(_02214__PTR38), .B(_02284__PTR6), .S(P2_StateBS16), .Z(_02214__PTR22) );
  MUX2_X1 U8299 ( .A(_02214__PTR39), .B(_02284__PTR7), .S(P2_StateBS16), .Z(_02214__PTR23) );
  MUX2_X1 U8300 ( .A(_02212__PTR32), .B(_02283__PTR0), .S(P2_StateBS16), .Z(_02212__PTR16) );
  MUX2_X1 U8301 ( .A(_02212__PTR33), .B(_02283__PTR1), .S(P2_StateBS16), .Z(_02212__PTR17) );
  MUX2_X1 U8302 ( .A(_02212__PTR34), .B(_02283__PTR2), .S(P2_StateBS16), .Z(_02212__PTR18) );
  MUX2_X1 U8303 ( .A(_02212__PTR35), .B(_02283__PTR3), .S(P2_StateBS16), .Z(_02212__PTR19) );
  MUX2_X1 U8304 ( .A(_02212__PTR36), .B(_02283__PTR4), .S(P2_StateBS16), .Z(_02212__PTR20) );
  MUX2_X1 U8305 ( .A(_02212__PTR37), .B(_02283__PTR5), .S(P2_StateBS16), .Z(_02212__PTR21) );
  MUX2_X1 U8306 ( .A(_02212__PTR38), .B(_02283__PTR6), .S(P2_StateBS16), .Z(_02212__PTR22) );
  MUX2_X1 U8307 ( .A(_02212__PTR39), .B(_02283__PTR7), .S(P2_StateBS16), .Z(_02212__PTR23) );
  MUX2_X1 U8308 ( .A(_02210__PTR32), .B(_02282__PTR0), .S(P2_StateBS16), .Z(_02210__PTR16) );
  MUX2_X1 U8309 ( .A(_02210__PTR33), .B(_02282__PTR1), .S(P2_StateBS16), .Z(_02210__PTR17) );
  MUX2_X1 U8310 ( .A(_02210__PTR34), .B(_02282__PTR2), .S(P2_StateBS16), .Z(_02210__PTR18) );
  MUX2_X1 U8311 ( .A(_02210__PTR35), .B(_02282__PTR3), .S(P2_StateBS16), .Z(_02210__PTR19) );
  MUX2_X1 U8312 ( .A(_02210__PTR36), .B(_02282__PTR4), .S(P2_StateBS16), .Z(_02210__PTR20) );
  MUX2_X1 U8313 ( .A(_02210__PTR37), .B(_02282__PTR5), .S(P2_StateBS16), .Z(_02210__PTR21) );
  MUX2_X1 U8314 ( .A(_02210__PTR38), .B(_02282__PTR6), .S(P2_StateBS16), .Z(_02210__PTR22) );
  MUX2_X1 U8315 ( .A(_02210__PTR39), .B(_02282__PTR7), .S(P2_StateBS16), .Z(_02210__PTR23) );
  MUX2_X1 U8316 ( .A(_02208__PTR32), .B(_02281__PTR0), .S(P2_StateBS16), .Z(_02208__PTR16) );
  MUX2_X1 U8317 ( .A(_02208__PTR33), .B(_02281__PTR1), .S(P2_StateBS16), .Z(_02208__PTR17) );
  MUX2_X1 U8318 ( .A(_02208__PTR34), .B(_02281__PTR2), .S(P2_StateBS16), .Z(_02208__PTR18) );
  MUX2_X1 U8319 ( .A(_02208__PTR35), .B(_02281__PTR3), .S(P2_StateBS16), .Z(_02208__PTR19) );
  MUX2_X1 U8320 ( .A(_02208__PTR36), .B(_02281__PTR4), .S(P2_StateBS16), .Z(_02208__PTR20) );
  MUX2_X1 U8321 ( .A(_02208__PTR37), .B(_02281__PTR5), .S(P2_StateBS16), .Z(_02208__PTR21) );
  MUX2_X1 U8322 ( .A(_02208__PTR38), .B(_02281__PTR6), .S(P2_StateBS16), .Z(_02208__PTR22) );
  MUX2_X1 U8323 ( .A(_02208__PTR39), .B(_02281__PTR7), .S(P2_StateBS16), .Z(_02208__PTR23) );
  MUX2_X1 U8324 ( .A(_02206__PTR32), .B(_02280__PTR0), .S(P2_StateBS16), .Z(_02206__PTR16) );
  MUX2_X1 U8325 ( .A(_02206__PTR33), .B(_02280__PTR1), .S(P2_StateBS16), .Z(_02206__PTR17) );
  MUX2_X1 U8326 ( .A(_02206__PTR34), .B(_02280__PTR2), .S(P2_StateBS16), .Z(_02206__PTR18) );
  MUX2_X1 U8327 ( .A(_02206__PTR35), .B(_02280__PTR3), .S(P2_StateBS16), .Z(_02206__PTR19) );
  MUX2_X1 U8328 ( .A(_02206__PTR36), .B(_02280__PTR4), .S(P2_StateBS16), .Z(_02206__PTR20) );
  MUX2_X1 U8329 ( .A(_02206__PTR37), .B(_02280__PTR5), .S(P2_StateBS16), .Z(_02206__PTR21) );
  MUX2_X1 U8330 ( .A(_02206__PTR38), .B(_02280__PTR6), .S(P2_StateBS16), .Z(_02206__PTR22) );
  MUX2_X1 U8331 ( .A(_02206__PTR39), .B(_02280__PTR7), .S(P2_StateBS16), .Z(_02206__PTR23) );
  MUX2_X1 U8332 ( .A(_02204__PTR32), .B(_02279__PTR0), .S(P2_StateBS16), .Z(_02204__PTR16) );
  MUX2_X1 U8333 ( .A(_02204__PTR33), .B(_02279__PTR1), .S(P2_StateBS16), .Z(_02204__PTR17) );
  MUX2_X1 U8334 ( .A(_02204__PTR34), .B(_02279__PTR2), .S(P2_StateBS16), .Z(_02204__PTR18) );
  MUX2_X1 U8335 ( .A(_02204__PTR35), .B(_02279__PTR3), .S(P2_StateBS16), .Z(_02204__PTR19) );
  MUX2_X1 U8336 ( .A(_02204__PTR36), .B(_02279__PTR4), .S(P2_StateBS16), .Z(_02204__PTR20) );
  MUX2_X1 U8337 ( .A(_02204__PTR37), .B(_02279__PTR5), .S(P2_StateBS16), .Z(_02204__PTR21) );
  MUX2_X1 U8338 ( .A(_02204__PTR38), .B(_02279__PTR6), .S(P2_StateBS16), .Z(_02204__PTR22) );
  MUX2_X1 U8339 ( .A(_02204__PTR39), .B(_02279__PTR7), .S(P2_StateBS16), .Z(_02204__PTR23) );
  MUX2_X1 U8340 ( .A(_02202__PTR32), .B(_02278__PTR0), .S(P2_StateBS16), .Z(_02202__PTR16) );
  MUX2_X1 U8341 ( .A(_02202__PTR33), .B(_02278__PTR1), .S(P2_StateBS16), .Z(_02202__PTR17) );
  MUX2_X1 U8342 ( .A(_02202__PTR34), .B(_02278__PTR2), .S(P2_StateBS16), .Z(_02202__PTR18) );
  MUX2_X1 U8343 ( .A(_02202__PTR35), .B(_02278__PTR3), .S(P2_StateBS16), .Z(_02202__PTR19) );
  MUX2_X1 U8344 ( .A(_02202__PTR36), .B(_02278__PTR4), .S(P2_StateBS16), .Z(_02202__PTR20) );
  MUX2_X1 U8345 ( .A(_02202__PTR37), .B(_02278__PTR5), .S(P2_StateBS16), .Z(_02202__PTR21) );
  MUX2_X1 U8346 ( .A(_02202__PTR38), .B(_02278__PTR6), .S(P2_StateBS16), .Z(_02202__PTR22) );
  MUX2_X1 U8347 ( .A(_02202__PTR39), .B(_02278__PTR7), .S(P2_StateBS16), .Z(_02202__PTR23) );
  MUX2_X1 U8348 ( .A(_02200__PTR32), .B(_02277__PTR0), .S(P2_StateBS16), .Z(_02200__PTR16) );
  MUX2_X1 U8349 ( .A(_02200__PTR33), .B(_02277__PTR1), .S(P2_StateBS16), .Z(_02200__PTR17) );
  MUX2_X1 U8350 ( .A(_02200__PTR34), .B(_02277__PTR2), .S(P2_StateBS16), .Z(_02200__PTR18) );
  MUX2_X1 U8351 ( .A(_02200__PTR35), .B(_02277__PTR3), .S(P2_StateBS16), .Z(_02200__PTR19) );
  MUX2_X1 U8352 ( .A(_02200__PTR36), .B(_02277__PTR4), .S(P2_StateBS16), .Z(_02200__PTR20) );
  MUX2_X1 U8353 ( .A(_02200__PTR37), .B(_02277__PTR5), .S(P2_StateBS16), .Z(_02200__PTR21) );
  MUX2_X1 U8354 ( .A(_02200__PTR38), .B(_02277__PTR6), .S(P2_StateBS16), .Z(_02200__PTR22) );
  MUX2_X1 U8355 ( .A(_02200__PTR39), .B(_02277__PTR7), .S(P2_StateBS16), .Z(_02200__PTR23) );
  MUX2_X1 U8356 ( .A(_02198__PTR32), .B(_02276__PTR0), .S(P2_StateBS16), .Z(_02198__PTR16) );
  MUX2_X1 U8357 ( .A(_02198__PTR33), .B(_02276__PTR1), .S(P2_StateBS16), .Z(_02198__PTR17) );
  MUX2_X1 U8358 ( .A(_02198__PTR34), .B(_02276__PTR2), .S(P2_StateBS16), .Z(_02198__PTR18) );
  MUX2_X1 U8359 ( .A(_02198__PTR35), .B(_02276__PTR3), .S(P2_StateBS16), .Z(_02198__PTR19) );
  MUX2_X1 U8360 ( .A(_02198__PTR36), .B(_02276__PTR4), .S(P2_StateBS16), .Z(_02198__PTR20) );
  MUX2_X1 U8361 ( .A(_02198__PTR37), .B(_02276__PTR5), .S(P2_StateBS16), .Z(_02198__PTR21) );
  MUX2_X1 U8362 ( .A(_02198__PTR38), .B(_02276__PTR6), .S(P2_StateBS16), .Z(_02198__PTR22) );
  MUX2_X1 U8363 ( .A(_02198__PTR39), .B(_02276__PTR7), .S(P2_StateBS16), .Z(_02198__PTR23) );
  MUX2_X1 U8364 ( .A(_02196__PTR32), .B(_02275__PTR0), .S(P2_StateBS16), .Z(_02196__PTR16) );
  MUX2_X1 U8365 ( .A(_02196__PTR33), .B(_02275__PTR1), .S(P2_StateBS16), .Z(_02196__PTR17) );
  MUX2_X1 U8366 ( .A(_02196__PTR34), .B(_02275__PTR2), .S(P2_StateBS16), .Z(_02196__PTR18) );
  MUX2_X1 U8367 ( .A(_02196__PTR35), .B(_02275__PTR3), .S(P2_StateBS16), .Z(_02196__PTR19) );
  MUX2_X1 U8368 ( .A(_02196__PTR36), .B(_02275__PTR4), .S(P2_StateBS16), .Z(_02196__PTR20) );
  MUX2_X1 U8369 ( .A(_02196__PTR37), .B(_02275__PTR5), .S(P2_StateBS16), .Z(_02196__PTR21) );
  MUX2_X1 U8370 ( .A(_02196__PTR38), .B(_02275__PTR6), .S(P2_StateBS16), .Z(_02196__PTR22) );
  MUX2_X1 U8371 ( .A(_02196__PTR39), .B(_02275__PTR7), .S(P2_StateBS16), .Z(_02196__PTR23) );
  MUX2_X1 U8372 ( .A(_02194__PTR32), .B(_02274__PTR0), .S(P2_StateBS16), .Z(_02194__PTR16) );
  MUX2_X1 U8373 ( .A(_02194__PTR33), .B(_02274__PTR1), .S(P2_StateBS16), .Z(_02194__PTR17) );
  MUX2_X1 U8374 ( .A(_02194__PTR34), .B(_02274__PTR2), .S(P2_StateBS16), .Z(_02194__PTR18) );
  MUX2_X1 U8375 ( .A(_02194__PTR35), .B(_02274__PTR3), .S(P2_StateBS16), .Z(_02194__PTR19) );
  MUX2_X1 U8376 ( .A(_02194__PTR36), .B(_02274__PTR4), .S(P2_StateBS16), .Z(_02194__PTR20) );
  MUX2_X1 U8377 ( .A(_02194__PTR37), .B(_02274__PTR5), .S(P2_StateBS16), .Z(_02194__PTR21) );
  MUX2_X1 U8378 ( .A(_02194__PTR38), .B(_02274__PTR6), .S(P2_StateBS16), .Z(_02194__PTR22) );
  MUX2_X1 U8379 ( .A(_02194__PTR39), .B(_02274__PTR7), .S(P2_StateBS16), .Z(_02194__PTR23) );
  MUX2_X1 U8380 ( .A(_02192__PTR32), .B(_02273__PTR0), .S(P2_StateBS16), .Z(_02192__PTR16) );
  MUX2_X1 U8381 ( .A(_02192__PTR33), .B(_02273__PTR1), .S(P2_StateBS16), .Z(_02192__PTR17) );
  MUX2_X1 U8382 ( .A(_02192__PTR34), .B(_02273__PTR2), .S(P2_StateBS16), .Z(_02192__PTR18) );
  MUX2_X1 U8383 ( .A(_02192__PTR35), .B(_02273__PTR3), .S(P2_StateBS16), .Z(_02192__PTR19) );
  MUX2_X1 U8384 ( .A(_02192__PTR36), .B(_02273__PTR4), .S(P2_StateBS16), .Z(_02192__PTR20) );
  MUX2_X1 U8385 ( .A(_02192__PTR37), .B(_02273__PTR5), .S(P2_StateBS16), .Z(_02192__PTR21) );
  MUX2_X1 U8386 ( .A(_02192__PTR38), .B(_02273__PTR6), .S(P2_StateBS16), .Z(_02192__PTR22) );
  MUX2_X1 U8387 ( .A(_02192__PTR39), .B(_02273__PTR7), .S(P2_StateBS16), .Z(_02192__PTR23) );
  MUX2_X1 U8388 ( .A(_02190__PTR32), .B(_02272__PTR0), .S(P2_StateBS16), .Z(_02190__PTR16) );
  MUX2_X1 U8389 ( .A(_02190__PTR33), .B(_02272__PTR1), .S(P2_StateBS16), .Z(_02190__PTR17) );
  MUX2_X1 U8390 ( .A(_02190__PTR34), .B(_02272__PTR2), .S(P2_StateBS16), .Z(_02190__PTR18) );
  MUX2_X1 U8391 ( .A(_02190__PTR35), .B(_02272__PTR3), .S(P2_StateBS16), .Z(_02190__PTR19) );
  MUX2_X1 U8392 ( .A(_02190__PTR36), .B(_02272__PTR4), .S(P2_StateBS16), .Z(_02190__PTR20) );
  MUX2_X1 U8393 ( .A(_02190__PTR37), .B(_02272__PTR5), .S(P2_StateBS16), .Z(_02190__PTR21) );
  MUX2_X1 U8394 ( .A(_02190__PTR38), .B(_02272__PTR6), .S(P2_StateBS16), .Z(_02190__PTR22) );
  MUX2_X1 U8395 ( .A(_02190__PTR39), .B(_02272__PTR7), .S(P2_StateBS16), .Z(_02190__PTR23) );
  MUX2_X1 U8396 ( .A(_03191__PTR1), .B(_02184__PTR129), .S(_02959__PTR31), .Z(_02288__PTR1) );
  MUX2_X1 U8397 ( .A(_03191__PTR2), .B(_02184__PTR130), .S(_02959__PTR31), .Z(_02288__PTR2) );
  MUX2_X1 U8398 ( .A(_03191__PTR3), .B(_02184__PTR131), .S(_02959__PTR31), .Z(_02288__PTR3) );
  MUX2_X1 U8399 ( .A(_03191__PTR4), .B(_02184__PTR132), .S(_02959__PTR31), .Z(_02288__PTR4) );
  MUX2_X1 U8400 ( .A(_03191__PTR5), .B(_02184__PTR133), .S(_02959__PTR31), .Z(_02288__PTR5) );
  MUX2_X1 U8401 ( .A(_03191__PTR6), .B(_02184__PTR134), .S(_02959__PTR31), .Z(_02288__PTR6) );
  MUX2_X1 U8402 ( .A(_03191__PTR7), .B(_02184__PTR135), .S(_02959__PTR31), .Z(_02288__PTR7) );
  MUX2_X1 U8403 ( .A(_03191__PTR8), .B(_02184__PTR136), .S(_02959__PTR31), .Z(_02288__PTR8) );
  MUX2_X1 U8404 ( .A(_03191__PTR9), .B(_02184__PTR137), .S(_02959__PTR31), .Z(_02288__PTR9) );
  MUX2_X1 U8405 ( .A(_03191__PTR10), .B(_02184__PTR138), .S(_02959__PTR31), .Z(_02288__PTR10) );
  MUX2_X1 U8406 ( .A(_03191__PTR11), .B(_02184__PTR139), .S(_02959__PTR31), .Z(_02288__PTR11) );
  MUX2_X1 U8407 ( .A(_03191__PTR12), .B(_02184__PTR140), .S(_02959__PTR31), .Z(_02288__PTR12) );
  MUX2_X1 U8408 ( .A(_03191__PTR13), .B(_02184__PTR141), .S(_02959__PTR31), .Z(_02288__PTR13) );
  MUX2_X1 U8409 ( .A(_03191__PTR14), .B(_02184__PTR142), .S(_02959__PTR31), .Z(_02288__PTR14) );
  MUX2_X1 U8410 ( .A(_03191__PTR15), .B(_02184__PTR143), .S(_02959__PTR31), .Z(_02288__PTR15) );
  MUX2_X1 U8411 ( .A(_03191__PTR16), .B(_02184__PTR144), .S(_02959__PTR31), .Z(_02288__PTR16) );
  MUX2_X1 U8412 ( .A(_03191__PTR17), .B(_02184__PTR145), .S(_02959__PTR31), .Z(_02288__PTR17) );
  MUX2_X1 U8413 ( .A(_03191__PTR18), .B(_02184__PTR146), .S(_02959__PTR31), .Z(_02288__PTR18) );
  MUX2_X1 U8414 ( .A(_03191__PTR19), .B(_02184__PTR147), .S(_02959__PTR31), .Z(_02288__PTR19) );
  MUX2_X1 U8415 ( .A(_03191__PTR20), .B(_02184__PTR148), .S(_02959__PTR31), .Z(_02288__PTR20) );
  MUX2_X1 U8416 ( .A(_03191__PTR21), .B(_02184__PTR149), .S(_02959__PTR31), .Z(_02288__PTR21) );
  MUX2_X1 U8417 ( .A(_03191__PTR22), .B(_02184__PTR150), .S(_02959__PTR31), .Z(_02288__PTR22) );
  MUX2_X1 U8418 ( .A(_03191__PTR23), .B(_02184__PTR151), .S(_02959__PTR31), .Z(_02288__PTR23) );
  MUX2_X1 U8419 ( .A(_03191__PTR24), .B(_02184__PTR152), .S(_02959__PTR31), .Z(_02288__PTR24) );
  MUX2_X1 U8420 ( .A(_03191__PTR25), .B(_02184__PTR153), .S(_02959__PTR31), .Z(_02288__PTR25) );
  MUX2_X1 U8421 ( .A(_03191__PTR26), .B(_02184__PTR154), .S(_02959__PTR31), .Z(_02288__PTR26) );
  MUX2_X1 U8422 ( .A(_03191__PTR27), .B(_02184__PTR155), .S(_02959__PTR31), .Z(_02288__PTR27) );
  MUX2_X1 U8423 ( .A(_03191__PTR28), .B(_02184__PTR156), .S(_02959__PTR31), .Z(_02288__PTR28) );
  MUX2_X1 U8424 ( .A(_03191__PTR29), .B(_02184__PTR157), .S(_02959__PTR31), .Z(_02288__PTR29) );
  MUX2_X1 U8425 ( .A(_03191__PTR30), .B(_02184__PTR158), .S(_02959__PTR31), .Z(_02288__PTR30) );
  MUX2_X1 U8426 ( .A(_03191__PTR31), .B(_02184__PTR159), .S(_02959__PTR31), .Z(_02288__PTR31) );
  MUX2_X1 U8427 ( .A(_02270__PTR0), .B(_03033__PTR0), .S(_02134__PTR0), .Z(_02287__PTR0) );
  MUX2_X1 U8428 ( .A(_02270__PTR1), .B(_03034__PTR1), .S(_02134__PTR0), .Z(_02287__PTR1) );
  MUX2_X1 U8429 ( .A(_02270__PTR2), .B(_03034__PTR2), .S(_02134__PTR0), .Z(_02287__PTR2) );
  MUX2_X1 U8430 ( .A(_02270__PTR3), .B(_03034__PTR3), .S(_02134__PTR0), .Z(_02287__PTR3) );
  MUX2_X1 U8431 ( .A(_02270__PTR4), .B(_03034__PTR4), .S(_02134__PTR0), .Z(_02287__PTR4) );
  MUX2_X1 U8432 ( .A(_02270__PTR5), .B(_03034__PTR5), .S(_02134__PTR0), .Z(_02287__PTR5) );
  MUX2_X1 U8433 ( .A(_02270__PTR6), .B(_03034__PTR6), .S(_02134__PTR0), .Z(_02287__PTR6) );
  MUX2_X1 U8434 ( .A(_02270__PTR7), .B(_03034__PTR7), .S(_02134__PTR0), .Z(_02287__PTR7) );
  MUX2_X1 U8435 ( .A(_02269__PTR0), .B(_03033__PTR0), .S(_02134__PTR1), .Z(_02286__PTR0) );
  MUX2_X1 U8436 ( .A(_02269__PTR1), .B(_03034__PTR1), .S(_02134__PTR1), .Z(_02286__PTR1) );
  MUX2_X1 U8437 ( .A(_02269__PTR2), .B(_03034__PTR2), .S(_02134__PTR1), .Z(_02286__PTR2) );
  MUX2_X1 U8438 ( .A(_02269__PTR3), .B(_03034__PTR3), .S(_02134__PTR1), .Z(_02286__PTR3) );
  MUX2_X1 U8439 ( .A(_02269__PTR4), .B(_03034__PTR4), .S(_02134__PTR1), .Z(_02286__PTR4) );
  MUX2_X1 U8440 ( .A(_02269__PTR5), .B(_03034__PTR5), .S(_02134__PTR1), .Z(_02286__PTR5) );
  MUX2_X1 U8441 ( .A(_02269__PTR6), .B(_03034__PTR6), .S(_02134__PTR1), .Z(_02286__PTR6) );
  MUX2_X1 U8442 ( .A(_02269__PTR7), .B(_03034__PTR7), .S(_02134__PTR1), .Z(_02286__PTR7) );
  MUX2_X1 U8443 ( .A(_02268__PTR0), .B(_03033__PTR0), .S(_02134__PTR2), .Z(_02285__PTR0) );
  MUX2_X1 U8444 ( .A(_02268__PTR1), .B(_03034__PTR1), .S(_02134__PTR2), .Z(_02285__PTR1) );
  MUX2_X1 U8445 ( .A(_02268__PTR2), .B(_03034__PTR2), .S(_02134__PTR2), .Z(_02285__PTR2) );
  MUX2_X1 U8446 ( .A(_02268__PTR3), .B(_03034__PTR3), .S(_02134__PTR2), .Z(_02285__PTR3) );
  MUX2_X1 U8447 ( .A(_02268__PTR4), .B(_03034__PTR4), .S(_02134__PTR2), .Z(_02285__PTR4) );
  MUX2_X1 U8448 ( .A(_02268__PTR5), .B(_03034__PTR5), .S(_02134__PTR2), .Z(_02285__PTR5) );
  MUX2_X1 U8449 ( .A(_02268__PTR6), .B(_03034__PTR6), .S(_02134__PTR2), .Z(_02285__PTR6) );
  MUX2_X1 U8450 ( .A(_02268__PTR7), .B(_03034__PTR7), .S(_02134__PTR2), .Z(_02285__PTR7) );
  MUX2_X1 U8451 ( .A(_02267__PTR0), .B(_03033__PTR0), .S(_02134__PTR3), .Z(_02284__PTR0) );
  MUX2_X1 U8452 ( .A(_02267__PTR1), .B(_03034__PTR1), .S(_02134__PTR3), .Z(_02284__PTR1) );
  MUX2_X1 U8453 ( .A(_02267__PTR2), .B(_03034__PTR2), .S(_02134__PTR3), .Z(_02284__PTR2) );
  MUX2_X1 U8454 ( .A(_02267__PTR3), .B(_03034__PTR3), .S(_02134__PTR3), .Z(_02284__PTR3) );
  MUX2_X1 U8455 ( .A(_02267__PTR4), .B(_03034__PTR4), .S(_02134__PTR3), .Z(_02284__PTR4) );
  MUX2_X1 U8456 ( .A(_02267__PTR5), .B(_03034__PTR5), .S(_02134__PTR3), .Z(_02284__PTR5) );
  MUX2_X1 U8457 ( .A(_02267__PTR6), .B(_03034__PTR6), .S(_02134__PTR3), .Z(_02284__PTR6) );
  MUX2_X1 U8458 ( .A(_02267__PTR7), .B(_03034__PTR7), .S(_02134__PTR3), .Z(_02284__PTR7) );
  MUX2_X1 U8459 ( .A(_02266__PTR0), .B(_03033__PTR0), .S(_02134__PTR4), .Z(_02283__PTR0) );
  MUX2_X1 U8460 ( .A(_02266__PTR1), .B(_03034__PTR1), .S(_02134__PTR4), .Z(_02283__PTR1) );
  MUX2_X1 U8461 ( .A(_02266__PTR2), .B(_03034__PTR2), .S(_02134__PTR4), .Z(_02283__PTR2) );
  MUX2_X1 U8462 ( .A(_02266__PTR3), .B(_03034__PTR3), .S(_02134__PTR4), .Z(_02283__PTR3) );
  MUX2_X1 U8463 ( .A(_02266__PTR4), .B(_03034__PTR4), .S(_02134__PTR4), .Z(_02283__PTR4) );
  MUX2_X1 U8464 ( .A(_02266__PTR5), .B(_03034__PTR5), .S(_02134__PTR4), .Z(_02283__PTR5) );
  MUX2_X1 U8465 ( .A(_02266__PTR6), .B(_03034__PTR6), .S(_02134__PTR4), .Z(_02283__PTR6) );
  MUX2_X1 U8466 ( .A(_02266__PTR7), .B(_03034__PTR7), .S(_02134__PTR4), .Z(_02283__PTR7) );
  MUX2_X1 U8467 ( .A(_02265__PTR0), .B(_03033__PTR0), .S(_02134__PTR5), .Z(_02282__PTR0) );
  MUX2_X1 U8468 ( .A(_02265__PTR1), .B(_03034__PTR1), .S(_02134__PTR5), .Z(_02282__PTR1) );
  MUX2_X1 U8469 ( .A(_02265__PTR2), .B(_03034__PTR2), .S(_02134__PTR5), .Z(_02282__PTR2) );
  MUX2_X1 U8470 ( .A(_02265__PTR3), .B(_03034__PTR3), .S(_02134__PTR5), .Z(_02282__PTR3) );
  MUX2_X1 U8471 ( .A(_02265__PTR4), .B(_03034__PTR4), .S(_02134__PTR5), .Z(_02282__PTR4) );
  MUX2_X1 U8472 ( .A(_02265__PTR5), .B(_03034__PTR5), .S(_02134__PTR5), .Z(_02282__PTR5) );
  MUX2_X1 U8473 ( .A(_02265__PTR6), .B(_03034__PTR6), .S(_02134__PTR5), .Z(_02282__PTR6) );
  MUX2_X1 U8474 ( .A(_02265__PTR7), .B(_03034__PTR7), .S(_02134__PTR5), .Z(_02282__PTR7) );
  MUX2_X1 U8475 ( .A(_02264__PTR0), .B(_03033__PTR0), .S(_02134__PTR6), .Z(_02281__PTR0) );
  MUX2_X1 U8476 ( .A(_02264__PTR1), .B(_03034__PTR1), .S(_02134__PTR6), .Z(_02281__PTR1) );
  MUX2_X1 U8477 ( .A(_02264__PTR2), .B(_03034__PTR2), .S(_02134__PTR6), .Z(_02281__PTR2) );
  MUX2_X1 U8478 ( .A(_02264__PTR3), .B(_03034__PTR3), .S(_02134__PTR6), .Z(_02281__PTR3) );
  MUX2_X1 U8479 ( .A(_02264__PTR4), .B(_03034__PTR4), .S(_02134__PTR6), .Z(_02281__PTR4) );
  MUX2_X1 U8480 ( .A(_02264__PTR5), .B(_03034__PTR5), .S(_02134__PTR6), .Z(_02281__PTR5) );
  MUX2_X1 U8481 ( .A(_02264__PTR6), .B(_03034__PTR6), .S(_02134__PTR6), .Z(_02281__PTR6) );
  MUX2_X1 U8482 ( .A(_02264__PTR7), .B(_03034__PTR7), .S(_02134__PTR6), .Z(_02281__PTR7) );
  MUX2_X1 U8483 ( .A(_02263__PTR0), .B(_03033__PTR0), .S(_02134__PTR7), .Z(_02280__PTR0) );
  MUX2_X1 U8484 ( .A(_02263__PTR1), .B(_03034__PTR1), .S(_02134__PTR7), .Z(_02280__PTR1) );
  MUX2_X1 U8485 ( .A(_02263__PTR2), .B(_03034__PTR2), .S(_02134__PTR7), .Z(_02280__PTR2) );
  MUX2_X1 U8486 ( .A(_02263__PTR3), .B(_03034__PTR3), .S(_02134__PTR7), .Z(_02280__PTR3) );
  MUX2_X1 U8487 ( .A(_02263__PTR4), .B(_03034__PTR4), .S(_02134__PTR7), .Z(_02280__PTR4) );
  MUX2_X1 U8488 ( .A(_02263__PTR5), .B(_03034__PTR5), .S(_02134__PTR7), .Z(_02280__PTR5) );
  MUX2_X1 U8489 ( .A(_02263__PTR6), .B(_03034__PTR6), .S(_02134__PTR7), .Z(_02280__PTR6) );
  MUX2_X1 U8490 ( .A(_02263__PTR7), .B(_03034__PTR7), .S(_02134__PTR7), .Z(_02280__PTR7) );
  MUX2_X1 U8491 ( .A(_02262__PTR0), .B(_03033__PTR0), .S(_02134__PTR8), .Z(_02279__PTR0) );
  MUX2_X1 U8492 ( .A(_02262__PTR1), .B(_03034__PTR1), .S(_02134__PTR8), .Z(_02279__PTR1) );
  MUX2_X1 U8493 ( .A(_02262__PTR2), .B(_03034__PTR2), .S(_02134__PTR8), .Z(_02279__PTR2) );
  MUX2_X1 U8494 ( .A(_02262__PTR3), .B(_03034__PTR3), .S(_02134__PTR8), .Z(_02279__PTR3) );
  MUX2_X1 U8495 ( .A(_02262__PTR4), .B(_03034__PTR4), .S(_02134__PTR8), .Z(_02279__PTR4) );
  MUX2_X1 U8496 ( .A(_02262__PTR5), .B(_03034__PTR5), .S(_02134__PTR8), .Z(_02279__PTR5) );
  MUX2_X1 U8497 ( .A(_02262__PTR6), .B(_03034__PTR6), .S(_02134__PTR8), .Z(_02279__PTR6) );
  MUX2_X1 U8498 ( .A(_02262__PTR7), .B(_03034__PTR7), .S(_02134__PTR8), .Z(_02279__PTR7) );
  MUX2_X1 U8499 ( .A(_02261__PTR0), .B(_03033__PTR0), .S(_02134__PTR9), .Z(_02278__PTR0) );
  MUX2_X1 U8500 ( .A(_02261__PTR1), .B(_03034__PTR1), .S(_02134__PTR9), .Z(_02278__PTR1) );
  MUX2_X1 U8501 ( .A(_02261__PTR2), .B(_03034__PTR2), .S(_02134__PTR9), .Z(_02278__PTR2) );
  MUX2_X1 U8502 ( .A(_02261__PTR3), .B(_03034__PTR3), .S(_02134__PTR9), .Z(_02278__PTR3) );
  MUX2_X1 U8503 ( .A(_02261__PTR4), .B(_03034__PTR4), .S(_02134__PTR9), .Z(_02278__PTR4) );
  MUX2_X1 U8504 ( .A(_02261__PTR5), .B(_03034__PTR5), .S(_02134__PTR9), .Z(_02278__PTR5) );
  MUX2_X1 U8505 ( .A(_02261__PTR6), .B(_03034__PTR6), .S(_02134__PTR9), .Z(_02278__PTR6) );
  MUX2_X1 U8506 ( .A(_02261__PTR7), .B(_03034__PTR7), .S(_02134__PTR9), .Z(_02278__PTR7) );
  MUX2_X1 U8507 ( .A(_02260__PTR0), .B(_03033__PTR0), .S(_02134__PTR10), .Z(_02277__PTR0) );
  MUX2_X1 U8508 ( .A(_02260__PTR1), .B(_03034__PTR1), .S(_02134__PTR10), .Z(_02277__PTR1) );
  MUX2_X1 U8509 ( .A(_02260__PTR2), .B(_03034__PTR2), .S(_02134__PTR10), .Z(_02277__PTR2) );
  MUX2_X1 U8510 ( .A(_02260__PTR3), .B(_03034__PTR3), .S(_02134__PTR10), .Z(_02277__PTR3) );
  MUX2_X1 U8511 ( .A(_02260__PTR4), .B(_03034__PTR4), .S(_02134__PTR10), .Z(_02277__PTR4) );
  MUX2_X1 U8512 ( .A(_02260__PTR5), .B(_03034__PTR5), .S(_02134__PTR10), .Z(_02277__PTR5) );
  MUX2_X1 U8513 ( .A(_02260__PTR6), .B(_03034__PTR6), .S(_02134__PTR10), .Z(_02277__PTR6) );
  MUX2_X1 U8514 ( .A(_02260__PTR7), .B(_03034__PTR7), .S(_02134__PTR10), .Z(_02277__PTR7) );
  MUX2_X1 U8515 ( .A(_02259__PTR0), .B(_03033__PTR0), .S(_02134__PTR11), .Z(_02276__PTR0) );
  MUX2_X1 U8516 ( .A(_02259__PTR1), .B(_03034__PTR1), .S(_02134__PTR11), .Z(_02276__PTR1) );
  MUX2_X1 U8517 ( .A(_02259__PTR2), .B(_03034__PTR2), .S(_02134__PTR11), .Z(_02276__PTR2) );
  MUX2_X1 U8518 ( .A(_02259__PTR3), .B(_03034__PTR3), .S(_02134__PTR11), .Z(_02276__PTR3) );
  MUX2_X1 U8519 ( .A(_02259__PTR4), .B(_03034__PTR4), .S(_02134__PTR11), .Z(_02276__PTR4) );
  MUX2_X1 U8520 ( .A(_02259__PTR5), .B(_03034__PTR5), .S(_02134__PTR11), .Z(_02276__PTR5) );
  MUX2_X1 U8521 ( .A(_02259__PTR6), .B(_03034__PTR6), .S(_02134__PTR11), .Z(_02276__PTR6) );
  MUX2_X1 U8522 ( .A(_02259__PTR7), .B(_03034__PTR7), .S(_02134__PTR11), .Z(_02276__PTR7) );
  MUX2_X1 U8523 ( .A(_02258__PTR0), .B(_03033__PTR0), .S(_02134__PTR12), .Z(_02275__PTR0) );
  MUX2_X1 U8524 ( .A(_02258__PTR1), .B(_03034__PTR1), .S(_02134__PTR12), .Z(_02275__PTR1) );
  MUX2_X1 U8525 ( .A(_02258__PTR2), .B(_03034__PTR2), .S(_02134__PTR12), .Z(_02275__PTR2) );
  MUX2_X1 U8526 ( .A(_02258__PTR3), .B(_03034__PTR3), .S(_02134__PTR12), .Z(_02275__PTR3) );
  MUX2_X1 U8527 ( .A(_02258__PTR4), .B(_03034__PTR4), .S(_02134__PTR12), .Z(_02275__PTR4) );
  MUX2_X1 U8528 ( .A(_02258__PTR5), .B(_03034__PTR5), .S(_02134__PTR12), .Z(_02275__PTR5) );
  MUX2_X1 U8529 ( .A(_02258__PTR6), .B(_03034__PTR6), .S(_02134__PTR12), .Z(_02275__PTR6) );
  MUX2_X1 U8530 ( .A(_02258__PTR7), .B(_03034__PTR7), .S(_02134__PTR12), .Z(_02275__PTR7) );
  MUX2_X1 U8531 ( .A(_02257__PTR0), .B(_03033__PTR0), .S(_02134__PTR13), .Z(_02274__PTR0) );
  MUX2_X1 U8532 ( .A(_02257__PTR1), .B(_03034__PTR1), .S(_02134__PTR13), .Z(_02274__PTR1) );
  MUX2_X1 U8533 ( .A(_02257__PTR2), .B(_03034__PTR2), .S(_02134__PTR13), .Z(_02274__PTR2) );
  MUX2_X1 U8534 ( .A(_02257__PTR3), .B(_03034__PTR3), .S(_02134__PTR13), .Z(_02274__PTR3) );
  MUX2_X1 U8535 ( .A(_02257__PTR4), .B(_03034__PTR4), .S(_02134__PTR13), .Z(_02274__PTR4) );
  MUX2_X1 U8536 ( .A(_02257__PTR5), .B(_03034__PTR5), .S(_02134__PTR13), .Z(_02274__PTR5) );
  MUX2_X1 U8537 ( .A(_02257__PTR6), .B(_03034__PTR6), .S(_02134__PTR13), .Z(_02274__PTR6) );
  MUX2_X1 U8538 ( .A(_02257__PTR7), .B(_03034__PTR7), .S(_02134__PTR13), .Z(_02274__PTR7) );
  MUX2_X1 U8539 ( .A(_02256__PTR0), .B(_03033__PTR0), .S(_02134__PTR14), .Z(_02273__PTR0) );
  MUX2_X1 U8540 ( .A(_02256__PTR1), .B(_03034__PTR1), .S(_02134__PTR14), .Z(_02273__PTR1) );
  MUX2_X1 U8541 ( .A(_02256__PTR2), .B(_03034__PTR2), .S(_02134__PTR14), .Z(_02273__PTR2) );
  MUX2_X1 U8542 ( .A(_02256__PTR3), .B(_03034__PTR3), .S(_02134__PTR14), .Z(_02273__PTR3) );
  MUX2_X1 U8543 ( .A(_02256__PTR4), .B(_03034__PTR4), .S(_02134__PTR14), .Z(_02273__PTR4) );
  MUX2_X1 U8544 ( .A(_02256__PTR5), .B(_03034__PTR5), .S(_02134__PTR14), .Z(_02273__PTR5) );
  MUX2_X1 U8545 ( .A(_02256__PTR6), .B(_03034__PTR6), .S(_02134__PTR14), .Z(_02273__PTR6) );
  MUX2_X1 U8546 ( .A(_02256__PTR7), .B(_03034__PTR7), .S(_02134__PTR14), .Z(_02273__PTR7) );
  MUX2_X1 U8547 ( .A(_02255__PTR0), .B(_03033__PTR0), .S(_02134__PTR15), .Z(_02272__PTR0) );
  MUX2_X1 U8548 ( .A(_02255__PTR1), .B(_03034__PTR1), .S(_02134__PTR15), .Z(_02272__PTR1) );
  MUX2_X1 U8549 ( .A(_02255__PTR2), .B(_03034__PTR2), .S(_02134__PTR15), .Z(_02272__PTR2) );
  MUX2_X1 U8550 ( .A(_02255__PTR3), .B(_03034__PTR3), .S(_02134__PTR15), .Z(_02272__PTR3) );
  MUX2_X1 U8551 ( .A(_02255__PTR4), .B(_03034__PTR4), .S(_02134__PTR15), .Z(_02272__PTR4) );
  MUX2_X1 U8552 ( .A(_02255__PTR5), .B(_03034__PTR5), .S(_02134__PTR15), .Z(_02272__PTR5) );
  MUX2_X1 U8553 ( .A(_02255__PTR6), .B(_03034__PTR6), .S(_02134__PTR15), .Z(_02272__PTR6) );
  MUX2_X1 U8554 ( .A(_02255__PTR7), .B(_03034__PTR7), .S(_02134__PTR15), .Z(_02272__PTR7) );
  MUX2_X1 U8555 ( .A(_02220__PTR32), .B(_03028__PTR0), .S(_02132__PTR0), .Z(_02270__PTR0) );
  MUX2_X1 U8556 ( .A(_02220__PTR33), .B(_03029__PTR1), .S(_02132__PTR0), .Z(_02270__PTR1) );
  MUX2_X1 U8557 ( .A(_02220__PTR34), .B(_03029__PTR2), .S(_02132__PTR0), .Z(_02270__PTR2) );
  MUX2_X1 U8558 ( .A(_02220__PTR35), .B(_03029__PTR3), .S(_02132__PTR0), .Z(_02270__PTR3) );
  MUX2_X1 U8559 ( .A(_02220__PTR36), .B(_03029__PTR4), .S(_02132__PTR0), .Z(_02270__PTR4) );
  MUX2_X1 U8560 ( .A(_02220__PTR37), .B(_03029__PTR5), .S(_02132__PTR0), .Z(_02270__PTR5) );
  MUX2_X1 U8561 ( .A(_02220__PTR38), .B(_03029__PTR6), .S(_02132__PTR0), .Z(_02270__PTR6) );
  MUX2_X1 U8562 ( .A(_02220__PTR39), .B(_03029__PTR7), .S(_02132__PTR0), .Z(_02270__PTR7) );
  MUX2_X1 U8563 ( .A(_02218__PTR32), .B(_03028__PTR0), .S(_02132__PTR1), .Z(_02269__PTR0) );
  MUX2_X1 U8564 ( .A(_02218__PTR33), .B(_03029__PTR1), .S(_02132__PTR1), .Z(_02269__PTR1) );
  MUX2_X1 U8565 ( .A(_02218__PTR34), .B(_03029__PTR2), .S(_02132__PTR1), .Z(_02269__PTR2) );
  MUX2_X1 U8566 ( .A(_02218__PTR35), .B(_03029__PTR3), .S(_02132__PTR1), .Z(_02269__PTR3) );
  MUX2_X1 U8567 ( .A(_02218__PTR36), .B(_03029__PTR4), .S(_02132__PTR1), .Z(_02269__PTR4) );
  MUX2_X1 U8568 ( .A(_02218__PTR37), .B(_03029__PTR5), .S(_02132__PTR1), .Z(_02269__PTR5) );
  MUX2_X1 U8569 ( .A(_02218__PTR38), .B(_03029__PTR6), .S(_02132__PTR1), .Z(_02269__PTR6) );
  MUX2_X1 U8570 ( .A(_02218__PTR39), .B(_03029__PTR7), .S(_02132__PTR1), .Z(_02269__PTR7) );
  MUX2_X1 U8571 ( .A(_02216__PTR32), .B(_03028__PTR0), .S(_02132__PTR2), .Z(_02268__PTR0) );
  MUX2_X1 U8572 ( .A(_02216__PTR33), .B(_03029__PTR1), .S(_02132__PTR2), .Z(_02268__PTR1) );
  MUX2_X1 U8573 ( .A(_02216__PTR34), .B(_03029__PTR2), .S(_02132__PTR2), .Z(_02268__PTR2) );
  MUX2_X1 U8574 ( .A(_02216__PTR35), .B(_03029__PTR3), .S(_02132__PTR2), .Z(_02268__PTR3) );
  MUX2_X1 U8575 ( .A(_02216__PTR36), .B(_03029__PTR4), .S(_02132__PTR2), .Z(_02268__PTR4) );
  MUX2_X1 U8576 ( .A(_02216__PTR37), .B(_03029__PTR5), .S(_02132__PTR2), .Z(_02268__PTR5) );
  MUX2_X1 U8577 ( .A(_02216__PTR38), .B(_03029__PTR6), .S(_02132__PTR2), .Z(_02268__PTR6) );
  MUX2_X1 U8578 ( .A(_02216__PTR39), .B(_03029__PTR7), .S(_02132__PTR2), .Z(_02268__PTR7) );
  MUX2_X1 U8579 ( .A(_02214__PTR32), .B(_03028__PTR0), .S(_02132__PTR3), .Z(_02267__PTR0) );
  MUX2_X1 U8580 ( .A(_02214__PTR33), .B(_03029__PTR1), .S(_02132__PTR3), .Z(_02267__PTR1) );
  MUX2_X1 U8581 ( .A(_02214__PTR34), .B(_03029__PTR2), .S(_02132__PTR3), .Z(_02267__PTR2) );
  MUX2_X1 U8582 ( .A(_02214__PTR35), .B(_03029__PTR3), .S(_02132__PTR3), .Z(_02267__PTR3) );
  MUX2_X1 U8583 ( .A(_02214__PTR36), .B(_03029__PTR4), .S(_02132__PTR3), .Z(_02267__PTR4) );
  MUX2_X1 U8584 ( .A(_02214__PTR37), .B(_03029__PTR5), .S(_02132__PTR3), .Z(_02267__PTR5) );
  MUX2_X1 U8585 ( .A(_02214__PTR38), .B(_03029__PTR6), .S(_02132__PTR3), .Z(_02267__PTR6) );
  MUX2_X1 U8586 ( .A(_02214__PTR39), .B(_03029__PTR7), .S(_02132__PTR3), .Z(_02267__PTR7) );
  MUX2_X1 U8587 ( .A(_02212__PTR32), .B(_03028__PTR0), .S(_02132__PTR4), .Z(_02266__PTR0) );
  MUX2_X1 U8588 ( .A(_02212__PTR33), .B(_03029__PTR1), .S(_02132__PTR4), .Z(_02266__PTR1) );
  MUX2_X1 U8589 ( .A(_02212__PTR34), .B(_03029__PTR2), .S(_02132__PTR4), .Z(_02266__PTR2) );
  MUX2_X1 U8590 ( .A(_02212__PTR35), .B(_03029__PTR3), .S(_02132__PTR4), .Z(_02266__PTR3) );
  MUX2_X1 U8591 ( .A(_02212__PTR36), .B(_03029__PTR4), .S(_02132__PTR4), .Z(_02266__PTR4) );
  MUX2_X1 U8592 ( .A(_02212__PTR37), .B(_03029__PTR5), .S(_02132__PTR4), .Z(_02266__PTR5) );
  MUX2_X1 U8593 ( .A(_02212__PTR38), .B(_03029__PTR6), .S(_02132__PTR4), .Z(_02266__PTR6) );
  MUX2_X1 U8594 ( .A(_02212__PTR39), .B(_03029__PTR7), .S(_02132__PTR4), .Z(_02266__PTR7) );
  MUX2_X1 U8595 ( .A(_02210__PTR32), .B(_03028__PTR0), .S(_02132__PTR5), .Z(_02265__PTR0) );
  MUX2_X1 U8596 ( .A(_02210__PTR33), .B(_03029__PTR1), .S(_02132__PTR5), .Z(_02265__PTR1) );
  MUX2_X1 U8597 ( .A(_02210__PTR34), .B(_03029__PTR2), .S(_02132__PTR5), .Z(_02265__PTR2) );
  MUX2_X1 U8598 ( .A(_02210__PTR35), .B(_03029__PTR3), .S(_02132__PTR5), .Z(_02265__PTR3) );
  MUX2_X1 U8599 ( .A(_02210__PTR36), .B(_03029__PTR4), .S(_02132__PTR5), .Z(_02265__PTR4) );
  MUX2_X1 U8600 ( .A(_02210__PTR37), .B(_03029__PTR5), .S(_02132__PTR5), .Z(_02265__PTR5) );
  MUX2_X1 U8601 ( .A(_02210__PTR38), .B(_03029__PTR6), .S(_02132__PTR5), .Z(_02265__PTR6) );
  MUX2_X1 U8602 ( .A(_02210__PTR39), .B(_03029__PTR7), .S(_02132__PTR5), .Z(_02265__PTR7) );
  MUX2_X1 U8603 ( .A(_02208__PTR32), .B(_03028__PTR0), .S(_02132__PTR6), .Z(_02264__PTR0) );
  MUX2_X1 U8604 ( .A(_02208__PTR33), .B(_03029__PTR1), .S(_02132__PTR6), .Z(_02264__PTR1) );
  MUX2_X1 U8605 ( .A(_02208__PTR34), .B(_03029__PTR2), .S(_02132__PTR6), .Z(_02264__PTR2) );
  MUX2_X1 U8606 ( .A(_02208__PTR35), .B(_03029__PTR3), .S(_02132__PTR6), .Z(_02264__PTR3) );
  MUX2_X1 U8607 ( .A(_02208__PTR36), .B(_03029__PTR4), .S(_02132__PTR6), .Z(_02264__PTR4) );
  MUX2_X1 U8608 ( .A(_02208__PTR37), .B(_03029__PTR5), .S(_02132__PTR6), .Z(_02264__PTR5) );
  MUX2_X1 U8609 ( .A(_02208__PTR38), .B(_03029__PTR6), .S(_02132__PTR6), .Z(_02264__PTR6) );
  MUX2_X1 U8610 ( .A(_02208__PTR39), .B(_03029__PTR7), .S(_02132__PTR6), .Z(_02264__PTR7) );
  MUX2_X1 U8611 ( .A(_02206__PTR32), .B(_03028__PTR0), .S(_02132__PTR7), .Z(_02263__PTR0) );
  MUX2_X1 U8612 ( .A(_02206__PTR33), .B(_03029__PTR1), .S(_02132__PTR7), .Z(_02263__PTR1) );
  MUX2_X1 U8613 ( .A(_02206__PTR34), .B(_03029__PTR2), .S(_02132__PTR7), .Z(_02263__PTR2) );
  MUX2_X1 U8614 ( .A(_02206__PTR35), .B(_03029__PTR3), .S(_02132__PTR7), .Z(_02263__PTR3) );
  MUX2_X1 U8615 ( .A(_02206__PTR36), .B(_03029__PTR4), .S(_02132__PTR7), .Z(_02263__PTR4) );
  MUX2_X1 U8616 ( .A(_02206__PTR37), .B(_03029__PTR5), .S(_02132__PTR7), .Z(_02263__PTR5) );
  MUX2_X1 U8617 ( .A(_02206__PTR38), .B(_03029__PTR6), .S(_02132__PTR7), .Z(_02263__PTR6) );
  MUX2_X1 U8618 ( .A(_02206__PTR39), .B(_03029__PTR7), .S(_02132__PTR7), .Z(_02263__PTR7) );
  MUX2_X1 U8619 ( .A(_02204__PTR32), .B(_03028__PTR0), .S(_02132__PTR8), .Z(_02262__PTR0) );
  MUX2_X1 U8620 ( .A(_02204__PTR33), .B(_03029__PTR1), .S(_02132__PTR8), .Z(_02262__PTR1) );
  MUX2_X1 U8621 ( .A(_02204__PTR34), .B(_03029__PTR2), .S(_02132__PTR8), .Z(_02262__PTR2) );
  MUX2_X1 U8622 ( .A(_02204__PTR35), .B(_03029__PTR3), .S(_02132__PTR8), .Z(_02262__PTR3) );
  MUX2_X1 U8623 ( .A(_02204__PTR36), .B(_03029__PTR4), .S(_02132__PTR8), .Z(_02262__PTR4) );
  MUX2_X1 U8624 ( .A(_02204__PTR37), .B(_03029__PTR5), .S(_02132__PTR8), .Z(_02262__PTR5) );
  MUX2_X1 U8625 ( .A(_02204__PTR38), .B(_03029__PTR6), .S(_02132__PTR8), .Z(_02262__PTR6) );
  MUX2_X1 U8626 ( .A(_02204__PTR39), .B(_03029__PTR7), .S(_02132__PTR8), .Z(_02262__PTR7) );
  MUX2_X1 U8627 ( .A(_02202__PTR32), .B(_03028__PTR0), .S(_02132__PTR9), .Z(_02261__PTR0) );
  MUX2_X1 U8628 ( .A(_02202__PTR33), .B(_03029__PTR1), .S(_02132__PTR9), .Z(_02261__PTR1) );
  MUX2_X1 U8629 ( .A(_02202__PTR34), .B(_03029__PTR2), .S(_02132__PTR9), .Z(_02261__PTR2) );
  MUX2_X1 U8630 ( .A(_02202__PTR35), .B(_03029__PTR3), .S(_02132__PTR9), .Z(_02261__PTR3) );
  MUX2_X1 U8631 ( .A(_02202__PTR36), .B(_03029__PTR4), .S(_02132__PTR9), .Z(_02261__PTR4) );
  MUX2_X1 U8632 ( .A(_02202__PTR37), .B(_03029__PTR5), .S(_02132__PTR9), .Z(_02261__PTR5) );
  MUX2_X1 U8633 ( .A(_02202__PTR38), .B(_03029__PTR6), .S(_02132__PTR9), .Z(_02261__PTR6) );
  MUX2_X1 U8634 ( .A(_02202__PTR39), .B(_03029__PTR7), .S(_02132__PTR9), .Z(_02261__PTR7) );
  MUX2_X1 U8635 ( .A(_02200__PTR32), .B(_03028__PTR0), .S(_02132__PTR10), .Z(_02260__PTR0) );
  MUX2_X1 U8636 ( .A(_02200__PTR33), .B(_03029__PTR1), .S(_02132__PTR10), .Z(_02260__PTR1) );
  MUX2_X1 U8637 ( .A(_02200__PTR34), .B(_03029__PTR2), .S(_02132__PTR10), .Z(_02260__PTR2) );
  MUX2_X1 U8638 ( .A(_02200__PTR35), .B(_03029__PTR3), .S(_02132__PTR10), .Z(_02260__PTR3) );
  MUX2_X1 U8639 ( .A(_02200__PTR36), .B(_03029__PTR4), .S(_02132__PTR10), .Z(_02260__PTR4) );
  MUX2_X1 U8640 ( .A(_02200__PTR37), .B(_03029__PTR5), .S(_02132__PTR10), .Z(_02260__PTR5) );
  MUX2_X1 U8641 ( .A(_02200__PTR38), .B(_03029__PTR6), .S(_02132__PTR10), .Z(_02260__PTR6) );
  MUX2_X1 U8642 ( .A(_02200__PTR39), .B(_03029__PTR7), .S(_02132__PTR10), .Z(_02260__PTR7) );
  MUX2_X1 U8643 ( .A(_02198__PTR32), .B(_03028__PTR0), .S(_02132__PTR11), .Z(_02259__PTR0) );
  MUX2_X1 U8644 ( .A(_02198__PTR33), .B(_03029__PTR1), .S(_02132__PTR11), .Z(_02259__PTR1) );
  MUX2_X1 U8645 ( .A(_02198__PTR34), .B(_03029__PTR2), .S(_02132__PTR11), .Z(_02259__PTR2) );
  MUX2_X1 U8646 ( .A(_02198__PTR35), .B(_03029__PTR3), .S(_02132__PTR11), .Z(_02259__PTR3) );
  MUX2_X1 U8647 ( .A(_02198__PTR36), .B(_03029__PTR4), .S(_02132__PTR11), .Z(_02259__PTR4) );
  MUX2_X1 U8648 ( .A(_02198__PTR37), .B(_03029__PTR5), .S(_02132__PTR11), .Z(_02259__PTR5) );
  MUX2_X1 U8649 ( .A(_02198__PTR38), .B(_03029__PTR6), .S(_02132__PTR11), .Z(_02259__PTR6) );
  MUX2_X1 U8650 ( .A(_02198__PTR39), .B(_03029__PTR7), .S(_02132__PTR11), .Z(_02259__PTR7) );
  MUX2_X1 U8651 ( .A(_02196__PTR32), .B(_03028__PTR0), .S(_02132__PTR12), .Z(_02258__PTR0) );
  MUX2_X1 U8652 ( .A(_02196__PTR33), .B(_03029__PTR1), .S(_02132__PTR12), .Z(_02258__PTR1) );
  MUX2_X1 U8653 ( .A(_02196__PTR34), .B(_03029__PTR2), .S(_02132__PTR12), .Z(_02258__PTR2) );
  MUX2_X1 U8654 ( .A(_02196__PTR35), .B(_03029__PTR3), .S(_02132__PTR12), .Z(_02258__PTR3) );
  MUX2_X1 U8655 ( .A(_02196__PTR36), .B(_03029__PTR4), .S(_02132__PTR12), .Z(_02258__PTR4) );
  MUX2_X1 U8656 ( .A(_02196__PTR37), .B(_03029__PTR5), .S(_02132__PTR12), .Z(_02258__PTR5) );
  MUX2_X1 U8657 ( .A(_02196__PTR38), .B(_03029__PTR6), .S(_02132__PTR12), .Z(_02258__PTR6) );
  MUX2_X1 U8658 ( .A(_02196__PTR39), .B(_03029__PTR7), .S(_02132__PTR12), .Z(_02258__PTR7) );
  MUX2_X1 U8659 ( .A(_02194__PTR32), .B(_03028__PTR0), .S(_02132__PTR13), .Z(_02257__PTR0) );
  MUX2_X1 U8660 ( .A(_02194__PTR33), .B(_03029__PTR1), .S(_02132__PTR13), .Z(_02257__PTR1) );
  MUX2_X1 U8661 ( .A(_02194__PTR34), .B(_03029__PTR2), .S(_02132__PTR13), .Z(_02257__PTR2) );
  MUX2_X1 U8662 ( .A(_02194__PTR35), .B(_03029__PTR3), .S(_02132__PTR13), .Z(_02257__PTR3) );
  MUX2_X1 U8663 ( .A(_02194__PTR36), .B(_03029__PTR4), .S(_02132__PTR13), .Z(_02257__PTR4) );
  MUX2_X1 U8664 ( .A(_02194__PTR37), .B(_03029__PTR5), .S(_02132__PTR13), .Z(_02257__PTR5) );
  MUX2_X1 U8665 ( .A(_02194__PTR38), .B(_03029__PTR6), .S(_02132__PTR13), .Z(_02257__PTR6) );
  MUX2_X1 U8666 ( .A(_02194__PTR39), .B(_03029__PTR7), .S(_02132__PTR13), .Z(_02257__PTR7) );
  MUX2_X1 U8667 ( .A(_02192__PTR32), .B(_03028__PTR0), .S(_02132__PTR14), .Z(_02256__PTR0) );
  MUX2_X1 U8668 ( .A(_02192__PTR33), .B(_03029__PTR1), .S(_02132__PTR14), .Z(_02256__PTR1) );
  MUX2_X1 U8669 ( .A(_02192__PTR34), .B(_03029__PTR2), .S(_02132__PTR14), .Z(_02256__PTR2) );
  MUX2_X1 U8670 ( .A(_02192__PTR35), .B(_03029__PTR3), .S(_02132__PTR14), .Z(_02256__PTR3) );
  MUX2_X1 U8671 ( .A(_02192__PTR36), .B(_03029__PTR4), .S(_02132__PTR14), .Z(_02256__PTR4) );
  MUX2_X1 U8672 ( .A(_02192__PTR37), .B(_03029__PTR5), .S(_02132__PTR14), .Z(_02256__PTR5) );
  MUX2_X1 U8673 ( .A(_02192__PTR38), .B(_03029__PTR6), .S(_02132__PTR14), .Z(_02256__PTR6) );
  MUX2_X1 U8674 ( .A(_02192__PTR39), .B(_03029__PTR7), .S(_02132__PTR14), .Z(_02256__PTR7) );
  MUX2_X1 U8675 ( .A(_02190__PTR32), .B(_03028__PTR0), .S(_02132__PTR15), .Z(_02255__PTR0) );
  MUX2_X1 U8676 ( .A(_02190__PTR33), .B(_03029__PTR1), .S(_02132__PTR15), .Z(_02255__PTR1) );
  MUX2_X1 U8677 ( .A(_02190__PTR34), .B(_03029__PTR2), .S(_02132__PTR15), .Z(_02255__PTR2) );
  MUX2_X1 U8678 ( .A(_02190__PTR35), .B(_03029__PTR3), .S(_02132__PTR15), .Z(_02255__PTR3) );
  MUX2_X1 U8679 ( .A(_02190__PTR36), .B(_03029__PTR4), .S(_02132__PTR15), .Z(_02255__PTR4) );
  MUX2_X1 U8680 ( .A(_02190__PTR37), .B(_03029__PTR5), .S(_02132__PTR15), .Z(_02255__PTR5) );
  MUX2_X1 U8681 ( .A(_02190__PTR38), .B(_03029__PTR6), .S(_02132__PTR15), .Z(_02255__PTR6) );
  MUX2_X1 U8682 ( .A(_02190__PTR39), .B(_03029__PTR7), .S(_02132__PTR15), .Z(_02255__PTR7) );
  MUX2_X1 U8683 ( .A(_02254__PTR0), .B(di2_PTR0), .S(_02130__PTR0), .Z(_02220__PTR32) );
  MUX2_X1 U8684 ( .A(_02254__PTR1), .B(di2_PTR1), .S(_02130__PTR0), .Z(_02220__PTR33) );
  MUX2_X1 U8685 ( .A(_02254__PTR2), .B(di2_PTR2), .S(_02130__PTR0), .Z(_02220__PTR34) );
  MUX2_X1 U8686 ( .A(_02254__PTR3), .B(di2_PTR3), .S(_02130__PTR0), .Z(_02220__PTR35) );
  MUX2_X1 U8687 ( .A(_02254__PTR4), .B(di2_PTR4), .S(_02130__PTR0), .Z(_02220__PTR36) );
  MUX2_X1 U8688 ( .A(_02254__PTR5), .B(di2_PTR5), .S(_02130__PTR0), .Z(_02220__PTR37) );
  MUX2_X1 U8689 ( .A(_02254__PTR6), .B(di2_PTR6), .S(_02130__PTR0), .Z(_02220__PTR38) );
  MUX2_X1 U8690 ( .A(_02254__PTR7), .B(di2_PTR7), .S(_02130__PTR0), .Z(_02220__PTR39) );
  MUX2_X1 U8691 ( .A(_02253__PTR0), .B(di2_PTR0), .S(_02130__PTR1), .Z(_02218__PTR32) );
  MUX2_X1 U8692 ( .A(_02253__PTR1), .B(di2_PTR1), .S(_02130__PTR1), .Z(_02218__PTR33) );
  MUX2_X1 U8693 ( .A(_02253__PTR2), .B(di2_PTR2), .S(_02130__PTR1), .Z(_02218__PTR34) );
  MUX2_X1 U8694 ( .A(_02253__PTR3), .B(di2_PTR3), .S(_02130__PTR1), .Z(_02218__PTR35) );
  MUX2_X1 U8695 ( .A(_02253__PTR4), .B(di2_PTR4), .S(_02130__PTR1), .Z(_02218__PTR36) );
  MUX2_X1 U8696 ( .A(_02253__PTR5), .B(di2_PTR5), .S(_02130__PTR1), .Z(_02218__PTR37) );
  MUX2_X1 U8697 ( .A(_02253__PTR6), .B(di2_PTR6), .S(_02130__PTR1), .Z(_02218__PTR38) );
  MUX2_X1 U8698 ( .A(_02253__PTR7), .B(di2_PTR7), .S(_02130__PTR1), .Z(_02218__PTR39) );
  MUX2_X1 U8699 ( .A(_02252__PTR0), .B(di2_PTR0), .S(_02130__PTR2), .Z(_02216__PTR32) );
  MUX2_X1 U8700 ( .A(_02252__PTR1), .B(di2_PTR1), .S(_02130__PTR2), .Z(_02216__PTR33) );
  MUX2_X1 U8701 ( .A(_02252__PTR2), .B(di2_PTR2), .S(_02130__PTR2), .Z(_02216__PTR34) );
  MUX2_X1 U8702 ( .A(_02252__PTR3), .B(di2_PTR3), .S(_02130__PTR2), .Z(_02216__PTR35) );
  MUX2_X1 U8703 ( .A(_02252__PTR4), .B(di2_PTR4), .S(_02130__PTR2), .Z(_02216__PTR36) );
  MUX2_X1 U8704 ( .A(_02252__PTR5), .B(di2_PTR5), .S(_02130__PTR2), .Z(_02216__PTR37) );
  MUX2_X1 U8705 ( .A(_02252__PTR6), .B(di2_PTR6), .S(_02130__PTR2), .Z(_02216__PTR38) );
  MUX2_X1 U8706 ( .A(_02252__PTR7), .B(di2_PTR7), .S(_02130__PTR2), .Z(_02216__PTR39) );
  MUX2_X1 U8707 ( .A(_02251__PTR0), .B(di2_PTR0), .S(_02130__PTR3), .Z(_02214__PTR32) );
  MUX2_X1 U8708 ( .A(_02251__PTR1), .B(di2_PTR1), .S(_02130__PTR3), .Z(_02214__PTR33) );
  MUX2_X1 U8709 ( .A(_02251__PTR2), .B(di2_PTR2), .S(_02130__PTR3), .Z(_02214__PTR34) );
  MUX2_X1 U8710 ( .A(_02251__PTR3), .B(di2_PTR3), .S(_02130__PTR3), .Z(_02214__PTR35) );
  MUX2_X1 U8711 ( .A(_02251__PTR4), .B(di2_PTR4), .S(_02130__PTR3), .Z(_02214__PTR36) );
  MUX2_X1 U8712 ( .A(_02251__PTR5), .B(di2_PTR5), .S(_02130__PTR3), .Z(_02214__PTR37) );
  MUX2_X1 U8713 ( .A(_02251__PTR6), .B(di2_PTR6), .S(_02130__PTR3), .Z(_02214__PTR38) );
  MUX2_X1 U8714 ( .A(_02251__PTR7), .B(di2_PTR7), .S(_02130__PTR3), .Z(_02214__PTR39) );
  MUX2_X1 U8715 ( .A(_02250__PTR0), .B(di2_PTR0), .S(_02130__PTR4), .Z(_02212__PTR32) );
  MUX2_X1 U8716 ( .A(_02250__PTR1), .B(di2_PTR1), .S(_02130__PTR4), .Z(_02212__PTR33) );
  MUX2_X1 U8717 ( .A(_02250__PTR2), .B(di2_PTR2), .S(_02130__PTR4), .Z(_02212__PTR34) );
  MUX2_X1 U8718 ( .A(_02250__PTR3), .B(di2_PTR3), .S(_02130__PTR4), .Z(_02212__PTR35) );
  MUX2_X1 U8719 ( .A(_02250__PTR4), .B(di2_PTR4), .S(_02130__PTR4), .Z(_02212__PTR36) );
  MUX2_X1 U8720 ( .A(_02250__PTR5), .B(di2_PTR5), .S(_02130__PTR4), .Z(_02212__PTR37) );
  MUX2_X1 U8721 ( .A(_02250__PTR6), .B(di2_PTR6), .S(_02130__PTR4), .Z(_02212__PTR38) );
  MUX2_X1 U8722 ( .A(_02250__PTR7), .B(di2_PTR7), .S(_02130__PTR4), .Z(_02212__PTR39) );
  MUX2_X1 U8723 ( .A(_02249__PTR0), .B(di2_PTR0), .S(_02130__PTR5), .Z(_02210__PTR32) );
  MUX2_X1 U8724 ( .A(_02249__PTR1), .B(di2_PTR1), .S(_02130__PTR5), .Z(_02210__PTR33) );
  MUX2_X1 U8725 ( .A(_02249__PTR2), .B(di2_PTR2), .S(_02130__PTR5), .Z(_02210__PTR34) );
  MUX2_X1 U8726 ( .A(_02249__PTR3), .B(di2_PTR3), .S(_02130__PTR5), .Z(_02210__PTR35) );
  MUX2_X1 U8727 ( .A(_02249__PTR4), .B(di2_PTR4), .S(_02130__PTR5), .Z(_02210__PTR36) );
  MUX2_X1 U8728 ( .A(_02249__PTR5), .B(di2_PTR5), .S(_02130__PTR5), .Z(_02210__PTR37) );
  MUX2_X1 U8729 ( .A(_02249__PTR6), .B(di2_PTR6), .S(_02130__PTR5), .Z(_02210__PTR38) );
  MUX2_X1 U8730 ( .A(_02249__PTR7), .B(di2_PTR7), .S(_02130__PTR5), .Z(_02210__PTR39) );
  MUX2_X1 U8731 ( .A(_02248__PTR0), .B(di2_PTR0), .S(_02130__PTR6), .Z(_02208__PTR32) );
  MUX2_X1 U8732 ( .A(_02248__PTR1), .B(di2_PTR1), .S(_02130__PTR6), .Z(_02208__PTR33) );
  MUX2_X1 U8733 ( .A(_02248__PTR2), .B(di2_PTR2), .S(_02130__PTR6), .Z(_02208__PTR34) );
  MUX2_X1 U8734 ( .A(_02248__PTR3), .B(di2_PTR3), .S(_02130__PTR6), .Z(_02208__PTR35) );
  MUX2_X1 U8735 ( .A(_02248__PTR4), .B(di2_PTR4), .S(_02130__PTR6), .Z(_02208__PTR36) );
  MUX2_X1 U8736 ( .A(_02248__PTR5), .B(di2_PTR5), .S(_02130__PTR6), .Z(_02208__PTR37) );
  MUX2_X1 U8737 ( .A(_02248__PTR6), .B(di2_PTR6), .S(_02130__PTR6), .Z(_02208__PTR38) );
  MUX2_X1 U8738 ( .A(_02248__PTR7), .B(di2_PTR7), .S(_02130__PTR6), .Z(_02208__PTR39) );
  MUX2_X1 U8739 ( .A(_02247__PTR0), .B(di2_PTR0), .S(_02130__PTR7), .Z(_02206__PTR32) );
  MUX2_X1 U8740 ( .A(_02247__PTR1), .B(di2_PTR1), .S(_02130__PTR7), .Z(_02206__PTR33) );
  MUX2_X1 U8741 ( .A(_02247__PTR2), .B(di2_PTR2), .S(_02130__PTR7), .Z(_02206__PTR34) );
  MUX2_X1 U8742 ( .A(_02247__PTR3), .B(di2_PTR3), .S(_02130__PTR7), .Z(_02206__PTR35) );
  MUX2_X1 U8743 ( .A(_02247__PTR4), .B(di2_PTR4), .S(_02130__PTR7), .Z(_02206__PTR36) );
  MUX2_X1 U8744 ( .A(_02247__PTR5), .B(di2_PTR5), .S(_02130__PTR7), .Z(_02206__PTR37) );
  MUX2_X1 U8745 ( .A(_02247__PTR6), .B(di2_PTR6), .S(_02130__PTR7), .Z(_02206__PTR38) );
  MUX2_X1 U8746 ( .A(_02247__PTR7), .B(di2_PTR7), .S(_02130__PTR7), .Z(_02206__PTR39) );
  MUX2_X1 U8747 ( .A(_02246__PTR0), .B(di2_PTR0), .S(_02130__PTR8), .Z(_02204__PTR32) );
  MUX2_X1 U8748 ( .A(_02246__PTR1), .B(di2_PTR1), .S(_02130__PTR8), .Z(_02204__PTR33) );
  MUX2_X1 U8749 ( .A(_02246__PTR2), .B(di2_PTR2), .S(_02130__PTR8), .Z(_02204__PTR34) );
  MUX2_X1 U8750 ( .A(_02246__PTR3), .B(di2_PTR3), .S(_02130__PTR8), .Z(_02204__PTR35) );
  MUX2_X1 U8751 ( .A(_02246__PTR4), .B(di2_PTR4), .S(_02130__PTR8), .Z(_02204__PTR36) );
  MUX2_X1 U8752 ( .A(_02246__PTR5), .B(di2_PTR5), .S(_02130__PTR8), .Z(_02204__PTR37) );
  MUX2_X1 U8753 ( .A(_02246__PTR6), .B(di2_PTR6), .S(_02130__PTR8), .Z(_02204__PTR38) );
  MUX2_X1 U8754 ( .A(_02246__PTR7), .B(di2_PTR7), .S(_02130__PTR8), .Z(_02204__PTR39) );
  MUX2_X1 U8755 ( .A(_02245__PTR0), .B(di2_PTR0), .S(_02130__PTR9), .Z(_02202__PTR32) );
  MUX2_X1 U8756 ( .A(_02245__PTR1), .B(di2_PTR1), .S(_02130__PTR9), .Z(_02202__PTR33) );
  MUX2_X1 U8757 ( .A(_02245__PTR2), .B(di2_PTR2), .S(_02130__PTR9), .Z(_02202__PTR34) );
  MUX2_X1 U8758 ( .A(_02245__PTR3), .B(di2_PTR3), .S(_02130__PTR9), .Z(_02202__PTR35) );
  MUX2_X1 U8759 ( .A(_02245__PTR4), .B(di2_PTR4), .S(_02130__PTR9), .Z(_02202__PTR36) );
  MUX2_X1 U8760 ( .A(_02245__PTR5), .B(di2_PTR5), .S(_02130__PTR9), .Z(_02202__PTR37) );
  MUX2_X1 U8761 ( .A(_02245__PTR6), .B(di2_PTR6), .S(_02130__PTR9), .Z(_02202__PTR38) );
  MUX2_X1 U8762 ( .A(_02245__PTR7), .B(di2_PTR7), .S(_02130__PTR9), .Z(_02202__PTR39) );
  MUX2_X1 U8763 ( .A(_02244__PTR0), .B(di2_PTR0), .S(_02130__PTR10), .Z(_02200__PTR32) );
  MUX2_X1 U8764 ( .A(_02244__PTR1), .B(di2_PTR1), .S(_02130__PTR10), .Z(_02200__PTR33) );
  MUX2_X1 U8765 ( .A(_02244__PTR2), .B(di2_PTR2), .S(_02130__PTR10), .Z(_02200__PTR34) );
  MUX2_X1 U8766 ( .A(_02244__PTR3), .B(di2_PTR3), .S(_02130__PTR10), .Z(_02200__PTR35) );
  MUX2_X1 U8767 ( .A(_02244__PTR4), .B(di2_PTR4), .S(_02130__PTR10), .Z(_02200__PTR36) );
  MUX2_X1 U8768 ( .A(_02244__PTR5), .B(di2_PTR5), .S(_02130__PTR10), .Z(_02200__PTR37) );
  MUX2_X1 U8769 ( .A(_02244__PTR6), .B(di2_PTR6), .S(_02130__PTR10), .Z(_02200__PTR38) );
  MUX2_X1 U8770 ( .A(_02244__PTR7), .B(di2_PTR7), .S(_02130__PTR10), .Z(_02200__PTR39) );
  MUX2_X1 U8771 ( .A(_02243__PTR0), .B(di2_PTR0), .S(_02130__PTR11), .Z(_02198__PTR32) );
  MUX2_X1 U8772 ( .A(_02243__PTR1), .B(di2_PTR1), .S(_02130__PTR11), .Z(_02198__PTR33) );
  MUX2_X1 U8773 ( .A(_02243__PTR2), .B(di2_PTR2), .S(_02130__PTR11), .Z(_02198__PTR34) );
  MUX2_X1 U8774 ( .A(_02243__PTR3), .B(di2_PTR3), .S(_02130__PTR11), .Z(_02198__PTR35) );
  MUX2_X1 U8775 ( .A(_02243__PTR4), .B(di2_PTR4), .S(_02130__PTR11), .Z(_02198__PTR36) );
  MUX2_X1 U8776 ( .A(_02243__PTR5), .B(di2_PTR5), .S(_02130__PTR11), .Z(_02198__PTR37) );
  MUX2_X1 U8777 ( .A(_02243__PTR6), .B(di2_PTR6), .S(_02130__PTR11), .Z(_02198__PTR38) );
  MUX2_X1 U8778 ( .A(_02243__PTR7), .B(di2_PTR7), .S(_02130__PTR11), .Z(_02198__PTR39) );
  MUX2_X1 U8779 ( .A(_02242__PTR0), .B(di2_PTR0), .S(_02130__PTR12), .Z(_02196__PTR32) );
  MUX2_X1 U8780 ( .A(_02242__PTR1), .B(di2_PTR1), .S(_02130__PTR12), .Z(_02196__PTR33) );
  MUX2_X1 U8781 ( .A(_02242__PTR2), .B(di2_PTR2), .S(_02130__PTR12), .Z(_02196__PTR34) );
  MUX2_X1 U8782 ( .A(_02242__PTR3), .B(di2_PTR3), .S(_02130__PTR12), .Z(_02196__PTR35) );
  MUX2_X1 U8783 ( .A(_02242__PTR4), .B(di2_PTR4), .S(_02130__PTR12), .Z(_02196__PTR36) );
  MUX2_X1 U8784 ( .A(_02242__PTR5), .B(di2_PTR5), .S(_02130__PTR12), .Z(_02196__PTR37) );
  MUX2_X1 U8785 ( .A(_02242__PTR6), .B(di2_PTR6), .S(_02130__PTR12), .Z(_02196__PTR38) );
  MUX2_X1 U8786 ( .A(_02242__PTR7), .B(di2_PTR7), .S(_02130__PTR12), .Z(_02196__PTR39) );
  MUX2_X1 U8787 ( .A(_02241__PTR0), .B(di2_PTR0), .S(_02130__PTR13), .Z(_02194__PTR32) );
  MUX2_X1 U8788 ( .A(_02241__PTR1), .B(di2_PTR1), .S(_02130__PTR13), .Z(_02194__PTR33) );
  MUX2_X1 U8789 ( .A(_02241__PTR2), .B(di2_PTR2), .S(_02130__PTR13), .Z(_02194__PTR34) );
  MUX2_X1 U8790 ( .A(_02241__PTR3), .B(di2_PTR3), .S(_02130__PTR13), .Z(_02194__PTR35) );
  MUX2_X1 U8791 ( .A(_02241__PTR4), .B(di2_PTR4), .S(_02130__PTR13), .Z(_02194__PTR36) );
  MUX2_X1 U8792 ( .A(_02241__PTR5), .B(di2_PTR5), .S(_02130__PTR13), .Z(_02194__PTR37) );
  MUX2_X1 U8793 ( .A(_02241__PTR6), .B(di2_PTR6), .S(_02130__PTR13), .Z(_02194__PTR38) );
  MUX2_X1 U8794 ( .A(_02241__PTR7), .B(di2_PTR7), .S(_02130__PTR13), .Z(_02194__PTR39) );
  MUX2_X1 U8795 ( .A(_02240__PTR0), .B(di2_PTR0), .S(_02130__PTR14), .Z(_02192__PTR32) );
  MUX2_X1 U8796 ( .A(_02240__PTR1), .B(di2_PTR1), .S(_02130__PTR14), .Z(_02192__PTR33) );
  MUX2_X1 U8797 ( .A(_02240__PTR2), .B(di2_PTR2), .S(_02130__PTR14), .Z(_02192__PTR34) );
  MUX2_X1 U8798 ( .A(_02240__PTR3), .B(di2_PTR3), .S(_02130__PTR14), .Z(_02192__PTR35) );
  MUX2_X1 U8799 ( .A(_02240__PTR4), .B(di2_PTR4), .S(_02130__PTR14), .Z(_02192__PTR36) );
  MUX2_X1 U8800 ( .A(_02240__PTR5), .B(di2_PTR5), .S(_02130__PTR14), .Z(_02192__PTR37) );
  MUX2_X1 U8801 ( .A(_02240__PTR6), .B(di2_PTR6), .S(_02130__PTR14), .Z(_02192__PTR38) );
  MUX2_X1 U8802 ( .A(_02240__PTR7), .B(di2_PTR7), .S(_02130__PTR14), .Z(_02192__PTR39) );
  MUX2_X1 U8803 ( .A(_02239__PTR0), .B(di2_PTR0), .S(_02130__PTR15), .Z(_02190__PTR32) );
  MUX2_X1 U8804 ( .A(_02239__PTR1), .B(di2_PTR1), .S(_02130__PTR15), .Z(_02190__PTR33) );
  MUX2_X1 U8805 ( .A(_02239__PTR2), .B(di2_PTR2), .S(_02130__PTR15), .Z(_02190__PTR34) );
  MUX2_X1 U8806 ( .A(_02239__PTR3), .B(di2_PTR3), .S(_02130__PTR15), .Z(_02190__PTR35) );
  MUX2_X1 U8807 ( .A(_02239__PTR4), .B(di2_PTR4), .S(_02130__PTR15), .Z(_02190__PTR36) );
  MUX2_X1 U8808 ( .A(_02239__PTR5), .B(di2_PTR5), .S(_02130__PTR15), .Z(_02190__PTR37) );
  MUX2_X1 U8809 ( .A(_02239__PTR6), .B(di2_PTR6), .S(_02130__PTR15), .Z(_02190__PTR38) );
  MUX2_X1 U8810 ( .A(_02239__PTR7), .B(di2_PTR7), .S(_02130__PTR15), .Z(_02190__PTR39) );
  MUX2_X1 U8811 ( .A(P2_P1_InstQueue_PTR0_PTR0), .B(di2_PTR0), .S(_02128__PTR0), .Z(_02254__PTR0) );
  MUX2_X1 U8812 ( .A(P2_P1_InstQueue_PTR0_PTR1), .B(di2_PTR1), .S(_02128__PTR0), .Z(_02254__PTR1) );
  MUX2_X1 U8813 ( .A(P2_P1_InstQueue_PTR0_PTR2), .B(di2_PTR2), .S(_02128__PTR0), .Z(_02254__PTR2) );
  MUX2_X1 U8814 ( .A(P2_P1_InstQueue_PTR0_PTR3), .B(di2_PTR3), .S(_02128__PTR0), .Z(_02254__PTR3) );
  MUX2_X1 U8815 ( .A(P2_P1_InstQueue_PTR0_PTR4), .B(di2_PTR4), .S(_02128__PTR0), .Z(_02254__PTR4) );
  MUX2_X1 U8816 ( .A(P2_P1_InstQueue_PTR0_PTR5), .B(di2_PTR5), .S(_02128__PTR0), .Z(_02254__PTR5) );
  MUX2_X1 U8817 ( .A(P2_P1_InstQueue_PTR0_PTR6), .B(di2_PTR6), .S(_02128__PTR0), .Z(_02254__PTR6) );
  MUX2_X1 U8818 ( .A(P2_P1_InstQueue_PTR0_PTR7), .B(di2_PTR7), .S(_02128__PTR0), .Z(_02254__PTR7) );
  MUX2_X1 U8819 ( .A(P2_P1_InstQueue_PTR1_PTR0), .B(di2_PTR0), .S(_02128__PTR1), .Z(_02253__PTR0) );
  MUX2_X1 U8820 ( .A(P2_P1_InstQueue_PTR1_PTR1), .B(di2_PTR1), .S(_02128__PTR1), .Z(_02253__PTR1) );
  MUX2_X1 U8821 ( .A(P2_P1_InstQueue_PTR1_PTR2), .B(di2_PTR2), .S(_02128__PTR1), .Z(_02253__PTR2) );
  MUX2_X1 U8822 ( .A(P2_P1_InstQueue_PTR1_PTR3), .B(di2_PTR3), .S(_02128__PTR1), .Z(_02253__PTR3) );
  MUX2_X1 U8823 ( .A(P2_P1_InstQueue_PTR1_PTR4), .B(di2_PTR4), .S(_02128__PTR1), .Z(_02253__PTR4) );
  MUX2_X1 U8824 ( .A(P2_P1_InstQueue_PTR1_PTR5), .B(di2_PTR5), .S(_02128__PTR1), .Z(_02253__PTR5) );
  MUX2_X1 U8825 ( .A(P2_P1_InstQueue_PTR1_PTR6), .B(di2_PTR6), .S(_02128__PTR1), .Z(_02253__PTR6) );
  MUX2_X1 U8826 ( .A(P2_P1_InstQueue_PTR1_PTR7), .B(di2_PTR7), .S(_02128__PTR1), .Z(_02253__PTR7) );
  MUX2_X1 U8827 ( .A(P2_P1_InstQueue_PTR2_PTR0), .B(di2_PTR0), .S(_02128__PTR2), .Z(_02252__PTR0) );
  MUX2_X1 U8828 ( .A(P2_P1_InstQueue_PTR2_PTR1), .B(di2_PTR1), .S(_02128__PTR2), .Z(_02252__PTR1) );
  MUX2_X1 U8829 ( .A(P2_P1_InstQueue_PTR2_PTR2), .B(di2_PTR2), .S(_02128__PTR2), .Z(_02252__PTR2) );
  MUX2_X1 U8830 ( .A(P2_P1_InstQueue_PTR2_PTR3), .B(di2_PTR3), .S(_02128__PTR2), .Z(_02252__PTR3) );
  MUX2_X1 U8831 ( .A(P2_P1_InstQueue_PTR2_PTR4), .B(di2_PTR4), .S(_02128__PTR2), .Z(_02252__PTR4) );
  MUX2_X1 U8832 ( .A(P2_P1_InstQueue_PTR2_PTR5), .B(di2_PTR5), .S(_02128__PTR2), .Z(_02252__PTR5) );
  MUX2_X1 U8833 ( .A(P2_P1_InstQueue_PTR2_PTR6), .B(di2_PTR6), .S(_02128__PTR2), .Z(_02252__PTR6) );
  MUX2_X1 U8834 ( .A(P2_P1_InstQueue_PTR2_PTR7), .B(di2_PTR7), .S(_02128__PTR2), .Z(_02252__PTR7) );
  MUX2_X1 U8835 ( .A(P2_P1_InstQueue_PTR3_PTR0), .B(di2_PTR0), .S(_02128__PTR3), .Z(_02251__PTR0) );
  MUX2_X1 U8836 ( .A(P2_P1_InstQueue_PTR3_PTR1), .B(di2_PTR1), .S(_02128__PTR3), .Z(_02251__PTR1) );
  MUX2_X1 U8837 ( .A(P2_P1_InstQueue_PTR3_PTR2), .B(di2_PTR2), .S(_02128__PTR3), .Z(_02251__PTR2) );
  MUX2_X1 U8838 ( .A(P2_P1_InstQueue_PTR3_PTR3), .B(di2_PTR3), .S(_02128__PTR3), .Z(_02251__PTR3) );
  MUX2_X1 U8839 ( .A(P2_P1_InstQueue_PTR3_PTR4), .B(di2_PTR4), .S(_02128__PTR3), .Z(_02251__PTR4) );
  MUX2_X1 U8840 ( .A(P2_P1_InstQueue_PTR3_PTR5), .B(di2_PTR5), .S(_02128__PTR3), .Z(_02251__PTR5) );
  MUX2_X1 U8841 ( .A(P2_P1_InstQueue_PTR3_PTR6), .B(di2_PTR6), .S(_02128__PTR3), .Z(_02251__PTR6) );
  MUX2_X1 U8842 ( .A(P2_P1_InstQueue_PTR3_PTR7), .B(di2_PTR7), .S(_02128__PTR3), .Z(_02251__PTR7) );
  MUX2_X1 U8843 ( .A(P2_P1_InstQueue_PTR4_PTR0), .B(di2_PTR0), .S(_02128__PTR4), .Z(_02250__PTR0) );
  MUX2_X1 U8844 ( .A(P2_P1_InstQueue_PTR4_PTR1), .B(di2_PTR1), .S(_02128__PTR4), .Z(_02250__PTR1) );
  MUX2_X1 U8845 ( .A(P2_P1_InstQueue_PTR4_PTR2), .B(di2_PTR2), .S(_02128__PTR4), .Z(_02250__PTR2) );
  MUX2_X1 U8846 ( .A(P2_P1_InstQueue_PTR4_PTR3), .B(di2_PTR3), .S(_02128__PTR4), .Z(_02250__PTR3) );
  MUX2_X1 U8847 ( .A(P2_P1_InstQueue_PTR4_PTR4), .B(di2_PTR4), .S(_02128__PTR4), .Z(_02250__PTR4) );
  MUX2_X1 U8848 ( .A(P2_P1_InstQueue_PTR4_PTR5), .B(di2_PTR5), .S(_02128__PTR4), .Z(_02250__PTR5) );
  MUX2_X1 U8849 ( .A(P2_P1_InstQueue_PTR4_PTR6), .B(di2_PTR6), .S(_02128__PTR4), .Z(_02250__PTR6) );
  MUX2_X1 U8850 ( .A(P2_P1_InstQueue_PTR4_PTR7), .B(di2_PTR7), .S(_02128__PTR4), .Z(_02250__PTR7) );
  MUX2_X1 U8851 ( .A(P2_P1_InstQueue_PTR5_PTR0), .B(di2_PTR0), .S(_02128__PTR5), .Z(_02249__PTR0) );
  MUX2_X1 U8852 ( .A(P2_P1_InstQueue_PTR5_PTR1), .B(di2_PTR1), .S(_02128__PTR5), .Z(_02249__PTR1) );
  MUX2_X1 U8853 ( .A(P2_P1_InstQueue_PTR5_PTR2), .B(di2_PTR2), .S(_02128__PTR5), .Z(_02249__PTR2) );
  MUX2_X1 U8854 ( .A(P2_P1_InstQueue_PTR5_PTR3), .B(di2_PTR3), .S(_02128__PTR5), .Z(_02249__PTR3) );
  MUX2_X1 U8855 ( .A(P2_P1_InstQueue_PTR5_PTR4), .B(di2_PTR4), .S(_02128__PTR5), .Z(_02249__PTR4) );
  MUX2_X1 U8856 ( .A(P2_P1_InstQueue_PTR5_PTR5), .B(di2_PTR5), .S(_02128__PTR5), .Z(_02249__PTR5) );
  MUX2_X1 U8857 ( .A(P2_P1_InstQueue_PTR5_PTR6), .B(di2_PTR6), .S(_02128__PTR5), .Z(_02249__PTR6) );
  MUX2_X1 U8858 ( .A(P2_P1_InstQueue_PTR5_PTR7), .B(di2_PTR7), .S(_02128__PTR5), .Z(_02249__PTR7) );
  MUX2_X1 U8859 ( .A(P2_P1_InstQueue_PTR6_PTR0), .B(di2_PTR0), .S(_02128__PTR6), .Z(_02248__PTR0) );
  MUX2_X1 U8860 ( .A(P2_P1_InstQueue_PTR6_PTR1), .B(di2_PTR1), .S(_02128__PTR6), .Z(_02248__PTR1) );
  MUX2_X1 U8861 ( .A(P2_P1_InstQueue_PTR6_PTR2), .B(di2_PTR2), .S(_02128__PTR6), .Z(_02248__PTR2) );
  MUX2_X1 U8862 ( .A(P2_P1_InstQueue_PTR6_PTR3), .B(di2_PTR3), .S(_02128__PTR6), .Z(_02248__PTR3) );
  MUX2_X1 U8863 ( .A(P2_P1_InstQueue_PTR6_PTR4), .B(di2_PTR4), .S(_02128__PTR6), .Z(_02248__PTR4) );
  MUX2_X1 U8864 ( .A(P2_P1_InstQueue_PTR6_PTR5), .B(di2_PTR5), .S(_02128__PTR6), .Z(_02248__PTR5) );
  MUX2_X1 U8865 ( .A(P2_P1_InstQueue_PTR6_PTR6), .B(di2_PTR6), .S(_02128__PTR6), .Z(_02248__PTR6) );
  MUX2_X1 U8866 ( .A(P2_P1_InstQueue_PTR6_PTR7), .B(di2_PTR7), .S(_02128__PTR6), .Z(_02248__PTR7) );
  MUX2_X1 U8867 ( .A(P2_P1_InstQueue_PTR7_PTR0), .B(di2_PTR0), .S(_02128__PTR7), .Z(_02247__PTR0) );
  MUX2_X1 U8868 ( .A(P2_P1_InstQueue_PTR7_PTR1), .B(di2_PTR1), .S(_02128__PTR7), .Z(_02247__PTR1) );
  MUX2_X1 U8869 ( .A(P2_P1_InstQueue_PTR7_PTR2), .B(di2_PTR2), .S(_02128__PTR7), .Z(_02247__PTR2) );
  MUX2_X1 U8870 ( .A(P2_P1_InstQueue_PTR7_PTR3), .B(di2_PTR3), .S(_02128__PTR7), .Z(_02247__PTR3) );
  MUX2_X1 U8871 ( .A(P2_P1_InstQueue_PTR7_PTR4), .B(di2_PTR4), .S(_02128__PTR7), .Z(_02247__PTR4) );
  MUX2_X1 U8872 ( .A(P2_P1_InstQueue_PTR7_PTR5), .B(di2_PTR5), .S(_02128__PTR7), .Z(_02247__PTR5) );
  MUX2_X1 U8873 ( .A(P2_P1_InstQueue_PTR7_PTR6), .B(di2_PTR6), .S(_02128__PTR7), .Z(_02247__PTR6) );
  MUX2_X1 U8874 ( .A(P2_P1_InstQueue_PTR7_PTR7), .B(di2_PTR7), .S(_02128__PTR7), .Z(_02247__PTR7) );
  MUX2_X1 U8875 ( .A(P2_P1_InstQueue_PTR8_PTR0), .B(di2_PTR0), .S(_02128__PTR8), .Z(_02246__PTR0) );
  MUX2_X1 U8876 ( .A(P2_P1_InstQueue_PTR8_PTR1), .B(di2_PTR1), .S(_02128__PTR8), .Z(_02246__PTR1) );
  MUX2_X1 U8877 ( .A(P2_P1_InstQueue_PTR8_PTR2), .B(di2_PTR2), .S(_02128__PTR8), .Z(_02246__PTR2) );
  MUX2_X1 U8878 ( .A(P2_P1_InstQueue_PTR8_PTR3), .B(di2_PTR3), .S(_02128__PTR8), .Z(_02246__PTR3) );
  MUX2_X1 U8879 ( .A(P2_P1_InstQueue_PTR8_PTR4), .B(di2_PTR4), .S(_02128__PTR8), .Z(_02246__PTR4) );
  MUX2_X1 U8880 ( .A(P2_P1_InstQueue_PTR8_PTR5), .B(di2_PTR5), .S(_02128__PTR8), .Z(_02246__PTR5) );
  MUX2_X1 U8881 ( .A(P2_P1_InstQueue_PTR8_PTR6), .B(di2_PTR6), .S(_02128__PTR8), .Z(_02246__PTR6) );
  MUX2_X1 U8882 ( .A(P2_P1_InstQueue_PTR8_PTR7), .B(di2_PTR7), .S(_02128__PTR8), .Z(_02246__PTR7) );
  MUX2_X1 U8883 ( .A(P2_P1_InstQueue_PTR9_PTR0), .B(di2_PTR0), .S(_02128__PTR9), .Z(_02245__PTR0) );
  MUX2_X1 U8884 ( .A(P2_P1_InstQueue_PTR9_PTR1), .B(di2_PTR1), .S(_02128__PTR9), .Z(_02245__PTR1) );
  MUX2_X1 U8885 ( .A(P2_P1_InstQueue_PTR9_PTR2), .B(di2_PTR2), .S(_02128__PTR9), .Z(_02245__PTR2) );
  MUX2_X1 U8886 ( .A(P2_P1_InstQueue_PTR9_PTR3), .B(di2_PTR3), .S(_02128__PTR9), .Z(_02245__PTR3) );
  MUX2_X1 U8887 ( .A(P2_P1_InstQueue_PTR9_PTR4), .B(di2_PTR4), .S(_02128__PTR9), .Z(_02245__PTR4) );
  MUX2_X1 U8888 ( .A(P2_P1_InstQueue_PTR9_PTR5), .B(di2_PTR5), .S(_02128__PTR9), .Z(_02245__PTR5) );
  MUX2_X1 U8889 ( .A(P2_P1_InstQueue_PTR9_PTR6), .B(di2_PTR6), .S(_02128__PTR9), .Z(_02245__PTR6) );
  MUX2_X1 U8890 ( .A(P2_P1_InstQueue_PTR9_PTR7), .B(di2_PTR7), .S(_02128__PTR9), .Z(_02245__PTR7) );
  MUX2_X1 U8891 ( .A(P2_P1_InstQueue_PTR10_PTR0), .B(di2_PTR0), .S(_02128__PTR10), .Z(_02244__PTR0) );
  MUX2_X1 U8892 ( .A(P2_P1_InstQueue_PTR10_PTR1), .B(di2_PTR1), .S(_02128__PTR10), .Z(_02244__PTR1) );
  MUX2_X1 U8893 ( .A(P2_P1_InstQueue_PTR10_PTR2), .B(di2_PTR2), .S(_02128__PTR10), .Z(_02244__PTR2) );
  MUX2_X1 U8894 ( .A(P2_P1_InstQueue_PTR10_PTR3), .B(di2_PTR3), .S(_02128__PTR10), .Z(_02244__PTR3) );
  MUX2_X1 U8895 ( .A(P2_P1_InstQueue_PTR10_PTR4), .B(di2_PTR4), .S(_02128__PTR10), .Z(_02244__PTR4) );
  MUX2_X1 U8896 ( .A(P2_P1_InstQueue_PTR10_PTR5), .B(di2_PTR5), .S(_02128__PTR10), .Z(_02244__PTR5) );
  MUX2_X1 U8897 ( .A(P2_P1_InstQueue_PTR10_PTR6), .B(di2_PTR6), .S(_02128__PTR10), .Z(_02244__PTR6) );
  MUX2_X1 U8898 ( .A(P2_P1_InstQueue_PTR10_PTR7), .B(di2_PTR7), .S(_02128__PTR10), .Z(_02244__PTR7) );
  MUX2_X1 U8899 ( .A(P2_P1_InstQueue_PTR11_PTR0), .B(di2_PTR0), .S(_02128__PTR11), .Z(_02243__PTR0) );
  MUX2_X1 U8900 ( .A(P2_P1_InstQueue_PTR11_PTR1), .B(di2_PTR1), .S(_02128__PTR11), .Z(_02243__PTR1) );
  MUX2_X1 U8901 ( .A(P2_P1_InstQueue_PTR11_PTR2), .B(di2_PTR2), .S(_02128__PTR11), .Z(_02243__PTR2) );
  MUX2_X1 U8902 ( .A(P2_P1_InstQueue_PTR11_PTR3), .B(di2_PTR3), .S(_02128__PTR11), .Z(_02243__PTR3) );
  MUX2_X1 U8903 ( .A(P2_P1_InstQueue_PTR11_PTR4), .B(di2_PTR4), .S(_02128__PTR11), .Z(_02243__PTR4) );
  MUX2_X1 U8904 ( .A(P2_P1_InstQueue_PTR11_PTR5), .B(di2_PTR5), .S(_02128__PTR11), .Z(_02243__PTR5) );
  MUX2_X1 U8905 ( .A(P2_P1_InstQueue_PTR11_PTR6), .B(di2_PTR6), .S(_02128__PTR11), .Z(_02243__PTR6) );
  MUX2_X1 U8906 ( .A(P2_P1_InstQueue_PTR11_PTR7), .B(di2_PTR7), .S(_02128__PTR11), .Z(_02243__PTR7) );
  MUX2_X1 U8907 ( .A(P2_P1_InstQueue_PTR12_PTR0), .B(di2_PTR0), .S(_02128__PTR12), .Z(_02242__PTR0) );
  MUX2_X1 U8908 ( .A(P2_P1_InstQueue_PTR12_PTR1), .B(di2_PTR1), .S(_02128__PTR12), .Z(_02242__PTR1) );
  MUX2_X1 U8909 ( .A(P2_P1_InstQueue_PTR12_PTR2), .B(di2_PTR2), .S(_02128__PTR12), .Z(_02242__PTR2) );
  MUX2_X1 U8910 ( .A(P2_P1_InstQueue_PTR12_PTR3), .B(di2_PTR3), .S(_02128__PTR12), .Z(_02242__PTR3) );
  MUX2_X1 U8911 ( .A(P2_P1_InstQueue_PTR12_PTR4), .B(di2_PTR4), .S(_02128__PTR12), .Z(_02242__PTR4) );
  MUX2_X1 U8912 ( .A(P2_P1_InstQueue_PTR12_PTR5), .B(di2_PTR5), .S(_02128__PTR12), .Z(_02242__PTR5) );
  MUX2_X1 U8913 ( .A(P2_P1_InstQueue_PTR12_PTR6), .B(di2_PTR6), .S(_02128__PTR12), .Z(_02242__PTR6) );
  MUX2_X1 U8914 ( .A(P2_P1_InstQueue_PTR12_PTR7), .B(di2_PTR7), .S(_02128__PTR12), .Z(_02242__PTR7) );
  MUX2_X1 U8915 ( .A(P2_P1_InstQueue_PTR13_PTR0), .B(di2_PTR0), .S(_02128__PTR13), .Z(_02241__PTR0) );
  MUX2_X1 U8916 ( .A(P2_P1_InstQueue_PTR13_PTR1), .B(di2_PTR1), .S(_02128__PTR13), .Z(_02241__PTR1) );
  MUX2_X1 U8917 ( .A(P2_P1_InstQueue_PTR13_PTR2), .B(di2_PTR2), .S(_02128__PTR13), .Z(_02241__PTR2) );
  MUX2_X1 U8918 ( .A(P2_P1_InstQueue_PTR13_PTR3), .B(di2_PTR3), .S(_02128__PTR13), .Z(_02241__PTR3) );
  MUX2_X1 U8919 ( .A(P2_P1_InstQueue_PTR13_PTR4), .B(di2_PTR4), .S(_02128__PTR13), .Z(_02241__PTR4) );
  MUX2_X1 U8920 ( .A(P2_P1_InstQueue_PTR13_PTR5), .B(di2_PTR5), .S(_02128__PTR13), .Z(_02241__PTR5) );
  MUX2_X1 U8921 ( .A(P2_P1_InstQueue_PTR13_PTR6), .B(di2_PTR6), .S(_02128__PTR13), .Z(_02241__PTR6) );
  MUX2_X1 U8922 ( .A(P2_P1_InstQueue_PTR13_PTR7), .B(di2_PTR7), .S(_02128__PTR13), .Z(_02241__PTR7) );
  MUX2_X1 U8923 ( .A(P2_P1_InstQueue_PTR14_PTR0), .B(di2_PTR0), .S(_02128__PTR14), .Z(_02240__PTR0) );
  MUX2_X1 U8924 ( .A(P2_P1_InstQueue_PTR14_PTR1), .B(di2_PTR1), .S(_02128__PTR14), .Z(_02240__PTR1) );
  MUX2_X1 U8925 ( .A(P2_P1_InstQueue_PTR14_PTR2), .B(di2_PTR2), .S(_02128__PTR14), .Z(_02240__PTR2) );
  MUX2_X1 U8926 ( .A(P2_P1_InstQueue_PTR14_PTR3), .B(di2_PTR3), .S(_02128__PTR14), .Z(_02240__PTR3) );
  MUX2_X1 U8927 ( .A(P2_P1_InstQueue_PTR14_PTR4), .B(di2_PTR4), .S(_02128__PTR14), .Z(_02240__PTR4) );
  MUX2_X1 U8928 ( .A(P2_P1_InstQueue_PTR14_PTR5), .B(di2_PTR5), .S(_02128__PTR14), .Z(_02240__PTR5) );
  MUX2_X1 U8929 ( .A(P2_P1_InstQueue_PTR14_PTR6), .B(di2_PTR6), .S(_02128__PTR14), .Z(_02240__PTR6) );
  MUX2_X1 U8930 ( .A(P2_P1_InstQueue_PTR14_PTR7), .B(di2_PTR7), .S(_02128__PTR14), .Z(_02240__PTR7) );
  MUX2_X1 U8931 ( .A(P2_P1_InstQueue_PTR15_PTR0), .B(di2_PTR0), .S(_02128__PTR15), .Z(_02239__PTR0) );
  MUX2_X1 U8932 ( .A(P2_P1_InstQueue_PTR15_PTR1), .B(di2_PTR1), .S(_02128__PTR15), .Z(_02239__PTR1) );
  MUX2_X1 U8933 ( .A(P2_P1_InstQueue_PTR15_PTR2), .B(di2_PTR2), .S(_02128__PTR15), .Z(_02239__PTR2) );
  MUX2_X1 U8934 ( .A(P2_P1_InstQueue_PTR15_PTR3), .B(di2_PTR3), .S(_02128__PTR15), .Z(_02239__PTR3) );
  MUX2_X1 U8935 ( .A(P2_P1_InstQueue_PTR15_PTR4), .B(di2_PTR4), .S(_02128__PTR15), .Z(_02239__PTR4) );
  MUX2_X1 U8936 ( .A(P2_P1_InstQueue_PTR15_PTR5), .B(di2_PTR5), .S(_02128__PTR15), .Z(_02239__PTR5) );
  MUX2_X1 U8937 ( .A(P2_P1_InstQueue_PTR15_PTR6), .B(di2_PTR6), .S(_02128__PTR15), .Z(_02239__PTR6) );
  MUX2_X1 U8938 ( .A(P2_P1_InstQueue_PTR15_PTR7), .B(di2_PTR7), .S(_02128__PTR15), .Z(_02239__PTR7) );
  MUX2_X1 U8939 ( .A(_02238__PTR0), .B(1'b0), .S(_02233_), .Z(_02169__PTR28) );
  MUX2_X1 U8940 ( .A(_02238__PTR1), .B(1'b1), .S(_02233_), .Z(_02169__PTR29) );
  MUX2_X1 U8941 ( .A(_02238__PTR2), .B(1'b1), .S(_02233_), .Z(_02169__PTR30) );
  MUX2_X1 U8942 ( .A(_02237__PTR0), .B(1'b1), .S(_02234_), .Z(_02238__PTR0) );
  MUX2_X1 U8943 ( .A(_02237__PTR1), .B(1'b0), .S(_02234_), .Z(_02238__PTR1) );
  MUX2_X1 U8944 ( .A(_02237__PTR2), .B(1'b1), .S(_02234_), .Z(_02238__PTR2) );
  INV_X1 U8945 ( .A(_01767__PTR4), .ZN(_02237__PTR0) );
  MUX2_X1 U8946 ( .A(_02236__PTR2), .B(1'b1), .S(_01767__PTR4), .Z(_02237__PTR1) );
  MUX2_X1 U8947 ( .A(_02236__PTR2), .B(1'b0), .S(_01767__PTR4), .Z(_02237__PTR2) );
  INV_X1 U8948 ( .A(_02235_), .ZN(_02236__PTR2) );
  MUX2_X1 U8949 ( .A(P2_EAX_PTR16), .B(_02334__PTR16), .S(_02296_), .Z(_02385__PTR80) );
  MUX2_X1 U8950 ( .A(P2_EAX_PTR17), .B(_02334__PTR17), .S(_02296_), .Z(_02385__PTR81) );
  MUX2_X1 U8951 ( .A(P2_EAX_PTR18), .B(_02334__PTR18), .S(_02296_), .Z(_02385__PTR82) );
  MUX2_X1 U8952 ( .A(P2_EAX_PTR19), .B(_02334__PTR19), .S(_02296_), .Z(_02385__PTR83) );
  MUX2_X1 U8953 ( .A(P2_EAX_PTR20), .B(_02334__PTR20), .S(_02296_), .Z(_02385__PTR84) );
  MUX2_X1 U8954 ( .A(P2_EAX_PTR21), .B(_02334__PTR21), .S(_02296_), .Z(_02385__PTR85) );
  MUX2_X1 U8955 ( .A(P2_EAX_PTR22), .B(_02334__PTR22), .S(_02296_), .Z(_02385__PTR86) );
  MUX2_X1 U8956 ( .A(P2_EAX_PTR23), .B(_02334__PTR23), .S(_02296_), .Z(_02385__PTR87) );
  MUX2_X1 U8957 ( .A(P2_EAX_PTR24), .B(_02334__PTR24), .S(_02296_), .Z(_02385__PTR88) );
  MUX2_X1 U8958 ( .A(P2_EAX_PTR25), .B(_02334__PTR25), .S(_02296_), .Z(_02385__PTR89) );
  MUX2_X1 U8959 ( .A(P2_EAX_PTR26), .B(_02334__PTR26), .S(_02296_), .Z(_02385__PTR90) );
  MUX2_X1 U8960 ( .A(P2_EAX_PTR27), .B(_02334__PTR27), .S(_02296_), .Z(_02385__PTR91) );
  MUX2_X1 U8961 ( .A(P2_EAX_PTR28), .B(_02334__PTR28), .S(_02296_), .Z(_02385__PTR92) );
  MUX2_X1 U8962 ( .A(P2_EAX_PTR29), .B(_02334__PTR29), .S(_02296_), .Z(_02385__PTR93) );
  MUX2_X1 U8963 ( .A(P2_EAX_PTR30), .B(_02334__PTR30), .S(_02296_), .Z(_02385__PTR94) );
  MUX2_X1 U8964 ( .A(P2_EAX_PTR31), .B(_02334__PTR31), .S(_02296_), .Z(_02385__PTR95) );
  MUX2_X1 U8965 ( .A(P2_EAX_PTR0), .B(_02306__PTR0), .S(_02296_), .Z(_02385__PTR96) );
  MUX2_X1 U8966 ( .A(P2_EAX_PTR1), .B(_02306__PTR1), .S(_02296_), .Z(_02385__PTR97) );
  MUX2_X1 U8967 ( .A(P2_EAX_PTR2), .B(_02306__PTR2), .S(_02296_), .Z(_02385__PTR98) );
  MUX2_X1 U8968 ( .A(P2_EAX_PTR3), .B(_02306__PTR3), .S(_02296_), .Z(_02385__PTR99) );
  MUX2_X1 U8969 ( .A(P2_EAX_PTR4), .B(_02306__PTR4), .S(_02296_), .Z(_02385__PTR100) );
  MUX2_X1 U8970 ( .A(P2_EAX_PTR5), .B(_02306__PTR5), .S(_02296_), .Z(_02385__PTR101) );
  MUX2_X1 U8971 ( .A(P2_EAX_PTR6), .B(_02306__PTR6), .S(_02296_), .Z(_02385__PTR102) );
  MUX2_X1 U8972 ( .A(P2_EAX_PTR7), .B(_02306__PTR7), .S(_02296_), .Z(_02385__PTR103) );
  MUX2_X1 U8973 ( .A(P2_EAX_PTR8), .B(_02306__PTR8), .S(_02296_), .Z(_02385__PTR104) );
  MUX2_X1 U8974 ( .A(P2_EAX_PTR9), .B(_02306__PTR9), .S(_02296_), .Z(_02385__PTR105) );
  MUX2_X1 U8975 ( .A(P2_EAX_PTR10), .B(_02306__PTR10), .S(_02296_), .Z(_02385__PTR106) );
  MUX2_X1 U8976 ( .A(P2_EAX_PTR11), .B(_02306__PTR11), .S(_02296_), .Z(_02385__PTR107) );
  MUX2_X1 U8977 ( .A(P2_EAX_PTR12), .B(_02306__PTR12), .S(_02296_), .Z(_02385__PTR108) );
  MUX2_X1 U8978 ( .A(P2_EAX_PTR13), .B(_02306__PTR13), .S(_02296_), .Z(_02385__PTR109) );
  MUX2_X1 U8979 ( .A(P2_EAX_PTR14), .B(_02306__PTR14), .S(_02296_), .Z(_02385__PTR110) );
  MUX2_X1 U8980 ( .A(P2_EAX_PTR15), .B(_02306__PTR15), .S(_02296_), .Z(_02385__PTR111) );
  MUX2_X1 U8981 ( .A(P2_EAX_PTR16), .B(_02306__PTR16), .S(_02296_), .Z(_02385__PTR112) );
  MUX2_X1 U8982 ( .A(P2_EAX_PTR17), .B(_02306__PTR17), .S(_02296_), .Z(_02385__PTR113) );
  MUX2_X1 U8983 ( .A(P2_EAX_PTR18), .B(_02306__PTR18), .S(_02296_), .Z(_02385__PTR114) );
  MUX2_X1 U8984 ( .A(P2_EAX_PTR19), .B(_02306__PTR19), .S(_02296_), .Z(_02385__PTR115) );
  MUX2_X1 U8985 ( .A(P2_EAX_PTR20), .B(_02306__PTR20), .S(_02296_), .Z(_02385__PTR116) );
  MUX2_X1 U8986 ( .A(P2_EAX_PTR21), .B(_02306__PTR21), .S(_02296_), .Z(_02385__PTR117) );
  MUX2_X1 U8987 ( .A(P2_EAX_PTR22), .B(_02306__PTR22), .S(_02296_), .Z(_02385__PTR118) );
  MUX2_X1 U8988 ( .A(P2_EAX_PTR23), .B(_02306__PTR23), .S(_02296_), .Z(_02385__PTR119) );
  MUX2_X1 U8989 ( .A(P2_EAX_PTR24), .B(_02306__PTR24), .S(_02296_), .Z(_02385__PTR120) );
  MUX2_X1 U8990 ( .A(P2_EAX_PTR25), .B(_02306__PTR25), .S(_02296_), .Z(_02385__PTR121) );
  MUX2_X1 U8991 ( .A(P2_EAX_PTR26), .B(_02306__PTR26), .S(_02296_), .Z(_02385__PTR122) );
  MUX2_X1 U8992 ( .A(P2_EAX_PTR27), .B(_02306__PTR27), .S(_02296_), .Z(_02385__PTR123) );
  MUX2_X1 U8993 ( .A(P2_EAX_PTR28), .B(_02306__PTR28), .S(_02296_), .Z(_02385__PTR124) );
  MUX2_X1 U8994 ( .A(P2_EAX_PTR29), .B(_02306__PTR29), .S(_02296_), .Z(_02385__PTR125) );
  MUX2_X1 U8995 ( .A(P2_EAX_PTR30), .B(_02306__PTR30), .S(_02296_), .Z(_02385__PTR126) );
  MUX2_X1 U8996 ( .A(P2_EAX_PTR31), .B(_02306__PTR31), .S(_02296_), .Z(_02385__PTR127) );
  INV_X1 U8997 ( .A(_02169__PTR21), .ZN(_02169__PTR20) );
  MUX2_X1 U8998 ( .A(_02231__PTR2), .B(1'b0), .S(_02169__PTR21), .Z(_02169__PTR22) );
  INV_X1 U8999 ( .A(_02301_), .ZN(_02231__PTR2) );
  INV_X1 U9000 ( .A(bs16), .ZN(_01878__PTR256) );
  MUX2_X1 U9001 ( .A(_02372__PTR1), .B(1'b0), .S(_02338_), .Z(_02169__PTR16) );
  MUX2_X1 U9002 ( .A(_02372__PTR1), .B(1'b1), .S(_02338_), .Z(_02169__PTR17) );
  MUX2_X1 U9003 ( .A(_02372__PTR2), .B(1'b1), .S(_02338_), .Z(_02169__PTR18) );
  MUX2_X1 U9004 ( .A(na), .B(1'b1), .S(_02349_), .Z(_02372__PTR1) );
  MUX2_X1 U9005 ( .A(_02003_), .B(1'b1), .S(_02349_), .Z(_02372__PTR2) );
  MUX2_X1 U9006 ( .A(_02333__PTR0), .B(1'b0), .S(_01767__PTR4), .Z(_02169__PTR12) );
  MUX2_X1 U9007 ( .A(_02333__PTR1), .B(1'b1), .S(_01767__PTR4), .Z(_02169__PTR13) );
  MUX2_X1 U9008 ( .A(_02333__PTR2), .B(1'b0), .S(_01767__PTR4), .Z(_02169__PTR14) );
  MUX2_X1 U9009 ( .A(_02332__PTR0), .B(1'b0), .S(_02292_), .Z(_02333__PTR0) );
  MUX2_X1 U9010 ( .A(_02332__PTR1), .B(1'b0), .S(_02292_), .Z(_02333__PTR1) );
  MUX2_X1 U9011 ( .A(_02332__PTR2), .B(1'b0), .S(_02292_), .Z(_02333__PTR2) );
  MUX2_X1 U9012 ( .A(_02331__PTR0), .B(1'b1), .S(_02295_), .Z(_02332__PTR0) );
  MUX2_X1 U9013 ( .A(_02331__PTR1), .B(1'b1), .S(_02295_), .Z(_02332__PTR1) );
  MUX2_X1 U9014 ( .A(_02331__PTR2), .B(1'b1), .S(_02295_), .Z(_02332__PTR2) );
  INV_X1 U9015 ( .A(_02298_), .ZN(_02331__PTR0) );
  MUX2_X1 U9016 ( .A(_02330__PTR1), .B(1'b1), .S(_02298_), .Z(_02331__PTR1) );
  MUX2_X1 U9017 ( .A(_02330__PTR2), .B(1'b1), .S(_02298_), .Z(_02331__PTR2) );
  MUX2_X1 U9018 ( .A(_02329__PTR1), .B(1'b0), .S(_02302_), .Z(_02330__PTR1) );
  MUX2_X1 U9019 ( .A(_02311_), .B(1'b0), .S(_02302_), .Z(_02330__PTR2) );
  INV_X1 U9020 ( .A(_02311_), .ZN(_02329__PTR1) );
  INV_X1 U9021 ( .A(P2_CodeFetch), .ZN(_02135__PTR6) );
  INV_X1 U9022 ( .A(P2_ReadRequest), .ZN(_02139__PTR6) );
  INV_X1 U9023 ( .A(P2_RequestPending), .ZN(_02169__PTR4) );
  MUX2_X1 U9024 ( .A(hold), .B(1'b0), .S(P2_RequestPending), .Z(_02169__PTR6) );
  MUX2_X1 U9025 ( .A(1'b0), .B(_02418__PTR0), .S(_01766__PTR2), .Z(_02511__PTR64) );
  MUX2_X1 U9026 ( .A(1'b0), .B(_02418__PTR1), .S(_01766__PTR2), .Z(_02511__PTR65) );
  MUX2_X1 U9027 ( .A(1'b0), .B(_02418__PTR2), .S(_01766__PTR2), .Z(_02511__PTR66) );
  MUX2_X1 U9028 ( .A(1'b0), .B(_02418__PTR3), .S(_01766__PTR2), .Z(_02511__PTR67) );
  MUX2_X1 U9029 ( .A(1'b0), .B(1'b0), .S(_01766__PTR2), .Z(_02511__PTR68) );
  MUX2_X1 U9030 ( .A(1'b0), .B(_02465__PTR3), .S(_01766__PTR2), .Z(_02513__PTR64) );
  MUX2_X1 U9031 ( .A(1'b0), .B(_02465__PTR4), .S(_01766__PTR2), .Z(_02513__PTR65) );
  MUX2_X1 U9032 ( .A(1'b0), .B(_02465__PTR5), .S(_01766__PTR2), .Z(_02513__PTR66) );
  MUX2_X1 U9033 ( .A(1'b0), .B(_02465__PTR6), .S(_01766__PTR2), .Z(_02513__PTR67) );
  MUX2_X1 U9034 ( .A(1'b0), .B(_02660__PTR0), .S(_01766__PTR2), .Z(_02509__PTR64) );
  MUX2_X1 U9035 ( .A(1'b0), .B(_02660__PTR1), .S(_01766__PTR2), .Z(_02509__PTR65) );
  MUX2_X1 U9036 ( .A(1'b0), .B(_02660__PTR2), .S(_01766__PTR2), .Z(_02509__PTR66) );
  MUX2_X1 U9037 ( .A(1'b0), .B(_02660__PTR3), .S(_01766__PTR2), .Z(_02509__PTR67) );
  MUX2_X1 U9038 ( .A(1'b0), .B(_02660__PTR4), .S(_01766__PTR2), .Z(_02509__PTR68) );
  MUX2_X1 U9039 ( .A(1'b0), .B(_02660__PTR5), .S(_01766__PTR2), .Z(_02509__PTR69) );
  MUX2_X1 U9040 ( .A(1'b0), .B(_02660__PTR6), .S(_01766__PTR2), .Z(_02509__PTR70) );
  MUX2_X1 U9041 ( .A(1'b0), .B(_02660__PTR7), .S(_01766__PTR2), .Z(_02509__PTR71) );
  MUX2_X1 U9042 ( .A(1'b0), .B(_02659__PTR0), .S(_01766__PTR2), .Z(_02507__PTR64) );
  MUX2_X1 U9043 ( .A(1'b0), .B(_02659__PTR1), .S(_01766__PTR2), .Z(_02507__PTR65) );
  MUX2_X1 U9044 ( .A(1'b0), .B(_02659__PTR2), .S(_01766__PTR2), .Z(_02507__PTR66) );
  MUX2_X1 U9045 ( .A(1'b0), .B(_02659__PTR3), .S(_01766__PTR2), .Z(_02507__PTR67) );
  MUX2_X1 U9046 ( .A(1'b0), .B(_02659__PTR4), .S(_01766__PTR2), .Z(_02507__PTR68) );
  MUX2_X1 U9047 ( .A(1'b0), .B(_02659__PTR5), .S(_01766__PTR2), .Z(_02507__PTR69) );
  MUX2_X1 U9048 ( .A(1'b0), .B(_02659__PTR6), .S(_01766__PTR2), .Z(_02507__PTR70) );
  MUX2_X1 U9049 ( .A(1'b0), .B(_02659__PTR7), .S(_01766__PTR2), .Z(_02507__PTR71) );
  MUX2_X1 U9050 ( .A(1'b0), .B(_02658__PTR0), .S(_01766__PTR2), .Z(_02505__PTR64) );
  MUX2_X1 U9051 ( .A(1'b0), .B(_02658__PTR1), .S(_01766__PTR2), .Z(_02505__PTR65) );
  MUX2_X1 U9052 ( .A(1'b0), .B(_02658__PTR2), .S(_01766__PTR2), .Z(_02505__PTR66) );
  MUX2_X1 U9053 ( .A(1'b0), .B(_02658__PTR3), .S(_01766__PTR2), .Z(_02505__PTR67) );
  MUX2_X1 U9054 ( .A(1'b0), .B(_02658__PTR4), .S(_01766__PTR2), .Z(_02505__PTR68) );
  MUX2_X1 U9055 ( .A(1'b0), .B(_02658__PTR5), .S(_01766__PTR2), .Z(_02505__PTR69) );
  MUX2_X1 U9056 ( .A(1'b0), .B(_02658__PTR6), .S(_01766__PTR2), .Z(_02505__PTR70) );
  MUX2_X1 U9057 ( .A(1'b0), .B(_02658__PTR7), .S(_01766__PTR2), .Z(_02505__PTR71) );
  MUX2_X1 U9058 ( .A(1'b0), .B(_02657__PTR0), .S(_01766__PTR2), .Z(_02503__PTR64) );
  MUX2_X1 U9059 ( .A(1'b0), .B(_02657__PTR1), .S(_01766__PTR2), .Z(_02503__PTR65) );
  MUX2_X1 U9060 ( .A(1'b0), .B(_02657__PTR2), .S(_01766__PTR2), .Z(_02503__PTR66) );
  MUX2_X1 U9061 ( .A(1'b0), .B(_02657__PTR3), .S(_01766__PTR2), .Z(_02503__PTR67) );
  MUX2_X1 U9062 ( .A(1'b0), .B(_02657__PTR4), .S(_01766__PTR2), .Z(_02503__PTR68) );
  MUX2_X1 U9063 ( .A(1'b0), .B(_02657__PTR5), .S(_01766__PTR2), .Z(_02503__PTR69) );
  MUX2_X1 U9064 ( .A(1'b0), .B(_02657__PTR6), .S(_01766__PTR2), .Z(_02503__PTR70) );
  MUX2_X1 U9065 ( .A(1'b0), .B(_02657__PTR7), .S(_01766__PTR2), .Z(_02503__PTR71) );
  MUX2_X1 U9066 ( .A(1'b0), .B(_02656__PTR0), .S(_01766__PTR2), .Z(_02501__PTR64) );
  MUX2_X1 U9067 ( .A(1'b0), .B(_02656__PTR1), .S(_01766__PTR2), .Z(_02501__PTR65) );
  MUX2_X1 U9068 ( .A(1'b0), .B(_02656__PTR2), .S(_01766__PTR2), .Z(_02501__PTR66) );
  MUX2_X1 U9069 ( .A(1'b0), .B(_02656__PTR3), .S(_01766__PTR2), .Z(_02501__PTR67) );
  MUX2_X1 U9070 ( .A(1'b0), .B(_02656__PTR4), .S(_01766__PTR2), .Z(_02501__PTR68) );
  MUX2_X1 U9071 ( .A(1'b0), .B(_02656__PTR5), .S(_01766__PTR2), .Z(_02501__PTR69) );
  MUX2_X1 U9072 ( .A(1'b0), .B(_02656__PTR6), .S(_01766__PTR2), .Z(_02501__PTR70) );
  MUX2_X1 U9073 ( .A(1'b0), .B(_02656__PTR7), .S(_01766__PTR2), .Z(_02501__PTR71) );
  MUX2_X1 U9074 ( .A(1'b0), .B(_02655__PTR0), .S(_01766__PTR2), .Z(_02499__PTR64) );
  MUX2_X1 U9075 ( .A(1'b0), .B(_02655__PTR1), .S(_01766__PTR2), .Z(_02499__PTR65) );
  MUX2_X1 U9076 ( .A(1'b0), .B(_02655__PTR2), .S(_01766__PTR2), .Z(_02499__PTR66) );
  MUX2_X1 U9077 ( .A(1'b0), .B(_02655__PTR3), .S(_01766__PTR2), .Z(_02499__PTR67) );
  MUX2_X1 U9078 ( .A(1'b0), .B(_02655__PTR4), .S(_01766__PTR2), .Z(_02499__PTR68) );
  MUX2_X1 U9079 ( .A(1'b0), .B(_02655__PTR5), .S(_01766__PTR2), .Z(_02499__PTR69) );
  MUX2_X1 U9080 ( .A(1'b0), .B(_02655__PTR6), .S(_01766__PTR2), .Z(_02499__PTR70) );
  MUX2_X1 U9081 ( .A(1'b0), .B(_02655__PTR7), .S(_01766__PTR2), .Z(_02499__PTR71) );
  MUX2_X1 U9082 ( .A(1'b0), .B(_02654__PTR0), .S(_01766__PTR2), .Z(_02497__PTR64) );
  MUX2_X1 U9083 ( .A(1'b0), .B(_02654__PTR1), .S(_01766__PTR2), .Z(_02497__PTR65) );
  MUX2_X1 U9084 ( .A(1'b0), .B(_02654__PTR2), .S(_01766__PTR2), .Z(_02497__PTR66) );
  MUX2_X1 U9085 ( .A(1'b0), .B(_02654__PTR3), .S(_01766__PTR2), .Z(_02497__PTR67) );
  MUX2_X1 U9086 ( .A(1'b0), .B(_02654__PTR4), .S(_01766__PTR2), .Z(_02497__PTR68) );
  MUX2_X1 U9087 ( .A(1'b0), .B(_02654__PTR5), .S(_01766__PTR2), .Z(_02497__PTR69) );
  MUX2_X1 U9088 ( .A(1'b0), .B(_02654__PTR6), .S(_01766__PTR2), .Z(_02497__PTR70) );
  MUX2_X1 U9089 ( .A(1'b0), .B(_02654__PTR7), .S(_01766__PTR2), .Z(_02497__PTR71) );
  MUX2_X1 U9090 ( .A(1'b0), .B(_02653__PTR0), .S(_01766__PTR2), .Z(_02495__PTR64) );
  MUX2_X1 U9091 ( .A(1'b0), .B(_02653__PTR1), .S(_01766__PTR2), .Z(_02495__PTR65) );
  MUX2_X1 U9092 ( .A(1'b0), .B(_02653__PTR2), .S(_01766__PTR2), .Z(_02495__PTR66) );
  MUX2_X1 U9093 ( .A(1'b0), .B(_02653__PTR3), .S(_01766__PTR2), .Z(_02495__PTR67) );
  MUX2_X1 U9094 ( .A(1'b0), .B(_02653__PTR4), .S(_01766__PTR2), .Z(_02495__PTR68) );
  MUX2_X1 U9095 ( .A(1'b0), .B(_02653__PTR5), .S(_01766__PTR2), .Z(_02495__PTR69) );
  MUX2_X1 U9096 ( .A(1'b0), .B(_02653__PTR6), .S(_01766__PTR2), .Z(_02495__PTR70) );
  MUX2_X1 U9097 ( .A(1'b0), .B(_02653__PTR7), .S(_01766__PTR2), .Z(_02495__PTR71) );
  MUX2_X1 U9098 ( .A(1'b0), .B(_02652__PTR0), .S(_01766__PTR2), .Z(_02493__PTR64) );
  MUX2_X1 U9099 ( .A(1'b0), .B(_02652__PTR1), .S(_01766__PTR2), .Z(_02493__PTR65) );
  MUX2_X1 U9100 ( .A(1'b0), .B(_02652__PTR2), .S(_01766__PTR2), .Z(_02493__PTR66) );
  MUX2_X1 U9101 ( .A(1'b0), .B(_02652__PTR3), .S(_01766__PTR2), .Z(_02493__PTR67) );
  MUX2_X1 U9102 ( .A(1'b0), .B(_02652__PTR4), .S(_01766__PTR2), .Z(_02493__PTR68) );
  MUX2_X1 U9103 ( .A(1'b0), .B(_02652__PTR5), .S(_01766__PTR2), .Z(_02493__PTR69) );
  MUX2_X1 U9104 ( .A(1'b0), .B(_02652__PTR6), .S(_01766__PTR2), .Z(_02493__PTR70) );
  MUX2_X1 U9105 ( .A(1'b0), .B(_02652__PTR7), .S(_01766__PTR2), .Z(_02493__PTR71) );
  MUX2_X1 U9106 ( .A(1'b0), .B(_02651__PTR0), .S(_01766__PTR2), .Z(_02491__PTR64) );
  MUX2_X1 U9107 ( .A(1'b0), .B(_02651__PTR1), .S(_01766__PTR2), .Z(_02491__PTR65) );
  MUX2_X1 U9108 ( .A(1'b0), .B(_02651__PTR2), .S(_01766__PTR2), .Z(_02491__PTR66) );
  MUX2_X1 U9109 ( .A(1'b0), .B(_02651__PTR3), .S(_01766__PTR2), .Z(_02491__PTR67) );
  MUX2_X1 U9110 ( .A(1'b0), .B(_02651__PTR4), .S(_01766__PTR2), .Z(_02491__PTR68) );
  MUX2_X1 U9111 ( .A(1'b0), .B(_02651__PTR5), .S(_01766__PTR2), .Z(_02491__PTR69) );
  MUX2_X1 U9112 ( .A(1'b0), .B(_02651__PTR6), .S(_01766__PTR2), .Z(_02491__PTR70) );
  MUX2_X1 U9113 ( .A(1'b0), .B(_02651__PTR7), .S(_01766__PTR2), .Z(_02491__PTR71) );
  MUX2_X1 U9114 ( .A(1'b0), .B(_02650__PTR0), .S(_01766__PTR2), .Z(_02489__PTR64) );
  MUX2_X1 U9115 ( .A(1'b0), .B(_02650__PTR1), .S(_01766__PTR2), .Z(_02489__PTR65) );
  MUX2_X1 U9116 ( .A(1'b0), .B(_02650__PTR2), .S(_01766__PTR2), .Z(_02489__PTR66) );
  MUX2_X1 U9117 ( .A(1'b0), .B(_02650__PTR3), .S(_01766__PTR2), .Z(_02489__PTR67) );
  MUX2_X1 U9118 ( .A(1'b0), .B(_02650__PTR4), .S(_01766__PTR2), .Z(_02489__PTR68) );
  MUX2_X1 U9119 ( .A(1'b0), .B(_02650__PTR5), .S(_01766__PTR2), .Z(_02489__PTR69) );
  MUX2_X1 U9120 ( .A(1'b0), .B(_02650__PTR6), .S(_01766__PTR2), .Z(_02489__PTR70) );
  MUX2_X1 U9121 ( .A(1'b0), .B(_02650__PTR7), .S(_01766__PTR2), .Z(_02489__PTR71) );
  MUX2_X1 U9122 ( .A(1'b0), .B(_02649__PTR0), .S(_01766__PTR2), .Z(_02487__PTR64) );
  MUX2_X1 U9123 ( .A(1'b0), .B(_02649__PTR1), .S(_01766__PTR2), .Z(_02487__PTR65) );
  MUX2_X1 U9124 ( .A(1'b0), .B(_02649__PTR2), .S(_01766__PTR2), .Z(_02487__PTR66) );
  MUX2_X1 U9125 ( .A(1'b0), .B(_02649__PTR3), .S(_01766__PTR2), .Z(_02487__PTR67) );
  MUX2_X1 U9126 ( .A(1'b0), .B(_02649__PTR4), .S(_01766__PTR2), .Z(_02487__PTR68) );
  MUX2_X1 U9127 ( .A(1'b0), .B(_02649__PTR5), .S(_01766__PTR2), .Z(_02487__PTR69) );
  MUX2_X1 U9128 ( .A(1'b0), .B(_02649__PTR6), .S(_01766__PTR2), .Z(_02487__PTR70) );
  MUX2_X1 U9129 ( .A(1'b0), .B(_02649__PTR7), .S(_01766__PTR2), .Z(_02487__PTR71) );
  MUX2_X1 U9130 ( .A(1'b0), .B(_02648__PTR0), .S(_01766__PTR2), .Z(_02485__PTR64) );
  MUX2_X1 U9131 ( .A(1'b0), .B(_02648__PTR1), .S(_01766__PTR2), .Z(_02485__PTR65) );
  MUX2_X1 U9132 ( .A(1'b0), .B(_02648__PTR2), .S(_01766__PTR2), .Z(_02485__PTR66) );
  MUX2_X1 U9133 ( .A(1'b0), .B(_02648__PTR3), .S(_01766__PTR2), .Z(_02485__PTR67) );
  MUX2_X1 U9134 ( .A(1'b0), .B(_02648__PTR4), .S(_01766__PTR2), .Z(_02485__PTR68) );
  MUX2_X1 U9135 ( .A(1'b0), .B(_02648__PTR5), .S(_01766__PTR2), .Z(_02485__PTR69) );
  MUX2_X1 U9136 ( .A(1'b0), .B(_02648__PTR6), .S(_01766__PTR2), .Z(_02485__PTR70) );
  MUX2_X1 U9137 ( .A(1'b0), .B(_02648__PTR7), .S(_01766__PTR2), .Z(_02485__PTR71) );
  MUX2_X1 U9138 ( .A(1'b0), .B(_02647__PTR0), .S(_01766__PTR2), .Z(_02483__PTR64) );
  MUX2_X1 U9139 ( .A(1'b0), .B(_02647__PTR1), .S(_01766__PTR2), .Z(_02483__PTR65) );
  MUX2_X1 U9140 ( .A(1'b0), .B(_02647__PTR2), .S(_01766__PTR2), .Z(_02483__PTR66) );
  MUX2_X1 U9141 ( .A(1'b0), .B(_02647__PTR3), .S(_01766__PTR2), .Z(_02483__PTR67) );
  MUX2_X1 U9142 ( .A(1'b0), .B(_02647__PTR4), .S(_01766__PTR2), .Z(_02483__PTR68) );
  MUX2_X1 U9143 ( .A(1'b0), .B(_02647__PTR5), .S(_01766__PTR2), .Z(_02483__PTR69) );
  MUX2_X1 U9144 ( .A(1'b0), .B(_02647__PTR6), .S(_01766__PTR2), .Z(_02483__PTR70) );
  MUX2_X1 U9145 ( .A(1'b0), .B(_02647__PTR7), .S(_01766__PTR2), .Z(_02483__PTR71) );
  MUX2_X1 U9146 ( .A(1'b0), .B(_02646__PTR0), .S(_01766__PTR2), .Z(_02481__PTR64) );
  MUX2_X1 U9147 ( .A(1'b0), .B(_02646__PTR1), .S(_01766__PTR2), .Z(_02481__PTR65) );
  MUX2_X1 U9148 ( .A(1'b0), .B(_02646__PTR2), .S(_01766__PTR2), .Z(_02481__PTR66) );
  MUX2_X1 U9149 ( .A(1'b0), .B(_02646__PTR3), .S(_01766__PTR2), .Z(_02481__PTR67) );
  MUX2_X1 U9150 ( .A(1'b0), .B(_02646__PTR4), .S(_01766__PTR2), .Z(_02481__PTR68) );
  MUX2_X1 U9151 ( .A(1'b0), .B(_02646__PTR5), .S(_01766__PTR2), .Z(_02481__PTR69) );
  MUX2_X1 U9152 ( .A(1'b0), .B(_02646__PTR6), .S(_01766__PTR2), .Z(_02481__PTR70) );
  MUX2_X1 U9153 ( .A(1'b0), .B(_02646__PTR7), .S(_01766__PTR2), .Z(_02481__PTR71) );
  MUX2_X1 U9154 ( .A(1'b0), .B(_02645__PTR0), .S(_01766__PTR2), .Z(_02479__PTR64) );
  MUX2_X1 U9155 ( .A(1'b0), .B(_02645__PTR1), .S(_01766__PTR2), .Z(_02479__PTR65) );
  MUX2_X1 U9156 ( .A(1'b0), .B(_02645__PTR2), .S(_01766__PTR2), .Z(_02479__PTR66) );
  MUX2_X1 U9157 ( .A(1'b0), .B(_02645__PTR3), .S(_01766__PTR2), .Z(_02479__PTR67) );
  MUX2_X1 U9158 ( .A(1'b0), .B(_02645__PTR4), .S(_01766__PTR2), .Z(_02479__PTR68) );
  MUX2_X1 U9159 ( .A(1'b0), .B(_02645__PTR5), .S(_01766__PTR2), .Z(_02479__PTR69) );
  MUX2_X1 U9160 ( .A(1'b0), .B(_02645__PTR6), .S(_01766__PTR2), .Z(_02479__PTR70) );
  MUX2_X1 U9161 ( .A(1'b0), .B(_02645__PTR7), .S(_01766__PTR2), .Z(_02479__PTR71) );
  MUX2_X1 U9162 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR0), .Z(_02660__PTR0) );
  MUX2_X1 U9163 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR0), .Z(_02660__PTR1) );
  MUX2_X1 U9164 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR0), .Z(_02660__PTR2) );
  MUX2_X1 U9165 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR0), .Z(_02660__PTR3) );
  MUX2_X1 U9166 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR0), .Z(_02660__PTR4) );
  MUX2_X1 U9167 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR0), .Z(_02660__PTR5) );
  MUX2_X1 U9168 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR0), .Z(_02660__PTR6) );
  MUX2_X1 U9169 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR0), .Z(_02660__PTR7) );
  MUX2_X1 U9170 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR1), .Z(_02659__PTR0) );
  MUX2_X1 U9171 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR1), .Z(_02659__PTR1) );
  MUX2_X1 U9172 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR1), .Z(_02659__PTR2) );
  MUX2_X1 U9173 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR1), .Z(_02659__PTR3) );
  MUX2_X1 U9174 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR1), .Z(_02659__PTR4) );
  MUX2_X1 U9175 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR1), .Z(_02659__PTR5) );
  MUX2_X1 U9176 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR1), .Z(_02659__PTR6) );
  MUX2_X1 U9177 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR1), .Z(_02659__PTR7) );
  MUX2_X1 U9178 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR2), .Z(_02658__PTR0) );
  MUX2_X1 U9179 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR2), .Z(_02658__PTR1) );
  MUX2_X1 U9180 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR2), .Z(_02658__PTR2) );
  MUX2_X1 U9181 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR2), .Z(_02658__PTR3) );
  MUX2_X1 U9182 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR2), .Z(_02658__PTR4) );
  MUX2_X1 U9183 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR2), .Z(_02658__PTR5) );
  MUX2_X1 U9184 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR2), .Z(_02658__PTR6) );
  MUX2_X1 U9185 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR2), .Z(_02658__PTR7) );
  MUX2_X1 U9186 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR3), .Z(_02657__PTR0) );
  MUX2_X1 U9187 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR3), .Z(_02657__PTR1) );
  MUX2_X1 U9188 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR3), .Z(_02657__PTR2) );
  MUX2_X1 U9189 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR3), .Z(_02657__PTR3) );
  MUX2_X1 U9190 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR3), .Z(_02657__PTR4) );
  MUX2_X1 U9191 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR3), .Z(_02657__PTR5) );
  MUX2_X1 U9192 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR3), .Z(_02657__PTR6) );
  MUX2_X1 U9193 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR3), .Z(_02657__PTR7) );
  MUX2_X1 U9194 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR4), .Z(_02656__PTR0) );
  MUX2_X1 U9195 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR4), .Z(_02656__PTR1) );
  MUX2_X1 U9196 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR4), .Z(_02656__PTR2) );
  MUX2_X1 U9197 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR4), .Z(_02656__PTR3) );
  MUX2_X1 U9198 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR4), .Z(_02656__PTR4) );
  MUX2_X1 U9199 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR4), .Z(_02656__PTR5) );
  MUX2_X1 U9200 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR4), .Z(_02656__PTR6) );
  MUX2_X1 U9201 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR4), .Z(_02656__PTR7) );
  MUX2_X1 U9202 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR5), .Z(_02655__PTR0) );
  MUX2_X1 U9203 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR5), .Z(_02655__PTR1) );
  MUX2_X1 U9204 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR5), .Z(_02655__PTR2) );
  MUX2_X1 U9205 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR5), .Z(_02655__PTR3) );
  MUX2_X1 U9206 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR5), .Z(_02655__PTR4) );
  MUX2_X1 U9207 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR5), .Z(_02655__PTR5) );
  MUX2_X1 U9208 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR5), .Z(_02655__PTR6) );
  MUX2_X1 U9209 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR5), .Z(_02655__PTR7) );
  MUX2_X1 U9210 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR6), .Z(_02654__PTR0) );
  MUX2_X1 U9211 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR6), .Z(_02654__PTR1) );
  MUX2_X1 U9212 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR6), .Z(_02654__PTR2) );
  MUX2_X1 U9213 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR6), .Z(_02654__PTR3) );
  MUX2_X1 U9214 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR6), .Z(_02654__PTR4) );
  MUX2_X1 U9215 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR6), .Z(_02654__PTR5) );
  MUX2_X1 U9216 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR6), .Z(_02654__PTR6) );
  MUX2_X1 U9217 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR6), .Z(_02654__PTR7) );
  MUX2_X1 U9218 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR7), .Z(_02653__PTR0) );
  MUX2_X1 U9219 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR7), .Z(_02653__PTR1) );
  MUX2_X1 U9220 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR7), .Z(_02653__PTR2) );
  MUX2_X1 U9221 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR7), .Z(_02653__PTR3) );
  MUX2_X1 U9222 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR7), .Z(_02653__PTR4) );
  MUX2_X1 U9223 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR7), .Z(_02653__PTR5) );
  MUX2_X1 U9224 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR7), .Z(_02653__PTR6) );
  MUX2_X1 U9225 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR7), .Z(_02653__PTR7) );
  MUX2_X1 U9226 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR8), .Z(_02652__PTR0) );
  MUX2_X1 U9227 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR8), .Z(_02652__PTR1) );
  MUX2_X1 U9228 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR8), .Z(_02652__PTR2) );
  MUX2_X1 U9229 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR8), .Z(_02652__PTR3) );
  MUX2_X1 U9230 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR8), .Z(_02652__PTR4) );
  MUX2_X1 U9231 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR8), .Z(_02652__PTR5) );
  MUX2_X1 U9232 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR8), .Z(_02652__PTR6) );
  MUX2_X1 U9233 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR8), .Z(_02652__PTR7) );
  MUX2_X1 U9234 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR9), .Z(_02651__PTR0) );
  MUX2_X1 U9235 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR9), .Z(_02651__PTR1) );
  MUX2_X1 U9236 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR9), .Z(_02651__PTR2) );
  MUX2_X1 U9237 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR9), .Z(_02651__PTR3) );
  MUX2_X1 U9238 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR9), .Z(_02651__PTR4) );
  MUX2_X1 U9239 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR9), .Z(_02651__PTR5) );
  MUX2_X1 U9240 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR9), .Z(_02651__PTR6) );
  MUX2_X1 U9241 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR9), .Z(_02651__PTR7) );
  MUX2_X1 U9242 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR10), .Z(_02650__PTR0) );
  MUX2_X1 U9243 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR10), .Z(_02650__PTR1) );
  MUX2_X1 U9244 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR10), .Z(_02650__PTR2) );
  MUX2_X1 U9245 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR10), .Z(_02650__PTR3) );
  MUX2_X1 U9246 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR10), .Z(_02650__PTR4) );
  MUX2_X1 U9247 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR10), .Z(_02650__PTR5) );
  MUX2_X1 U9248 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR10), .Z(_02650__PTR6) );
  MUX2_X1 U9249 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR10), .Z(_02650__PTR7) );
  MUX2_X1 U9250 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR11), .Z(_02649__PTR0) );
  MUX2_X1 U9251 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR11), .Z(_02649__PTR1) );
  MUX2_X1 U9252 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR11), .Z(_02649__PTR2) );
  MUX2_X1 U9253 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR11), .Z(_02649__PTR3) );
  MUX2_X1 U9254 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR11), .Z(_02649__PTR4) );
  MUX2_X1 U9255 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR11), .Z(_02649__PTR5) );
  MUX2_X1 U9256 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR11), .Z(_02649__PTR6) );
  MUX2_X1 U9257 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR11), .Z(_02649__PTR7) );
  MUX2_X1 U9258 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR12), .Z(_02648__PTR0) );
  MUX2_X1 U9259 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR12), .Z(_02648__PTR1) );
  MUX2_X1 U9260 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR12), .Z(_02648__PTR2) );
  MUX2_X1 U9261 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR12), .Z(_02648__PTR3) );
  MUX2_X1 U9262 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR12), .Z(_02648__PTR4) );
  MUX2_X1 U9263 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR12), .Z(_02648__PTR5) );
  MUX2_X1 U9264 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR12), .Z(_02648__PTR6) );
  MUX2_X1 U9265 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR12), .Z(_02648__PTR7) );
  MUX2_X1 U9266 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR13), .Z(_02647__PTR0) );
  MUX2_X1 U9267 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR13), .Z(_02647__PTR1) );
  MUX2_X1 U9268 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR13), .Z(_02647__PTR2) );
  MUX2_X1 U9269 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR13), .Z(_02647__PTR3) );
  MUX2_X1 U9270 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR13), .Z(_02647__PTR4) );
  MUX2_X1 U9271 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR13), .Z(_02647__PTR5) );
  MUX2_X1 U9272 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR13), .Z(_02647__PTR6) );
  MUX2_X1 U9273 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR13), .Z(_02647__PTR7) );
  MUX2_X1 U9274 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR14), .Z(_02646__PTR0) );
  MUX2_X1 U9275 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR14), .Z(_02646__PTR1) );
  MUX2_X1 U9276 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR14), .Z(_02646__PTR2) );
  MUX2_X1 U9277 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR14), .Z(_02646__PTR3) );
  MUX2_X1 U9278 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR14), .Z(_02646__PTR4) );
  MUX2_X1 U9279 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR14), .Z(_02646__PTR5) );
  MUX2_X1 U9280 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR14), .Z(_02646__PTR6) );
  MUX2_X1 U9281 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR14), .Z(_02646__PTR7) );
  MUX2_X1 U9282 ( .A(1'b0), .B(_02464__PTR0), .S(_02417__PTR15), .Z(_02645__PTR0) );
  MUX2_X1 U9283 ( .A(1'b0), .B(_02464__PTR1), .S(_02417__PTR15), .Z(_02645__PTR1) );
  MUX2_X1 U9284 ( .A(1'b0), .B(_02464__PTR2), .S(_02417__PTR15), .Z(_02645__PTR2) );
  MUX2_X1 U9285 ( .A(1'b0), .B(_02464__PTR3), .S(_02417__PTR15), .Z(_02645__PTR3) );
  MUX2_X1 U9286 ( .A(1'b0), .B(_02464__PTR4), .S(_02417__PTR15), .Z(_02645__PTR4) );
  MUX2_X1 U9287 ( .A(1'b0), .B(_02464__PTR5), .S(_02417__PTR15), .Z(_02645__PTR5) );
  MUX2_X1 U9288 ( .A(1'b0), .B(_02464__PTR6), .S(_02417__PTR15), .Z(_02645__PTR6) );
  MUX2_X1 U9289 ( .A(1'b0), .B(_02464__PTR7), .S(_02417__PTR15), .Z(_02645__PTR7) );
  MUX2_X1 U9290 ( .A(1'b0), .B(_02644__PTR0), .S(_02475__PTR28), .Z(_02511__PTR56) );
  MUX2_X1 U9291 ( .A(1'b0), .B(_02644__PTR4), .S(_02475__PTR28), .Z(_02511__PTR60) );
  MUX2_X1 U9292 ( .A(1'b0), .B(1'b1), .S(P3_P1_Flush), .Z(_02644__PTR0) );
  MUX2_X1 U9293 ( .A(1'b0), .B(1'b0), .S(P3_P1_Flush), .Z(_02644__PTR4) );
  MUX2_X1 U9294 ( .A(P3_P1_InstQueueRd_Addr_PTR0), .B(_02643__PTR0), .S(P3_P1_Flush), .Z(_02513__PTR56) );
  MUX2_X1 U9295 ( .A(P3_P1_InstQueueRd_Addr_PTR1), .B(_02643__PTR1), .S(P3_P1_Flush), .Z(_02513__PTR57) );
  MUX2_X1 U9296 ( .A(P3_P1_InstQueueRd_Addr_PTR2), .B(_02643__PTR2), .S(P3_P1_Flush), .Z(_02513__PTR58) );
  MUX2_X1 U9297 ( .A(P3_P1_InstQueueRd_Addr_PTR3), .B(1'b0), .S(P3_P1_Flush), .Z(_02513__PTR59) );
  MUX2_X1 U9298 ( .A(P3_P1_InstQueueRd_Addr_PTR4), .B(1'b0), .S(P3_P1_Flush), .Z(_02513__PTR60) );
  MUX2_X1 U9299 ( .A(1'b1), .B(_02662__PTR0), .S(P3_P1_InstAddrPointer_PTR0), .Z(_02643__PTR0) );
  MUX2_X1 U9300 ( .A(1'b0), .B(_03321__PTR1), .S(P3_P1_InstAddrPointer_PTR0), .Z(_02643__PTR1) );
  MUX2_X1 U9301 ( .A(1'b0), .B(_03320__PTR1), .S(P3_P1_InstAddrPointer_PTR0), .Z(_02643__PTR2) );
  MUX2_X1 U9302 ( .A(_03439__PTR1), .B(P3_P1_InstAddrPointer_PTR1), .S(_03234__PTR31), .Z(_03319__PTR1) );
  MUX2_X1 U9303 ( .A(1'b1), .B(1'b0), .S(P3_READY_n), .Z(_02475__PTR26) );
  MUX2_X1 U9304 ( .A(1'b0), .B(1'b0), .S(P3_READY_n), .Z(_02431__PTR6) );
  MUX2_X1 U9305 ( .A(_02699__PTR0), .B(1'b1), .S(_02642_), .Z(_02475__PTR20) );
  MUX2_X1 U9306 ( .A(_02699__PTR1), .B(1'b1), .S(_02642_), .Z(_02475__PTR21) );
  MUX2_X1 U9307 ( .A(_02699__PTR2), .B(1'b1), .S(_02642_), .Z(_02475__PTR22) );
  MUX2_X1 U9308 ( .A(_02699__PTR3), .B(1'b0), .S(_02642_), .Z(_02475__PTR23) );
  MUX2_X1 U9309 ( .A(P3_Datao_PTR16), .B(_02625__PTR16), .S(_02585_), .Z(_02692__PTR48) );
  MUX2_X1 U9310 ( .A(P3_Datao_PTR17), .B(_02625__PTR17), .S(_02585_), .Z(_02692__PTR49) );
  MUX2_X1 U9311 ( .A(P3_Datao_PTR18), .B(_02625__PTR18), .S(_02585_), .Z(_02692__PTR50) );
  MUX2_X1 U9312 ( .A(P3_Datao_PTR19), .B(_02625__PTR19), .S(_02585_), .Z(_02692__PTR51) );
  MUX2_X1 U9313 ( .A(P3_Datao_PTR20), .B(_02625__PTR20), .S(_02585_), .Z(_02692__PTR52) );
  MUX2_X1 U9314 ( .A(P3_Datao_PTR21), .B(_02625__PTR21), .S(_02585_), .Z(_02692__PTR53) );
  MUX2_X1 U9315 ( .A(P3_Datao_PTR22), .B(_02625__PTR22), .S(_02585_), .Z(_02692__PTR54) );
  MUX2_X1 U9316 ( .A(P3_Datao_PTR23), .B(_02625__PTR23), .S(_02585_), .Z(_02692__PTR55) );
  MUX2_X1 U9317 ( .A(P3_Datao_PTR24), .B(_02625__PTR24), .S(_02585_), .Z(_02692__PTR56) );
  MUX2_X1 U9318 ( .A(P3_Datao_PTR25), .B(_02625__PTR25), .S(_02585_), .Z(_02692__PTR57) );
  MUX2_X1 U9319 ( .A(P3_Datao_PTR26), .B(_02625__PTR26), .S(_02585_), .Z(_02692__PTR58) );
  MUX2_X1 U9320 ( .A(P3_Datao_PTR27), .B(_02625__PTR27), .S(_02585_), .Z(_02692__PTR59) );
  MUX2_X1 U9321 ( .A(P3_Datao_PTR28), .B(_02625__PTR28), .S(_02585_), .Z(_02692__PTR60) );
  MUX2_X1 U9322 ( .A(P3_Datao_PTR29), .B(_02625__PTR29), .S(_02585_), .Z(_02692__PTR61) );
  MUX2_X1 U9323 ( .A(P3_Datao_PTR30), .B(_02625__PTR30), .S(_02585_), .Z(_02692__PTR62) );
  MUX2_X1 U9324 ( .A(P3_Datao_PTR31), .B(_02610__PTR31), .S(_02585_), .Z(_02692__PTR95) );
  MUX2_X1 U9325 ( .A(P3_Datao_PTR0), .B(_02610__PTR0), .S(_02585_), .Z(_02692__PTR64) );
  MUX2_X1 U9326 ( .A(P3_Datao_PTR1), .B(_02610__PTR1), .S(_02585_), .Z(_02692__PTR65) );
  MUX2_X1 U9327 ( .A(P3_Datao_PTR2), .B(_02610__PTR2), .S(_02585_), .Z(_02692__PTR66) );
  MUX2_X1 U9328 ( .A(P3_Datao_PTR3), .B(_02610__PTR3), .S(_02585_), .Z(_02692__PTR67) );
  MUX2_X1 U9329 ( .A(P3_Datao_PTR4), .B(_02610__PTR4), .S(_02585_), .Z(_02692__PTR68) );
  MUX2_X1 U9330 ( .A(P3_Datao_PTR5), .B(_02610__PTR5), .S(_02585_), .Z(_02692__PTR69) );
  MUX2_X1 U9331 ( .A(P3_Datao_PTR6), .B(_02610__PTR6), .S(_02585_), .Z(_02692__PTR70) );
  MUX2_X1 U9332 ( .A(P3_Datao_PTR7), .B(_02610__PTR7), .S(_02585_), .Z(_02692__PTR71) );
  MUX2_X1 U9333 ( .A(P3_Datao_PTR8), .B(_02610__PTR8), .S(_02585_), .Z(_02692__PTR72) );
  MUX2_X1 U9334 ( .A(P3_Datao_PTR9), .B(_02610__PTR9), .S(_02585_), .Z(_02692__PTR73) );
  MUX2_X1 U9335 ( .A(P3_Datao_PTR10), .B(_02610__PTR10), .S(_02585_), .Z(_02692__PTR74) );
  MUX2_X1 U9336 ( .A(P3_Datao_PTR11), .B(_02610__PTR11), .S(_02585_), .Z(_02692__PTR75) );
  MUX2_X1 U9337 ( .A(P3_Datao_PTR12), .B(_02610__PTR12), .S(_02585_), .Z(_02692__PTR76) );
  MUX2_X1 U9338 ( .A(P3_Datao_PTR13), .B(_02610__PTR13), .S(_02585_), .Z(_02692__PTR77) );
  MUX2_X1 U9339 ( .A(P3_Datao_PTR14), .B(_02610__PTR14), .S(_02585_), .Z(_02692__PTR78) );
  MUX2_X1 U9340 ( .A(P3_Datao_PTR15), .B(_02610__PTR15), .S(_02585_), .Z(_02692__PTR79) );
  MUX2_X1 U9341 ( .A(P3_Datao_PTR16), .B(_02610__PTR16), .S(_02585_), .Z(_02692__PTR80) );
  MUX2_X1 U9342 ( .A(P3_Datao_PTR17), .B(_02610__PTR17), .S(_02585_), .Z(_02692__PTR81) );
  MUX2_X1 U9343 ( .A(P3_Datao_PTR18), .B(_02610__PTR18), .S(_02585_), .Z(_02692__PTR82) );
  MUX2_X1 U9344 ( .A(P3_Datao_PTR19), .B(_02610__PTR19), .S(_02585_), .Z(_02692__PTR83) );
  MUX2_X1 U9345 ( .A(P3_Datao_PTR20), .B(_02610__PTR20), .S(_02585_), .Z(_02692__PTR84) );
  MUX2_X1 U9346 ( .A(P3_Datao_PTR21), .B(_02610__PTR21), .S(_02585_), .Z(_02692__PTR85) );
  MUX2_X1 U9347 ( .A(P3_Datao_PTR22), .B(_02610__PTR22), .S(_02585_), .Z(_02692__PTR86) );
  MUX2_X1 U9348 ( .A(P3_Datao_PTR23), .B(_02610__PTR23), .S(_02585_), .Z(_02692__PTR87) );
  MUX2_X1 U9349 ( .A(P3_Datao_PTR24), .B(_02610__PTR24), .S(_02585_), .Z(_02692__PTR88) );
  MUX2_X1 U9350 ( .A(P3_Datao_PTR25), .B(_02610__PTR25), .S(_02585_), .Z(_02692__PTR89) );
  MUX2_X1 U9351 ( .A(P3_Datao_PTR26), .B(_02610__PTR26), .S(_02585_), .Z(_02692__PTR90) );
  MUX2_X1 U9352 ( .A(P3_Datao_PTR27), .B(_02610__PTR27), .S(_02585_), .Z(_02692__PTR91) );
  MUX2_X1 U9353 ( .A(P3_Datao_PTR28), .B(_02610__PTR28), .S(_02585_), .Z(_02692__PTR92) );
  MUX2_X1 U9354 ( .A(P3_Datao_PTR29), .B(_02610__PTR29), .S(_02585_), .Z(_02692__PTR93) );
  MUX2_X1 U9355 ( .A(P3_Datao_PTR30), .B(_02610__PTR30), .S(_02585_), .Z(_02692__PTR94) );
  MUX2_X1 U9356 ( .A(P3_RequestPending), .B(_02626_), .S(_02585_), .Z(_02443__PTR0) );
  MUX2_X1 U9357 ( .A(1'b1), .B(P3_READY_n), .S(_02604_), .Z(_02626_) );
  MUX2_X1 U9358 ( .A(P3_MemoryFetch), .B(1'b0), .S(_02585_), .Z(_02450__PTR0) );
  MUX2_X1 U9359 ( .A(1'b0), .B(_02615_), .S(_02585_), .Z(_02435__PTR0) );
  MUX2_X1 U9360 ( .A(1'b1), .B(_02614_), .S(_02585_), .Z(_02439__PTR0) );
  MUX2_X1 U9361 ( .A(P3_P1_State2_PTR0), .B(_02613__PTR0), .S(_02585_), .Z(_02696__PTR4) );
  MUX2_X1 U9362 ( .A(P3_P1_State2_PTR1), .B(_02613__PTR1), .S(_02585_), .Z(_02696__PTR5) );
  MUX2_X1 U9363 ( .A(P3_P1_State2_PTR2), .B(_02613__PTR2), .S(_02585_), .Z(_02696__PTR6) );
  MUX2_X1 U9364 ( .A(P3_P1_State2_PTR3), .B(_02613__PTR3), .S(_02585_), .Z(_02696__PTR7) );
  MUX2_X1 U9365 ( .A(P3_Datao_PTR16), .B(1'b0), .S(_02604_), .Z(_02625__PTR16) );
  MUX2_X1 U9366 ( .A(P3_Datao_PTR17), .B(1'b0), .S(_02604_), .Z(_02625__PTR17) );
  MUX2_X1 U9367 ( .A(P3_Datao_PTR18), .B(1'b0), .S(_02604_), .Z(_02625__PTR18) );
  MUX2_X1 U9368 ( .A(P3_Datao_PTR19), .B(1'b0), .S(_02604_), .Z(_02625__PTR19) );
  MUX2_X1 U9369 ( .A(P3_Datao_PTR20), .B(1'b0), .S(_02604_), .Z(_02625__PTR20) );
  MUX2_X1 U9370 ( .A(P3_Datao_PTR21), .B(1'b0), .S(_02604_), .Z(_02625__PTR21) );
  MUX2_X1 U9371 ( .A(P3_Datao_PTR22), .B(1'b0), .S(_02604_), .Z(_02625__PTR22) );
  MUX2_X1 U9372 ( .A(P3_Datao_PTR23), .B(1'b0), .S(_02604_), .Z(_02625__PTR23) );
  MUX2_X1 U9373 ( .A(P3_Datao_PTR24), .B(1'b0), .S(_02604_), .Z(_02625__PTR24) );
  MUX2_X1 U9374 ( .A(P3_Datao_PTR25), .B(1'b0), .S(_02604_), .Z(_02625__PTR25) );
  MUX2_X1 U9375 ( .A(P3_Datao_PTR26), .B(1'b0), .S(_02604_), .Z(_02625__PTR26) );
  MUX2_X1 U9376 ( .A(P3_Datao_PTR27), .B(1'b0), .S(_02604_), .Z(_02625__PTR27) );
  MUX2_X1 U9377 ( .A(P3_Datao_PTR28), .B(1'b0), .S(_02604_), .Z(_02625__PTR28) );
  MUX2_X1 U9378 ( .A(P3_Datao_PTR29), .B(1'b0), .S(_02604_), .Z(_02625__PTR29) );
  MUX2_X1 U9379 ( .A(P3_Datao_PTR30), .B(1'b0), .S(_02604_), .Z(_02625__PTR30) );
  MUX2_X1 U9380 ( .A(P3_Datao_PTR31), .B(1'b0), .S(_02604_), .Z(_02610__PTR31) );
  MUX2_X1 U9381 ( .A(P3_Datao_PTR0), .B(P3_EAX_PTR0), .S(_02604_), .Z(_02610__PTR0) );
  MUX2_X1 U9382 ( .A(P3_Datao_PTR1), .B(P3_EAX_PTR1), .S(_02604_), .Z(_02610__PTR1) );
  MUX2_X1 U9383 ( .A(P3_Datao_PTR2), .B(P3_EAX_PTR2), .S(_02604_), .Z(_02610__PTR2) );
  MUX2_X1 U9384 ( .A(P3_Datao_PTR3), .B(P3_EAX_PTR3), .S(_02604_), .Z(_02610__PTR3) );
  MUX2_X1 U9385 ( .A(P3_Datao_PTR4), .B(P3_EAX_PTR4), .S(_02604_), .Z(_02610__PTR4) );
  MUX2_X1 U9386 ( .A(P3_Datao_PTR5), .B(P3_EAX_PTR5), .S(_02604_), .Z(_02610__PTR5) );
  MUX2_X1 U9387 ( .A(P3_Datao_PTR6), .B(P3_EAX_PTR6), .S(_02604_), .Z(_02610__PTR6) );
  MUX2_X1 U9388 ( .A(P3_Datao_PTR7), .B(P3_EAX_PTR7), .S(_02604_), .Z(_02610__PTR7) );
  MUX2_X1 U9389 ( .A(P3_Datao_PTR8), .B(P3_EAX_PTR8), .S(_02604_), .Z(_02610__PTR8) );
  MUX2_X1 U9390 ( .A(P3_Datao_PTR9), .B(P3_EAX_PTR9), .S(_02604_), .Z(_02610__PTR9) );
  MUX2_X1 U9391 ( .A(P3_Datao_PTR10), .B(P3_EAX_PTR10), .S(_02604_), .Z(_02610__PTR10) );
  MUX2_X1 U9392 ( .A(P3_Datao_PTR11), .B(P3_EAX_PTR11), .S(_02604_), .Z(_02610__PTR11) );
  MUX2_X1 U9393 ( .A(P3_Datao_PTR12), .B(P3_EAX_PTR12), .S(_02604_), .Z(_02610__PTR12) );
  MUX2_X1 U9394 ( .A(P3_Datao_PTR13), .B(P3_EAX_PTR13), .S(_02604_), .Z(_02610__PTR13) );
  MUX2_X1 U9395 ( .A(P3_Datao_PTR14), .B(P3_EAX_PTR14), .S(_02604_), .Z(_02610__PTR14) );
  MUX2_X1 U9396 ( .A(P3_Datao_PTR15), .B(P3_EAX_PTR15), .S(_02604_), .Z(_02610__PTR15) );
  MUX2_X1 U9397 ( .A(P3_Datao_PTR16), .B(_03315__PTR0), .S(_02604_), .Z(_02610__PTR16) );
  MUX2_X1 U9398 ( .A(P3_Datao_PTR17), .B(_03316__PTR1), .S(_02604_), .Z(_02610__PTR17) );
  MUX2_X1 U9399 ( .A(P3_Datao_PTR18), .B(_03316__PTR2), .S(_02604_), .Z(_02610__PTR18) );
  MUX2_X1 U9400 ( .A(P3_Datao_PTR19), .B(_03316__PTR3), .S(_02604_), .Z(_02610__PTR19) );
  MUX2_X1 U9401 ( .A(P3_Datao_PTR20), .B(_03316__PTR4), .S(_02604_), .Z(_02610__PTR20) );
  MUX2_X1 U9402 ( .A(P3_Datao_PTR21), .B(_03316__PTR5), .S(_02604_), .Z(_02610__PTR21) );
  MUX2_X1 U9403 ( .A(P3_Datao_PTR22), .B(_03316__PTR6), .S(_02604_), .Z(_02610__PTR22) );
  MUX2_X1 U9404 ( .A(P3_Datao_PTR23), .B(_03316__PTR7), .S(_02604_), .Z(_02610__PTR23) );
  MUX2_X1 U9405 ( .A(P3_Datao_PTR24), .B(_03316__PTR8), .S(_02604_), .Z(_02610__PTR24) );
  MUX2_X1 U9406 ( .A(P3_Datao_PTR25), .B(_03316__PTR9), .S(_02604_), .Z(_02610__PTR25) );
  MUX2_X1 U9407 ( .A(P3_Datao_PTR26), .B(_03316__PTR10), .S(_02604_), .Z(_02610__PTR26) );
  MUX2_X1 U9408 ( .A(P3_Datao_PTR27), .B(_03316__PTR11), .S(_02604_), .Z(_02610__PTR27) );
  MUX2_X1 U9409 ( .A(P3_Datao_PTR28), .B(_03316__PTR12), .S(_02604_), .Z(_02610__PTR28) );
  MUX2_X1 U9410 ( .A(P3_Datao_PTR29), .B(_03316__PTR13), .S(_02604_), .Z(_02610__PTR29) );
  MUX2_X1 U9411 ( .A(P3_Datao_PTR30), .B(_03316__PTR14), .S(_02604_), .Z(_02610__PTR30) );
  MUX2_X1 U9412 ( .A(P3_ReadRequest), .B(1'b0), .S(_02585_), .Z(_02447__PTR0) );
  MUX2_X1 U9413 ( .A(P3_RequestPending), .B(_02611_), .S(_02585_), .Z(_02443__PTR2) );
  MUX2_X1 U9414 ( .A(P3_P1_InstQueueRd_Addr_PTR1), .B(_02599__PTR1), .S(_02604_), .Z(_02617__PTR1) );
  MUX2_X1 U9415 ( .A(P3_P1_InstQueueRd_Addr_PTR2), .B(_02599__PTR2), .S(_02604_), .Z(_02617__PTR2) );
  MUX2_X1 U9416 ( .A(P3_P1_InstQueueRd_Addr_PTR3), .B(_02599__PTR3), .S(_02604_), .Z(_02617__PTR3) );
  MUX2_X1 U9417 ( .A(P3_P1_InstQueueRd_Addr_PTR4), .B(_02599__PTR4), .S(_02604_), .Z(_02617__PTR4) );
  MUX2_X1 U9418 ( .A(P3_P1_InstAddrPointer_PTR1), .B(_02598__PTR1), .S(_02604_), .Z(_02616__PTR1) );
  MUX2_X1 U9419 ( .A(P3_P1_InstAddrPointer_PTR2), .B(_02598__PTR2), .S(_02604_), .Z(_02616__PTR2) );
  MUX2_X1 U9420 ( .A(P3_P1_InstAddrPointer_PTR3), .B(_02598__PTR3), .S(_02604_), .Z(_02616__PTR3) );
  MUX2_X1 U9421 ( .A(P3_P1_InstAddrPointer_PTR4), .B(_02598__PTR4), .S(_02604_), .Z(_02616__PTR4) );
  MUX2_X1 U9422 ( .A(P3_P1_InstAddrPointer_PTR5), .B(_02598__PTR5), .S(_02604_), .Z(_02616__PTR5) );
  MUX2_X1 U9423 ( .A(P3_P1_InstAddrPointer_PTR6), .B(_02598__PTR6), .S(_02604_), .Z(_02616__PTR6) );
  MUX2_X1 U9424 ( .A(P3_P1_InstAddrPointer_PTR7), .B(_02598__PTR7), .S(_02604_), .Z(_02616__PTR7) );
  MUX2_X1 U9425 ( .A(P3_P1_InstAddrPointer_PTR8), .B(_02598__PTR8), .S(_02604_), .Z(_02616__PTR8) );
  MUX2_X1 U9426 ( .A(P3_P1_InstAddrPointer_PTR9), .B(_02598__PTR9), .S(_02604_), .Z(_02616__PTR9) );
  MUX2_X1 U9427 ( .A(P3_P1_InstAddrPointer_PTR10), .B(_02598__PTR10), .S(_02604_), .Z(_02616__PTR10) );
  MUX2_X1 U9428 ( .A(P3_P1_InstAddrPointer_PTR11), .B(_02598__PTR11), .S(_02604_), .Z(_02616__PTR11) );
  MUX2_X1 U9429 ( .A(P3_P1_InstAddrPointer_PTR12), .B(_02598__PTR12), .S(_02604_), .Z(_02616__PTR12) );
  MUX2_X1 U9430 ( .A(P3_P1_InstAddrPointer_PTR13), .B(_02598__PTR13), .S(_02604_), .Z(_02616__PTR13) );
  MUX2_X1 U9431 ( .A(P3_P1_InstAddrPointer_PTR14), .B(_02598__PTR14), .S(_02604_), .Z(_02616__PTR14) );
  MUX2_X1 U9432 ( .A(P3_P1_InstAddrPointer_PTR15), .B(_02598__PTR15), .S(_02604_), .Z(_02616__PTR15) );
  MUX2_X1 U9433 ( .A(P3_P1_InstAddrPointer_PTR16), .B(_02598__PTR16), .S(_02604_), .Z(_02616__PTR16) );
  MUX2_X1 U9434 ( .A(P3_P1_InstAddrPointer_PTR17), .B(_02598__PTR17), .S(_02604_), .Z(_02616__PTR17) );
  MUX2_X1 U9435 ( .A(P3_P1_InstAddrPointer_PTR18), .B(_02598__PTR18), .S(_02604_), .Z(_02616__PTR18) );
  MUX2_X1 U9436 ( .A(P3_P1_InstAddrPointer_PTR19), .B(_02598__PTR19), .S(_02604_), .Z(_02616__PTR19) );
  MUX2_X1 U9437 ( .A(P3_P1_InstAddrPointer_PTR20), .B(_02598__PTR20), .S(_02604_), .Z(_02616__PTR20) );
  MUX2_X1 U9438 ( .A(P3_P1_InstAddrPointer_PTR21), .B(_02598__PTR21), .S(_02604_), .Z(_02616__PTR21) );
  MUX2_X1 U9439 ( .A(P3_P1_InstAddrPointer_PTR22), .B(_02598__PTR22), .S(_02604_), .Z(_02616__PTR22) );
  MUX2_X1 U9440 ( .A(P3_P1_InstAddrPointer_PTR23), .B(_02598__PTR23), .S(_02604_), .Z(_02616__PTR23) );
  MUX2_X1 U9441 ( .A(P3_P1_InstAddrPointer_PTR24), .B(_02598__PTR24), .S(_02604_), .Z(_02616__PTR24) );
  MUX2_X1 U9442 ( .A(P3_P1_InstAddrPointer_PTR25), .B(_02598__PTR25), .S(_02604_), .Z(_02616__PTR25) );
  MUX2_X1 U9443 ( .A(P3_P1_InstAddrPointer_PTR26), .B(_02598__PTR26), .S(_02604_), .Z(_02616__PTR26) );
  MUX2_X1 U9444 ( .A(P3_P1_InstAddrPointer_PTR27), .B(_02598__PTR27), .S(_02604_), .Z(_02616__PTR27) );
  MUX2_X1 U9445 ( .A(P3_P1_InstAddrPointer_PTR28), .B(_02598__PTR28), .S(_02604_), .Z(_02616__PTR28) );
  MUX2_X1 U9446 ( .A(P3_P1_InstAddrPointer_PTR29), .B(_02598__PTR29), .S(_02604_), .Z(_02616__PTR29) );
  MUX2_X1 U9447 ( .A(P3_P1_InstAddrPointer_PTR30), .B(_02598__PTR30), .S(_02604_), .Z(_02616__PTR30) );
  MUX2_X1 U9448 ( .A(P3_P1_InstAddrPointer_PTR31), .B(_02598__PTR31), .S(_02604_), .Z(_02616__PTR31) );
  MUX2_X1 U9449 ( .A(P3_P1_Flush), .B(_02597_), .S(_02604_), .Z(_02615_) );
  MUX2_X1 U9450 ( .A(P3_P1_More), .B(_02596_), .S(_02604_), .Z(_02614_) );
  MUX2_X1 U9451 ( .A(P3_P1_State2_PTR0), .B(_02609__PTR0), .S(_02604_), .Z(_02613__PTR0) );
  MUX2_X1 U9452 ( .A(P3_P1_State2_PTR1), .B(_02609__PTR1), .S(_02604_), .Z(_02613__PTR1) );
  MUX2_X1 U9453 ( .A(P3_P1_State2_PTR2), .B(_02609__PTR2), .S(_02604_), .Z(_02613__PTR2) );
  MUX2_X1 U9454 ( .A(P3_P1_State2_PTR3), .B(_02609__PTR3), .S(_02604_), .Z(_02613__PTR3) );
  MUX2_X1 U9455 ( .A(P3_EBX_PTR0), .B(_02594__PTR0), .S(_02604_), .Z(_02612__PTR0) );
  MUX2_X1 U9456 ( .A(P3_EBX_PTR1), .B(_02608__PTR1), .S(_02604_), .Z(_02612__PTR1) );
  MUX2_X1 U9457 ( .A(P3_EBX_PTR2), .B(_02608__PTR2), .S(_02604_), .Z(_02612__PTR2) );
  MUX2_X1 U9458 ( .A(P3_EBX_PTR3), .B(_02608__PTR3), .S(_02604_), .Z(_02612__PTR3) );
  MUX2_X1 U9459 ( .A(P3_EBX_PTR4), .B(_02608__PTR4), .S(_02604_), .Z(_02612__PTR4) );
  MUX2_X1 U9460 ( .A(P3_EBX_PTR5), .B(_02608__PTR5), .S(_02604_), .Z(_02612__PTR5) );
  MUX2_X1 U9461 ( .A(P3_EBX_PTR6), .B(_02608__PTR6), .S(_02604_), .Z(_02612__PTR6) );
  MUX2_X1 U9462 ( .A(P3_EBX_PTR7), .B(_02608__PTR7), .S(_02604_), .Z(_02612__PTR7) );
  MUX2_X1 U9463 ( .A(P3_EBX_PTR8), .B(_02608__PTR8), .S(_02604_), .Z(_02612__PTR8) );
  MUX2_X1 U9464 ( .A(P3_EBX_PTR9), .B(_02608__PTR9), .S(_02604_), .Z(_02612__PTR9) );
  MUX2_X1 U9465 ( .A(P3_EBX_PTR10), .B(_02608__PTR10), .S(_02604_), .Z(_02612__PTR10) );
  MUX2_X1 U9466 ( .A(P3_EBX_PTR11), .B(_02608__PTR11), .S(_02604_), .Z(_02612__PTR11) );
  MUX2_X1 U9467 ( .A(P3_EBX_PTR12), .B(_02608__PTR12), .S(_02604_), .Z(_02612__PTR12) );
  MUX2_X1 U9468 ( .A(P3_EBX_PTR13), .B(_02608__PTR13), .S(_02604_), .Z(_02612__PTR13) );
  MUX2_X1 U9469 ( .A(P3_EBX_PTR14), .B(_02608__PTR14), .S(_02604_), .Z(_02612__PTR14) );
  MUX2_X1 U9470 ( .A(P3_EBX_PTR15), .B(_02608__PTR15), .S(_02604_), .Z(_02612__PTR15) );
  MUX2_X1 U9471 ( .A(P3_EBX_PTR16), .B(_02608__PTR16), .S(_02604_), .Z(_02612__PTR16) );
  MUX2_X1 U9472 ( .A(P3_EBX_PTR17), .B(_02608__PTR17), .S(_02604_), .Z(_02612__PTR17) );
  MUX2_X1 U9473 ( .A(P3_EBX_PTR18), .B(_02608__PTR18), .S(_02604_), .Z(_02612__PTR18) );
  MUX2_X1 U9474 ( .A(P3_EBX_PTR19), .B(_02608__PTR19), .S(_02604_), .Z(_02612__PTR19) );
  MUX2_X1 U9475 ( .A(P3_EBX_PTR20), .B(_02608__PTR20), .S(_02604_), .Z(_02612__PTR20) );
  MUX2_X1 U9476 ( .A(P3_EBX_PTR21), .B(_02608__PTR21), .S(_02604_), .Z(_02612__PTR21) );
  MUX2_X1 U9477 ( .A(P3_EBX_PTR22), .B(_02608__PTR22), .S(_02604_), .Z(_02612__PTR22) );
  MUX2_X1 U9478 ( .A(P3_EBX_PTR23), .B(_02608__PTR23), .S(_02604_), .Z(_02612__PTR23) );
  MUX2_X1 U9479 ( .A(P3_EBX_PTR24), .B(_02608__PTR24), .S(_02604_), .Z(_02612__PTR24) );
  MUX2_X1 U9480 ( .A(P3_EBX_PTR25), .B(_02608__PTR25), .S(_02604_), .Z(_02612__PTR25) );
  MUX2_X1 U9481 ( .A(P3_EBX_PTR26), .B(_02608__PTR26), .S(_02604_), .Z(_02612__PTR26) );
  MUX2_X1 U9482 ( .A(P3_EBX_PTR27), .B(_02608__PTR27), .S(_02604_), .Z(_02612__PTR27) );
  MUX2_X1 U9483 ( .A(P3_EBX_PTR28), .B(_02608__PTR28), .S(_02604_), .Z(_02612__PTR28) );
  MUX2_X1 U9484 ( .A(P3_EBX_PTR29), .B(_02608__PTR29), .S(_02604_), .Z(_02612__PTR29) );
  MUX2_X1 U9485 ( .A(P3_EBX_PTR30), .B(_02608__PTR30), .S(_02604_), .Z(_02612__PTR30) );
  MUX2_X1 U9486 ( .A(P3_EBX_PTR31), .B(_02608__PTR31), .S(_02604_), .Z(_02612__PTR31) );
  MUX2_X1 U9487 ( .A(1'b1), .B(_02607_), .S(_02604_), .Z(_02611_) );
  MUX2_X1 U9488 ( .A(_02606__PTR0), .B(P3_P1_State2_PTR0), .S(P3_READY_n), .Z(_02609__PTR0) );
  MUX2_X1 U9489 ( .A(_02606__PTR1), .B(P3_P1_State2_PTR1), .S(P3_READY_n), .Z(_02609__PTR1) );
  MUX2_X1 U9490 ( .A(_02606__PTR2), .B(P3_P1_State2_PTR2), .S(P3_READY_n), .Z(_02609__PTR2) );
  MUX2_X1 U9491 ( .A(_02606__PTR3), .B(P3_P1_State2_PTR3), .S(P3_READY_n), .Z(_02609__PTR3) );
  MUX2_X1 U9492 ( .A(_02605__PTR1), .B(P3_EBX_PTR1), .S(P3_READY_n), .Z(_02608__PTR1) );
  MUX2_X1 U9493 ( .A(_02605__PTR2), .B(P3_EBX_PTR2), .S(P3_READY_n), .Z(_02608__PTR2) );
  MUX2_X1 U9494 ( .A(_02605__PTR3), .B(P3_EBX_PTR3), .S(P3_READY_n), .Z(_02608__PTR3) );
  MUX2_X1 U9495 ( .A(_02605__PTR4), .B(P3_EBX_PTR4), .S(P3_READY_n), .Z(_02608__PTR4) );
  MUX2_X1 U9496 ( .A(_02605__PTR5), .B(P3_EBX_PTR5), .S(P3_READY_n), .Z(_02608__PTR5) );
  MUX2_X1 U9497 ( .A(_02605__PTR6), .B(P3_EBX_PTR6), .S(P3_READY_n), .Z(_02608__PTR6) );
  MUX2_X1 U9498 ( .A(_02605__PTR7), .B(P3_EBX_PTR7), .S(P3_READY_n), .Z(_02608__PTR7) );
  MUX2_X1 U9499 ( .A(_02605__PTR8), .B(P3_EBX_PTR8), .S(P3_READY_n), .Z(_02608__PTR8) );
  MUX2_X1 U9500 ( .A(_02605__PTR9), .B(P3_EBX_PTR9), .S(P3_READY_n), .Z(_02608__PTR9) );
  MUX2_X1 U9501 ( .A(_02605__PTR10), .B(P3_EBX_PTR10), .S(P3_READY_n), .Z(_02608__PTR10) );
  MUX2_X1 U9502 ( .A(_02605__PTR11), .B(P3_EBX_PTR11), .S(P3_READY_n), .Z(_02608__PTR11) );
  MUX2_X1 U9503 ( .A(_02605__PTR12), .B(P3_EBX_PTR12), .S(P3_READY_n), .Z(_02608__PTR12) );
  MUX2_X1 U9504 ( .A(_02605__PTR13), .B(P3_EBX_PTR13), .S(P3_READY_n), .Z(_02608__PTR13) );
  MUX2_X1 U9505 ( .A(_02605__PTR14), .B(P3_EBX_PTR14), .S(P3_READY_n), .Z(_02608__PTR14) );
  MUX2_X1 U9506 ( .A(_02605__PTR15), .B(P3_EBX_PTR15), .S(P3_READY_n), .Z(_02608__PTR15) );
  MUX2_X1 U9507 ( .A(_02605__PTR16), .B(P3_EBX_PTR16), .S(P3_READY_n), .Z(_02608__PTR16) );
  MUX2_X1 U9508 ( .A(_02605__PTR17), .B(P3_EBX_PTR17), .S(P3_READY_n), .Z(_02608__PTR17) );
  MUX2_X1 U9509 ( .A(_02605__PTR18), .B(P3_EBX_PTR18), .S(P3_READY_n), .Z(_02608__PTR18) );
  MUX2_X1 U9510 ( .A(_02605__PTR19), .B(P3_EBX_PTR19), .S(P3_READY_n), .Z(_02608__PTR19) );
  MUX2_X1 U9511 ( .A(_02605__PTR20), .B(P3_EBX_PTR20), .S(P3_READY_n), .Z(_02608__PTR20) );
  MUX2_X1 U9512 ( .A(_02605__PTR21), .B(P3_EBX_PTR21), .S(P3_READY_n), .Z(_02608__PTR21) );
  MUX2_X1 U9513 ( .A(_02605__PTR22), .B(P3_EBX_PTR22), .S(P3_READY_n), .Z(_02608__PTR22) );
  MUX2_X1 U9514 ( .A(_02605__PTR23), .B(P3_EBX_PTR23), .S(P3_READY_n), .Z(_02608__PTR23) );
  MUX2_X1 U9515 ( .A(_02605__PTR24), .B(P3_EBX_PTR24), .S(P3_READY_n), .Z(_02608__PTR24) );
  MUX2_X1 U9516 ( .A(_02605__PTR25), .B(P3_EBX_PTR25), .S(P3_READY_n), .Z(_02608__PTR25) );
  MUX2_X1 U9517 ( .A(_02605__PTR26), .B(P3_EBX_PTR26), .S(P3_READY_n), .Z(_02608__PTR26) );
  MUX2_X1 U9518 ( .A(_02605__PTR27), .B(P3_EBX_PTR27), .S(P3_READY_n), .Z(_02608__PTR27) );
  MUX2_X1 U9519 ( .A(_02605__PTR28), .B(P3_EBX_PTR28), .S(P3_READY_n), .Z(_02608__PTR28) );
  MUX2_X1 U9520 ( .A(_02605__PTR29), .B(P3_EBX_PTR29), .S(P3_READY_n), .Z(_02608__PTR29) );
  MUX2_X1 U9521 ( .A(_02605__PTR30), .B(P3_EBX_PTR30), .S(P3_READY_n), .Z(_02608__PTR30) );
  MUX2_X1 U9522 ( .A(_02605__PTR31), .B(P3_EBX_PTR31), .S(P3_READY_n), .Z(_02608__PTR31) );
  MUX2_X1 U9523 ( .A(_02475__PTR9), .B(1'b1), .S(P3_READY_n), .Z(_02607_) );
  MUX2_X1 U9524 ( .A(1'b0), .B(P3_P1_State2_PTR0), .S(P3_StateBS16), .Z(_02606__PTR0) );
  MUX2_X1 U9525 ( .A(1'b1), .B(P3_P1_State2_PTR1), .S(P3_StateBS16), .Z(_02606__PTR1) );
  MUX2_X1 U9526 ( .A(1'b1), .B(P3_P1_State2_PTR2), .S(P3_StateBS16), .Z(_02606__PTR2) );
  MUX2_X1 U9527 ( .A(1'b0), .B(P3_P1_State2_PTR3), .S(P3_StateBS16), .Z(_02606__PTR3) );
  MUX2_X1 U9528 ( .A(_02463__PTR7), .B(P3_EBX_PTR1), .S(P3_StateBS16), .Z(_02605__PTR1) );
  MUX2_X1 U9529 ( .A(_03312__PTR1), .B(P3_EBX_PTR2), .S(P3_StateBS16), .Z(_02605__PTR2) );
  MUX2_X1 U9530 ( .A(_03312__PTR2), .B(P3_EBX_PTR3), .S(P3_StateBS16), .Z(_02605__PTR3) );
  MUX2_X1 U9531 ( .A(_03312__PTR3), .B(P3_EBX_PTR4), .S(P3_StateBS16), .Z(_02605__PTR4) );
  MUX2_X1 U9532 ( .A(_03312__PTR4), .B(P3_EBX_PTR5), .S(P3_StateBS16), .Z(_02605__PTR5) );
  MUX2_X1 U9533 ( .A(_03312__PTR5), .B(P3_EBX_PTR6), .S(P3_StateBS16), .Z(_02605__PTR6) );
  MUX2_X1 U9534 ( .A(_03312__PTR6), .B(P3_EBX_PTR7), .S(P3_StateBS16), .Z(_02605__PTR7) );
  MUX2_X1 U9535 ( .A(_03312__PTR7), .B(P3_EBX_PTR8), .S(P3_StateBS16), .Z(_02605__PTR8) );
  MUX2_X1 U9536 ( .A(_03312__PTR8), .B(P3_EBX_PTR9), .S(P3_StateBS16), .Z(_02605__PTR9) );
  MUX2_X1 U9537 ( .A(_03312__PTR9), .B(P3_EBX_PTR10), .S(P3_StateBS16), .Z(_02605__PTR10) );
  MUX2_X1 U9538 ( .A(_03312__PTR10), .B(P3_EBX_PTR11), .S(P3_StateBS16), .Z(_02605__PTR11) );
  MUX2_X1 U9539 ( .A(_03312__PTR11), .B(P3_EBX_PTR12), .S(P3_StateBS16), .Z(_02605__PTR12) );
  MUX2_X1 U9540 ( .A(_03312__PTR12), .B(P3_EBX_PTR13), .S(P3_StateBS16), .Z(_02605__PTR13) );
  MUX2_X1 U9541 ( .A(_03312__PTR13), .B(P3_EBX_PTR14), .S(P3_StateBS16), .Z(_02605__PTR14) );
  MUX2_X1 U9542 ( .A(_03312__PTR14), .B(P3_EBX_PTR15), .S(P3_StateBS16), .Z(_02605__PTR15) );
  MUX2_X1 U9543 ( .A(_03312__PTR15), .B(P3_EBX_PTR16), .S(P3_StateBS16), .Z(_02605__PTR16) );
  MUX2_X1 U9544 ( .A(_03312__PTR16), .B(P3_EBX_PTR17), .S(P3_StateBS16), .Z(_02605__PTR17) );
  MUX2_X1 U9545 ( .A(_03312__PTR17), .B(P3_EBX_PTR18), .S(P3_StateBS16), .Z(_02605__PTR18) );
  MUX2_X1 U9546 ( .A(_03312__PTR18), .B(P3_EBX_PTR19), .S(P3_StateBS16), .Z(_02605__PTR19) );
  MUX2_X1 U9547 ( .A(_03312__PTR19), .B(P3_EBX_PTR20), .S(P3_StateBS16), .Z(_02605__PTR20) );
  MUX2_X1 U9548 ( .A(_03312__PTR20), .B(P3_EBX_PTR21), .S(P3_StateBS16), .Z(_02605__PTR21) );
  MUX2_X1 U9549 ( .A(_03312__PTR21), .B(P3_EBX_PTR22), .S(P3_StateBS16), .Z(_02605__PTR22) );
  MUX2_X1 U9550 ( .A(_03312__PTR22), .B(P3_EBX_PTR23), .S(P3_StateBS16), .Z(_02605__PTR23) );
  MUX2_X1 U9551 ( .A(_03312__PTR23), .B(P3_EBX_PTR24), .S(P3_StateBS16), .Z(_02605__PTR24) );
  MUX2_X1 U9552 ( .A(_03312__PTR24), .B(P3_EBX_PTR25), .S(P3_StateBS16), .Z(_02605__PTR25) );
  MUX2_X1 U9553 ( .A(_03312__PTR25), .B(P3_EBX_PTR26), .S(P3_StateBS16), .Z(_02605__PTR26) );
  MUX2_X1 U9554 ( .A(_03312__PTR26), .B(P3_EBX_PTR27), .S(P3_StateBS16), .Z(_02605__PTR27) );
  MUX2_X1 U9555 ( .A(_03312__PTR27), .B(P3_EBX_PTR28), .S(P3_StateBS16), .Z(_02605__PTR28) );
  MUX2_X1 U9556 ( .A(_03312__PTR28), .B(P3_EBX_PTR29), .S(P3_StateBS16), .Z(_02605__PTR29) );
  MUX2_X1 U9557 ( .A(_03312__PTR29), .B(P3_EBX_PTR30), .S(P3_StateBS16), .Z(_02605__PTR30) );
  MUX2_X1 U9558 ( .A(_03312__PTR30), .B(P3_EBX_PTR31), .S(P3_StateBS16), .Z(_02605__PTR31) );
  MUX2_X1 U9559 ( .A(_03308__PTR3), .B(P3_P1_InstQueueRd_Addr_PTR4), .S(P3_READY_n), .Z(_02624__PTR4) );
  MUX2_X1 U9560 ( .A(_02471__PTR4), .B(P3_P1_InstQueueRd_Addr_PTR1), .S(P3_READY_n), .Z(_02599__PTR1) );
  MUX2_X1 U9561 ( .A(_02471__PTR5), .B(P3_P1_InstQueueRd_Addr_PTR2), .S(P3_READY_n), .Z(_02599__PTR2) );
  MUX2_X1 U9562 ( .A(_02471__PTR6), .B(P3_P1_InstQueueRd_Addr_PTR3), .S(P3_READY_n), .Z(_02599__PTR3) );
  MUX2_X1 U9563 ( .A(1'b0), .B(P3_P1_InstQueueRd_Addr_PTR4), .S(P3_READY_n), .Z(_02599__PTR4) );
  MUX2_X1 U9564 ( .A(P3_P1_lWord_PTR0), .B(P3_EAX_PTR0), .S(_02585_), .Z(_02689__PTR16) );
  MUX2_X1 U9565 ( .A(P3_P1_lWord_PTR1), .B(P3_EAX_PTR1), .S(_02585_), .Z(_02689__PTR17) );
  MUX2_X1 U9566 ( .A(P3_P1_lWord_PTR2), .B(P3_EAX_PTR2), .S(_02585_), .Z(_02689__PTR18) );
  MUX2_X1 U9567 ( .A(P3_P1_lWord_PTR3), .B(P3_EAX_PTR3), .S(_02585_), .Z(_02689__PTR19) );
  MUX2_X1 U9568 ( .A(P3_P1_lWord_PTR4), .B(P3_EAX_PTR4), .S(_02585_), .Z(_02689__PTR20) );
  MUX2_X1 U9569 ( .A(P3_P1_lWord_PTR5), .B(P3_EAX_PTR5), .S(_02585_), .Z(_02689__PTR21) );
  MUX2_X1 U9570 ( .A(P3_P1_lWord_PTR6), .B(P3_EAX_PTR6), .S(_02585_), .Z(_02689__PTR22) );
  MUX2_X1 U9571 ( .A(P3_P1_lWord_PTR7), .B(P3_EAX_PTR7), .S(_02585_), .Z(_02689__PTR23) );
  MUX2_X1 U9572 ( .A(P3_P1_lWord_PTR8), .B(P3_EAX_PTR8), .S(_02585_), .Z(_02689__PTR24) );
  MUX2_X1 U9573 ( .A(P3_P1_lWord_PTR9), .B(P3_EAX_PTR9), .S(_02585_), .Z(_02689__PTR25) );
  MUX2_X1 U9574 ( .A(P3_P1_lWord_PTR10), .B(P3_EAX_PTR10), .S(_02585_), .Z(_02689__PTR26) );
  MUX2_X1 U9575 ( .A(P3_P1_lWord_PTR11), .B(P3_EAX_PTR11), .S(_02585_), .Z(_02689__PTR27) );
  MUX2_X1 U9576 ( .A(P3_P1_lWord_PTR12), .B(P3_EAX_PTR12), .S(_02585_), .Z(_02689__PTR28) );
  MUX2_X1 U9577 ( .A(P3_P1_lWord_PTR13), .B(P3_EAX_PTR13), .S(_02585_), .Z(_02689__PTR29) );
  MUX2_X1 U9578 ( .A(P3_P1_lWord_PTR14), .B(P3_EAX_PTR14), .S(_02585_), .Z(_02689__PTR30) );
  MUX2_X1 U9579 ( .A(P3_P1_lWord_PTR15), .B(P3_EAX_PTR15), .S(_02585_), .Z(_02689__PTR31) );
  MUX2_X1 U9580 ( .A(P3_P1_lWord_PTR0), .B(_02593__PTR0), .S(_02585_), .Z(_02689__PTR32) );
  MUX2_X1 U9581 ( .A(P3_P1_lWord_PTR1), .B(_02593__PTR1), .S(_02585_), .Z(_02689__PTR33) );
  MUX2_X1 U9582 ( .A(P3_P1_lWord_PTR2), .B(_02593__PTR2), .S(_02585_), .Z(_02689__PTR34) );
  MUX2_X1 U9583 ( .A(P3_P1_lWord_PTR3), .B(_02593__PTR3), .S(_02585_), .Z(_02689__PTR35) );
  MUX2_X1 U9584 ( .A(P3_P1_lWord_PTR4), .B(_02593__PTR4), .S(_02585_), .Z(_02689__PTR36) );
  MUX2_X1 U9585 ( .A(P3_P1_lWord_PTR5), .B(_02593__PTR5), .S(_02585_), .Z(_02689__PTR37) );
  MUX2_X1 U9586 ( .A(P3_P1_lWord_PTR6), .B(_02593__PTR6), .S(_02585_), .Z(_02689__PTR38) );
  MUX2_X1 U9587 ( .A(P3_P1_lWord_PTR7), .B(_02593__PTR7), .S(_02585_), .Z(_02689__PTR39) );
  MUX2_X1 U9588 ( .A(P3_P1_lWord_PTR8), .B(_02593__PTR8), .S(_02585_), .Z(_02689__PTR40) );
  MUX2_X1 U9589 ( .A(P3_P1_lWord_PTR9), .B(_02593__PTR9), .S(_02585_), .Z(_02689__PTR41) );
  MUX2_X1 U9590 ( .A(P3_P1_lWord_PTR10), .B(_02593__PTR10), .S(_02585_), .Z(_02689__PTR42) );
  MUX2_X1 U9591 ( .A(P3_P1_lWord_PTR11), .B(_02593__PTR11), .S(_02585_), .Z(_02689__PTR43) );
  MUX2_X1 U9592 ( .A(P3_P1_lWord_PTR12), .B(_02593__PTR12), .S(_02585_), .Z(_02689__PTR44) );
  MUX2_X1 U9593 ( .A(P3_P1_lWord_PTR13), .B(_02593__PTR13), .S(_02585_), .Z(_02689__PTR45) );
  MUX2_X1 U9594 ( .A(P3_P1_lWord_PTR14), .B(_02593__PTR14), .S(_02585_), .Z(_02689__PTR46) );
  MUX2_X1 U9595 ( .A(P3_P1_lWord_PTR15), .B(_02593__PTR15), .S(_02585_), .Z(_02689__PTR47) );
  MUX2_X1 U9596 ( .A(1'b0), .B(_02597_), .S(_02585_), .Z(_02435__PTR1) );
  MUX2_X1 U9597 ( .A(1'b1), .B(_02596_), .S(_02585_), .Z(_02439__PTR1) );
  MUX2_X1 U9598 ( .A(buf2_PTR16), .B(P3_EAX_PTR16), .S(P3_READY_n), .Z(_02623__PTR16) );
  MUX2_X1 U9599 ( .A(buf2_PTR17), .B(P3_EAX_PTR17), .S(P3_READY_n), .Z(_02623__PTR17) );
  MUX2_X1 U9600 ( .A(buf2_PTR18), .B(P3_EAX_PTR18), .S(P3_READY_n), .Z(_02623__PTR18) );
  MUX2_X1 U9601 ( .A(buf2_PTR19), .B(P3_EAX_PTR19), .S(P3_READY_n), .Z(_02623__PTR19) );
  MUX2_X1 U9602 ( .A(buf2_PTR20), .B(P3_EAX_PTR20), .S(P3_READY_n), .Z(_02623__PTR20) );
  MUX2_X1 U9603 ( .A(buf2_PTR21), .B(P3_EAX_PTR21), .S(P3_READY_n), .Z(_02623__PTR21) );
  MUX2_X1 U9604 ( .A(buf2_PTR22), .B(P3_EAX_PTR22), .S(P3_READY_n), .Z(_02623__PTR22) );
  MUX2_X1 U9605 ( .A(buf2_PTR23), .B(P3_EAX_PTR23), .S(P3_READY_n), .Z(_02623__PTR23) );
  MUX2_X1 U9606 ( .A(buf2_PTR24), .B(P3_EAX_PTR24), .S(P3_READY_n), .Z(_02623__PTR24) );
  MUX2_X1 U9607 ( .A(buf2_PTR25), .B(P3_EAX_PTR25), .S(P3_READY_n), .Z(_02623__PTR25) );
  MUX2_X1 U9608 ( .A(buf2_PTR26), .B(P3_EAX_PTR26), .S(P3_READY_n), .Z(_02623__PTR26) );
  MUX2_X1 U9609 ( .A(buf2_PTR27), .B(P3_EAX_PTR27), .S(P3_READY_n), .Z(_02623__PTR27) );
  MUX2_X1 U9610 ( .A(buf2_PTR28), .B(P3_EAX_PTR28), .S(P3_READY_n), .Z(_02623__PTR28) );
  MUX2_X1 U9611 ( .A(buf2_PTR29), .B(P3_EAX_PTR29), .S(P3_READY_n), .Z(_02623__PTR29) );
  MUX2_X1 U9612 ( .A(buf2_PTR30), .B(P3_EAX_PTR30), .S(P3_READY_n), .Z(_02623__PTR30) );
  MUX2_X1 U9613 ( .A(buf2_PTR31), .B(P3_EAX_PTR31), .S(P3_READY_n), .Z(_02623__PTR31) );
  MUX2_X1 U9614 ( .A(buf2_PTR0), .B(P3_EAX_PTR0), .S(P3_READY_n), .Z(_02595__PTR0) );
  MUX2_X1 U9615 ( .A(buf2_PTR1), .B(P3_EAX_PTR1), .S(P3_READY_n), .Z(_02595__PTR1) );
  MUX2_X1 U9616 ( .A(buf2_PTR2), .B(P3_EAX_PTR2), .S(P3_READY_n), .Z(_02595__PTR2) );
  MUX2_X1 U9617 ( .A(buf2_PTR3), .B(P3_EAX_PTR3), .S(P3_READY_n), .Z(_02595__PTR3) );
  MUX2_X1 U9618 ( .A(buf2_PTR4), .B(P3_EAX_PTR4), .S(P3_READY_n), .Z(_02595__PTR4) );
  MUX2_X1 U9619 ( .A(buf2_PTR5), .B(P3_EAX_PTR5), .S(P3_READY_n), .Z(_02595__PTR5) );
  MUX2_X1 U9620 ( .A(buf2_PTR6), .B(P3_EAX_PTR6), .S(P3_READY_n), .Z(_02595__PTR6) );
  MUX2_X1 U9621 ( .A(buf2_PTR7), .B(P3_EAX_PTR7), .S(P3_READY_n), .Z(_02595__PTR7) );
  MUX2_X1 U9622 ( .A(buf2_PTR8), .B(P3_EAX_PTR8), .S(P3_READY_n), .Z(_02595__PTR8) );
  MUX2_X1 U9623 ( .A(buf2_PTR9), .B(P3_EAX_PTR9), .S(P3_READY_n), .Z(_02595__PTR9) );
  MUX2_X1 U9624 ( .A(buf2_PTR10), .B(P3_EAX_PTR10), .S(P3_READY_n), .Z(_02595__PTR10) );
  MUX2_X1 U9625 ( .A(buf2_PTR11), .B(P3_EAX_PTR11), .S(P3_READY_n), .Z(_02595__PTR11) );
  MUX2_X1 U9626 ( .A(buf2_PTR12), .B(P3_EAX_PTR12), .S(P3_READY_n), .Z(_02595__PTR12) );
  MUX2_X1 U9627 ( .A(buf2_PTR13), .B(P3_EAX_PTR13), .S(P3_READY_n), .Z(_02595__PTR13) );
  MUX2_X1 U9628 ( .A(buf2_PTR14), .B(P3_EAX_PTR14), .S(P3_READY_n), .Z(_02595__PTR14) );
  MUX2_X1 U9629 ( .A(buf2_PTR15), .B(P3_EAX_PTR15), .S(P3_READY_n), .Z(_02595__PTR15) );
  MUX2_X1 U9630 ( .A(buf2_PTR0), .B(P3_EAX_PTR16), .S(P3_READY_n), .Z(_02595__PTR16) );
  MUX2_X1 U9631 ( .A(buf2_PTR1), .B(P3_EAX_PTR17), .S(P3_READY_n), .Z(_02595__PTR17) );
  MUX2_X1 U9632 ( .A(buf2_PTR2), .B(P3_EAX_PTR18), .S(P3_READY_n), .Z(_02595__PTR18) );
  MUX2_X1 U9633 ( .A(buf2_PTR3), .B(P3_EAX_PTR19), .S(P3_READY_n), .Z(_02595__PTR19) );
  MUX2_X1 U9634 ( .A(buf2_PTR4), .B(P3_EAX_PTR20), .S(P3_READY_n), .Z(_02595__PTR20) );
  MUX2_X1 U9635 ( .A(buf2_PTR5), .B(P3_EAX_PTR21), .S(P3_READY_n), .Z(_02595__PTR21) );
  MUX2_X1 U9636 ( .A(buf2_PTR6), .B(P3_EAX_PTR22), .S(P3_READY_n), .Z(_02595__PTR22) );
  MUX2_X1 U9637 ( .A(buf2_PTR7), .B(P3_EAX_PTR23), .S(P3_READY_n), .Z(_02595__PTR23) );
  MUX2_X1 U9638 ( .A(buf2_PTR8), .B(P3_EAX_PTR24), .S(P3_READY_n), .Z(_02595__PTR24) );
  MUX2_X1 U9639 ( .A(buf2_PTR9), .B(P3_EAX_PTR25), .S(P3_READY_n), .Z(_02595__PTR25) );
  MUX2_X1 U9640 ( .A(buf2_PTR10), .B(P3_EAX_PTR26), .S(P3_READY_n), .Z(_02595__PTR26) );
  MUX2_X1 U9641 ( .A(buf2_PTR11), .B(P3_EAX_PTR27), .S(P3_READY_n), .Z(_02595__PTR27) );
  MUX2_X1 U9642 ( .A(buf2_PTR12), .B(P3_EAX_PTR28), .S(P3_READY_n), .Z(_02595__PTR28) );
  MUX2_X1 U9643 ( .A(buf2_PTR13), .B(P3_EAX_PTR29), .S(P3_READY_n), .Z(_02595__PTR29) );
  MUX2_X1 U9644 ( .A(buf2_PTR14), .B(P3_EAX_PTR30), .S(P3_READY_n), .Z(_02595__PTR30) );
  MUX2_X1 U9645 ( .A(1'b0), .B(P3_EAX_PTR31), .S(P3_READY_n), .Z(_02595__PTR31) );
  MUX2_X1 U9646 ( .A(P3_P1_uWord_PTR0), .B(_03315__PTR0), .S(_02585_), .Z(_02685__PTR15) );
  MUX2_X1 U9647 ( .A(P3_P1_uWord_PTR1), .B(_03316__PTR1), .S(_02585_), .Z(_02685__PTR16) );
  MUX2_X1 U9648 ( .A(P3_P1_uWord_PTR2), .B(_03316__PTR2), .S(_02585_), .Z(_02685__PTR17) );
  MUX2_X1 U9649 ( .A(P3_P1_uWord_PTR3), .B(_03316__PTR3), .S(_02585_), .Z(_02685__PTR18) );
  MUX2_X1 U9650 ( .A(P3_P1_uWord_PTR4), .B(_03316__PTR4), .S(_02585_), .Z(_02685__PTR19) );
  MUX2_X1 U9651 ( .A(P3_P1_uWord_PTR5), .B(_03316__PTR5), .S(_02585_), .Z(_02685__PTR20) );
  MUX2_X1 U9652 ( .A(P3_P1_uWord_PTR6), .B(_03316__PTR6), .S(_02585_), .Z(_02685__PTR21) );
  MUX2_X1 U9653 ( .A(P3_P1_uWord_PTR7), .B(_03316__PTR7), .S(_02585_), .Z(_02685__PTR22) );
  MUX2_X1 U9654 ( .A(P3_P1_uWord_PTR8), .B(_03316__PTR8), .S(_02585_), .Z(_02685__PTR23) );
  MUX2_X1 U9655 ( .A(P3_P1_uWord_PTR9), .B(_03316__PTR9), .S(_02585_), .Z(_02685__PTR24) );
  MUX2_X1 U9656 ( .A(P3_P1_uWord_PTR10), .B(_03316__PTR10), .S(_02585_), .Z(_02685__PTR25) );
  MUX2_X1 U9657 ( .A(P3_P1_uWord_PTR11), .B(_03316__PTR11), .S(_02585_), .Z(_02685__PTR26) );
  MUX2_X1 U9658 ( .A(P3_P1_uWord_PTR12), .B(_03316__PTR12), .S(_02585_), .Z(_02685__PTR27) );
  MUX2_X1 U9659 ( .A(P3_P1_uWord_PTR13), .B(_03316__PTR13), .S(_02585_), .Z(_02685__PTR28) );
  MUX2_X1 U9660 ( .A(P3_P1_uWord_PTR14), .B(_03316__PTR14), .S(_02585_), .Z(_02685__PTR29) );
  MUX2_X1 U9661 ( .A(P3_P1_uWord_PTR0), .B(_02592__PTR0), .S(_02585_), .Z(_02685__PTR30) );
  MUX2_X1 U9662 ( .A(P3_P1_uWord_PTR1), .B(_02592__PTR1), .S(_02585_), .Z(_02685__PTR31) );
  MUX2_X1 U9663 ( .A(P3_P1_uWord_PTR2), .B(_02592__PTR2), .S(_02585_), .Z(_02685__PTR32) );
  MUX2_X1 U9664 ( .A(P3_P1_uWord_PTR3), .B(_02592__PTR3), .S(_02585_), .Z(_02685__PTR33) );
  MUX2_X1 U9665 ( .A(P3_P1_uWord_PTR4), .B(_02592__PTR4), .S(_02585_), .Z(_02685__PTR34) );
  MUX2_X1 U9666 ( .A(P3_P1_uWord_PTR5), .B(_02592__PTR5), .S(_02585_), .Z(_02685__PTR35) );
  MUX2_X1 U9667 ( .A(P3_P1_uWord_PTR6), .B(_02592__PTR6), .S(_02585_), .Z(_02685__PTR36) );
  MUX2_X1 U9668 ( .A(P3_P1_uWord_PTR7), .B(_02592__PTR7), .S(_02585_), .Z(_02685__PTR37) );
  MUX2_X1 U9669 ( .A(P3_P1_uWord_PTR8), .B(_02592__PTR8), .S(_02585_), .Z(_02685__PTR38) );
  MUX2_X1 U9670 ( .A(P3_P1_uWord_PTR9), .B(_02592__PTR9), .S(_02585_), .Z(_02685__PTR39) );
  MUX2_X1 U9671 ( .A(P3_P1_uWord_PTR10), .B(_02592__PTR10), .S(_02585_), .Z(_02685__PTR40) );
  MUX2_X1 U9672 ( .A(P3_P1_uWord_PTR11), .B(_02592__PTR11), .S(_02585_), .Z(_02685__PTR41) );
  MUX2_X1 U9673 ( .A(P3_P1_uWord_PTR12), .B(_02592__PTR12), .S(_02585_), .Z(_02685__PTR42) );
  MUX2_X1 U9674 ( .A(P3_P1_uWord_PTR13), .B(_02592__PTR13), .S(_02585_), .Z(_02685__PTR43) );
  MUX2_X1 U9675 ( .A(P3_P1_uWord_PTR14), .B(_02592__PTR14), .S(_02585_), .Z(_02685__PTR44) );
  MUX2_X1 U9676 ( .A(P3_CodeFetch), .B(1'b0), .S(_02585_), .Z(_02454__PTR0) );
  MUX2_X1 U9677 ( .A(P3_MemoryFetch), .B(1'b1), .S(_02585_), .Z(_02450__PTR1) );
  MUX2_X1 U9678 ( .A(P3_ReadRequest), .B(1'b1), .S(_02585_), .Z(_02447__PTR1) );
  MUX2_X1 U9679 ( .A(P3_RequestPending), .B(P3_READY_n), .S(_02585_), .Z(_02443__PTR1) );
  MUX2_X1 U9680 ( .A(P3_P1_InstQueueRd_Addr_PTR4), .B(_02624__PTR4), .S(_02585_), .Z(_02666__PTR19) );
  MUX2_X1 U9681 ( .A(P3_P1_InstQueueRd_Addr_PTR1), .B(_02617__PTR1), .S(_02585_), .Z(_02666__PTR11) );
  MUX2_X1 U9682 ( .A(P3_P1_InstQueueRd_Addr_PTR2), .B(_02617__PTR2), .S(_02585_), .Z(_02666__PTR12) );
  MUX2_X1 U9683 ( .A(P3_P1_InstQueueRd_Addr_PTR3), .B(_02617__PTR3), .S(_02585_), .Z(_02666__PTR13) );
  MUX2_X1 U9684 ( .A(P3_P1_InstQueueRd_Addr_PTR4), .B(_02617__PTR4), .S(_02585_), .Z(_02666__PTR14) );
  MUX2_X1 U9685 ( .A(P3_P1_InstQueueRd_Addr_PTR1), .B(_02599__PTR1), .S(_02585_), .Z(_02666__PTR21) );
  MUX2_X1 U9686 ( .A(P3_P1_InstQueueRd_Addr_PTR2), .B(_02599__PTR2), .S(_02585_), .Z(_02666__PTR22) );
  MUX2_X1 U9687 ( .A(P3_P1_InstQueueRd_Addr_PTR3), .B(_02599__PTR3), .S(_02585_), .Z(_02666__PTR23) );
  MUX2_X1 U9688 ( .A(P3_P1_InstQueueRd_Addr_PTR4), .B(_02599__PTR4), .S(_02585_), .Z(_02666__PTR24) );
  MUX2_X1 U9689 ( .A(_02662__PTR33), .B(P3_P1_InstAddrPointer_PTR1), .S(P3_READY_n), .Z(_02598__PTR1) );
  MUX2_X1 U9690 ( .A(_02662__PTR34), .B(P3_P1_InstAddrPointer_PTR2), .S(P3_READY_n), .Z(_02598__PTR2) );
  MUX2_X1 U9691 ( .A(_02662__PTR35), .B(P3_P1_InstAddrPointer_PTR3), .S(P3_READY_n), .Z(_02598__PTR3) );
  MUX2_X1 U9692 ( .A(_02662__PTR36), .B(P3_P1_InstAddrPointer_PTR4), .S(P3_READY_n), .Z(_02598__PTR4) );
  MUX2_X1 U9693 ( .A(_02662__PTR37), .B(P3_P1_InstAddrPointer_PTR5), .S(P3_READY_n), .Z(_02598__PTR5) );
  MUX2_X1 U9694 ( .A(_02662__PTR38), .B(P3_P1_InstAddrPointer_PTR6), .S(P3_READY_n), .Z(_02598__PTR6) );
  MUX2_X1 U9695 ( .A(_02662__PTR39), .B(P3_P1_InstAddrPointer_PTR7), .S(P3_READY_n), .Z(_02598__PTR7) );
  MUX2_X1 U9696 ( .A(_02662__PTR40), .B(P3_P1_InstAddrPointer_PTR8), .S(P3_READY_n), .Z(_02598__PTR8) );
  MUX2_X1 U9697 ( .A(_02662__PTR41), .B(P3_P1_InstAddrPointer_PTR9), .S(P3_READY_n), .Z(_02598__PTR9) );
  MUX2_X1 U9698 ( .A(_02662__PTR42), .B(P3_P1_InstAddrPointer_PTR10), .S(P3_READY_n), .Z(_02598__PTR10) );
  MUX2_X1 U9699 ( .A(_02662__PTR43), .B(P3_P1_InstAddrPointer_PTR11), .S(P3_READY_n), .Z(_02598__PTR11) );
  MUX2_X1 U9700 ( .A(_02662__PTR44), .B(P3_P1_InstAddrPointer_PTR12), .S(P3_READY_n), .Z(_02598__PTR12) );
  MUX2_X1 U9701 ( .A(_02662__PTR45), .B(P3_P1_InstAddrPointer_PTR13), .S(P3_READY_n), .Z(_02598__PTR13) );
  MUX2_X1 U9702 ( .A(_02662__PTR46), .B(P3_P1_InstAddrPointer_PTR14), .S(P3_READY_n), .Z(_02598__PTR14) );
  MUX2_X1 U9703 ( .A(_02662__PTR47), .B(P3_P1_InstAddrPointer_PTR15), .S(P3_READY_n), .Z(_02598__PTR15) );
  MUX2_X1 U9704 ( .A(_02662__PTR48), .B(P3_P1_InstAddrPointer_PTR16), .S(P3_READY_n), .Z(_02598__PTR16) );
  MUX2_X1 U9705 ( .A(_02662__PTR49), .B(P3_P1_InstAddrPointer_PTR17), .S(P3_READY_n), .Z(_02598__PTR17) );
  MUX2_X1 U9706 ( .A(_02662__PTR50), .B(P3_P1_InstAddrPointer_PTR18), .S(P3_READY_n), .Z(_02598__PTR18) );
  MUX2_X1 U9707 ( .A(_02662__PTR51), .B(P3_P1_InstAddrPointer_PTR19), .S(P3_READY_n), .Z(_02598__PTR19) );
  MUX2_X1 U9708 ( .A(_02662__PTR52), .B(P3_P1_InstAddrPointer_PTR20), .S(P3_READY_n), .Z(_02598__PTR20) );
  MUX2_X1 U9709 ( .A(_02662__PTR53), .B(P3_P1_InstAddrPointer_PTR21), .S(P3_READY_n), .Z(_02598__PTR21) );
  MUX2_X1 U9710 ( .A(_02662__PTR54), .B(P3_P1_InstAddrPointer_PTR22), .S(P3_READY_n), .Z(_02598__PTR22) );
  MUX2_X1 U9711 ( .A(_02662__PTR55), .B(P3_P1_InstAddrPointer_PTR23), .S(P3_READY_n), .Z(_02598__PTR23) );
  MUX2_X1 U9712 ( .A(_02662__PTR56), .B(P3_P1_InstAddrPointer_PTR24), .S(P3_READY_n), .Z(_02598__PTR24) );
  MUX2_X1 U9713 ( .A(_02662__PTR57), .B(P3_P1_InstAddrPointer_PTR25), .S(P3_READY_n), .Z(_02598__PTR25) );
  MUX2_X1 U9714 ( .A(_02662__PTR58), .B(P3_P1_InstAddrPointer_PTR26), .S(P3_READY_n), .Z(_02598__PTR26) );
  MUX2_X1 U9715 ( .A(_02662__PTR59), .B(P3_P1_InstAddrPointer_PTR27), .S(P3_READY_n), .Z(_02598__PTR27) );
  MUX2_X1 U9716 ( .A(_02662__PTR60), .B(P3_P1_InstAddrPointer_PTR28), .S(P3_READY_n), .Z(_02598__PTR28) );
  MUX2_X1 U9717 ( .A(_02662__PTR61), .B(P3_P1_InstAddrPointer_PTR29), .S(P3_READY_n), .Z(_02598__PTR29) );
  MUX2_X1 U9718 ( .A(_02662__PTR62), .B(P3_P1_InstAddrPointer_PTR30), .S(P3_READY_n), .Z(_02598__PTR30) );
  MUX2_X1 U9719 ( .A(_02662__PTR63), .B(P3_P1_InstAddrPointer_PTR31), .S(P3_READY_n), .Z(_02598__PTR31) );
  MUX2_X1 U9720 ( .A(1'b0), .B(P3_P1_Flush), .S(P3_READY_n), .Z(_02597_) );
  MUX2_X1 U9721 ( .A(1'b0), .B(P3_P1_More), .S(P3_READY_n), .Z(_02596_) );
  MUX2_X1 U9722 ( .A(_02589__PTR0), .B(P3_EBX_PTR0), .S(P3_READY_n), .Z(_02594__PTR0) );
  MUX2_X1 U9723 ( .A(_02589__PTR1), .B(_02588__PTR1), .S(P3_READY_n), .Z(_02594__PTR1) );
  MUX2_X1 U9724 ( .A(_02589__PTR2), .B(_02588__PTR2), .S(P3_READY_n), .Z(_02594__PTR2) );
  MUX2_X1 U9725 ( .A(_02589__PTR3), .B(_02588__PTR3), .S(P3_READY_n), .Z(_02594__PTR3) );
  MUX2_X1 U9726 ( .A(_02589__PTR4), .B(_02588__PTR4), .S(P3_READY_n), .Z(_02594__PTR4) );
  MUX2_X1 U9727 ( .A(_02589__PTR5), .B(_02588__PTR5), .S(P3_READY_n), .Z(_02594__PTR5) );
  MUX2_X1 U9728 ( .A(_02589__PTR6), .B(_02588__PTR6), .S(P3_READY_n), .Z(_02594__PTR6) );
  MUX2_X1 U9729 ( .A(_02589__PTR7), .B(_02588__PTR7), .S(P3_READY_n), .Z(_02594__PTR7) );
  MUX2_X1 U9730 ( .A(_02589__PTR8), .B(_02588__PTR8), .S(P3_READY_n), .Z(_02594__PTR8) );
  MUX2_X1 U9731 ( .A(_02589__PTR9), .B(_02588__PTR9), .S(P3_READY_n), .Z(_02594__PTR9) );
  MUX2_X1 U9732 ( .A(_02589__PTR10), .B(_02588__PTR10), .S(P3_READY_n), .Z(_02594__PTR10) );
  MUX2_X1 U9733 ( .A(_02589__PTR11), .B(_02588__PTR11), .S(P3_READY_n), .Z(_02594__PTR11) );
  MUX2_X1 U9734 ( .A(_02589__PTR12), .B(_02588__PTR12), .S(P3_READY_n), .Z(_02594__PTR12) );
  MUX2_X1 U9735 ( .A(_02589__PTR13), .B(_02588__PTR13), .S(P3_READY_n), .Z(_02594__PTR13) );
  MUX2_X1 U9736 ( .A(_02589__PTR14), .B(_02588__PTR14), .S(P3_READY_n), .Z(_02594__PTR14) );
  MUX2_X1 U9737 ( .A(_02589__PTR15), .B(_02588__PTR15), .S(P3_READY_n), .Z(_02594__PTR15) );
  MUX2_X1 U9738 ( .A(_02589__PTR16), .B(_02588__PTR16), .S(P3_READY_n), .Z(_02594__PTR16) );
  MUX2_X1 U9739 ( .A(_02589__PTR17), .B(_02588__PTR17), .S(P3_READY_n), .Z(_02594__PTR17) );
  MUX2_X1 U9740 ( .A(_02589__PTR18), .B(_02588__PTR18), .S(P3_READY_n), .Z(_02594__PTR18) );
  MUX2_X1 U9741 ( .A(_02589__PTR19), .B(_02588__PTR19), .S(P3_READY_n), .Z(_02594__PTR19) );
  MUX2_X1 U9742 ( .A(_02589__PTR20), .B(_02588__PTR20), .S(P3_READY_n), .Z(_02594__PTR20) );
  MUX2_X1 U9743 ( .A(_02589__PTR21), .B(_02588__PTR21), .S(P3_READY_n), .Z(_02594__PTR21) );
  MUX2_X1 U9744 ( .A(_02589__PTR22), .B(_02588__PTR22), .S(P3_READY_n), .Z(_02594__PTR22) );
  MUX2_X1 U9745 ( .A(_02589__PTR23), .B(_02588__PTR23), .S(P3_READY_n), .Z(_02594__PTR23) );
  MUX2_X1 U9746 ( .A(_02589__PTR24), .B(_02588__PTR24), .S(P3_READY_n), .Z(_02594__PTR24) );
  MUX2_X1 U9747 ( .A(_02589__PTR25), .B(_02588__PTR25), .S(P3_READY_n), .Z(_02594__PTR25) );
  MUX2_X1 U9748 ( .A(_02589__PTR26), .B(_02588__PTR26), .S(P3_READY_n), .Z(_02594__PTR26) );
  MUX2_X1 U9749 ( .A(_02589__PTR27), .B(_02588__PTR27), .S(P3_READY_n), .Z(_02594__PTR27) );
  MUX2_X1 U9750 ( .A(_02589__PTR28), .B(_02588__PTR28), .S(P3_READY_n), .Z(_02594__PTR28) );
  MUX2_X1 U9751 ( .A(_02589__PTR29), .B(_02588__PTR29), .S(P3_READY_n), .Z(_02594__PTR29) );
  MUX2_X1 U9752 ( .A(_02589__PTR30), .B(_02588__PTR30), .S(P3_READY_n), .Z(_02594__PTR30) );
  MUX2_X1 U9753 ( .A(_02589__PTR31), .B(_02588__PTR31), .S(P3_READY_n), .Z(_02594__PTR31) );
  MUX2_X1 U9754 ( .A(buf2_PTR0), .B(P3_P1_lWord_PTR0), .S(P3_READY_n), .Z(_02593__PTR0) );
  MUX2_X1 U9755 ( .A(buf2_PTR1), .B(P3_P1_lWord_PTR1), .S(P3_READY_n), .Z(_02593__PTR1) );
  MUX2_X1 U9756 ( .A(buf2_PTR2), .B(P3_P1_lWord_PTR2), .S(P3_READY_n), .Z(_02593__PTR2) );
  MUX2_X1 U9757 ( .A(buf2_PTR3), .B(P3_P1_lWord_PTR3), .S(P3_READY_n), .Z(_02593__PTR3) );
  MUX2_X1 U9758 ( .A(buf2_PTR4), .B(P3_P1_lWord_PTR4), .S(P3_READY_n), .Z(_02593__PTR4) );
  MUX2_X1 U9759 ( .A(buf2_PTR5), .B(P3_P1_lWord_PTR5), .S(P3_READY_n), .Z(_02593__PTR5) );
  MUX2_X1 U9760 ( .A(buf2_PTR6), .B(P3_P1_lWord_PTR6), .S(P3_READY_n), .Z(_02593__PTR6) );
  MUX2_X1 U9761 ( .A(buf2_PTR7), .B(P3_P1_lWord_PTR7), .S(P3_READY_n), .Z(_02593__PTR7) );
  MUX2_X1 U9762 ( .A(buf2_PTR8), .B(P3_P1_lWord_PTR8), .S(P3_READY_n), .Z(_02593__PTR8) );
  MUX2_X1 U9763 ( .A(buf2_PTR9), .B(P3_P1_lWord_PTR9), .S(P3_READY_n), .Z(_02593__PTR9) );
  MUX2_X1 U9764 ( .A(buf2_PTR10), .B(P3_P1_lWord_PTR10), .S(P3_READY_n), .Z(_02593__PTR10) );
  MUX2_X1 U9765 ( .A(buf2_PTR11), .B(P3_P1_lWord_PTR11), .S(P3_READY_n), .Z(_02593__PTR11) );
  MUX2_X1 U9766 ( .A(buf2_PTR12), .B(P3_P1_lWord_PTR12), .S(P3_READY_n), .Z(_02593__PTR12) );
  MUX2_X1 U9767 ( .A(buf2_PTR13), .B(P3_P1_lWord_PTR13), .S(P3_READY_n), .Z(_02593__PTR13) );
  MUX2_X1 U9768 ( .A(buf2_PTR14), .B(P3_P1_lWord_PTR14), .S(P3_READY_n), .Z(_02593__PTR14) );
  MUX2_X1 U9769 ( .A(buf2_PTR15), .B(P3_P1_lWord_PTR15), .S(P3_READY_n), .Z(_02593__PTR15) );
  MUX2_X1 U9770 ( .A(buf2_PTR0), .B(P3_P1_uWord_PTR0), .S(P3_READY_n), .Z(_02592__PTR0) );
  MUX2_X1 U9771 ( .A(buf2_PTR1), .B(P3_P1_uWord_PTR1), .S(P3_READY_n), .Z(_02592__PTR1) );
  MUX2_X1 U9772 ( .A(buf2_PTR2), .B(P3_P1_uWord_PTR2), .S(P3_READY_n), .Z(_02592__PTR2) );
  MUX2_X1 U9773 ( .A(buf2_PTR3), .B(P3_P1_uWord_PTR3), .S(P3_READY_n), .Z(_02592__PTR3) );
  MUX2_X1 U9774 ( .A(buf2_PTR4), .B(P3_P1_uWord_PTR4), .S(P3_READY_n), .Z(_02592__PTR4) );
  MUX2_X1 U9775 ( .A(buf2_PTR5), .B(P3_P1_uWord_PTR5), .S(P3_READY_n), .Z(_02592__PTR5) );
  MUX2_X1 U9776 ( .A(buf2_PTR6), .B(P3_P1_uWord_PTR6), .S(P3_READY_n), .Z(_02592__PTR6) );
  MUX2_X1 U9777 ( .A(buf2_PTR7), .B(P3_P1_uWord_PTR7), .S(P3_READY_n), .Z(_02592__PTR7) );
  MUX2_X1 U9778 ( .A(buf2_PTR8), .B(P3_P1_uWord_PTR8), .S(P3_READY_n), .Z(_02592__PTR8) );
  MUX2_X1 U9779 ( .A(buf2_PTR9), .B(P3_P1_uWord_PTR9), .S(P3_READY_n), .Z(_02592__PTR9) );
  MUX2_X1 U9780 ( .A(buf2_PTR10), .B(P3_P1_uWord_PTR10), .S(P3_READY_n), .Z(_02592__PTR10) );
  MUX2_X1 U9781 ( .A(buf2_PTR11), .B(P3_P1_uWord_PTR11), .S(P3_READY_n), .Z(_02592__PTR11) );
  MUX2_X1 U9782 ( .A(buf2_PTR12), .B(P3_P1_uWord_PTR12), .S(P3_READY_n), .Z(_02592__PTR12) );
  MUX2_X1 U9783 ( .A(buf2_PTR13), .B(P3_P1_uWord_PTR13), .S(P3_READY_n), .Z(_02592__PTR13) );
  MUX2_X1 U9784 ( .A(buf2_PTR14), .B(P3_P1_uWord_PTR14), .S(P3_READY_n), .Z(_02592__PTR14) );
  MUX2_X1 U9785 ( .A(P3_P1_InstAddrPointer_PTR0), .B(_02662__PTR0), .S(_02435__PTR2), .Z(_02662__PTR128) );
  MUX2_X1 U9786 ( .A(P3_P1_InstAddrPointer_PTR1), .B(_02662__PTR1), .S(_02435__PTR2), .Z(_02662__PTR129) );
  MUX2_X1 U9787 ( .A(P3_P1_InstAddrPointer_PTR2), .B(_03297__PTR2), .S(_02435__PTR2), .Z(_02662__PTR130) );
  MUX2_X1 U9788 ( .A(P3_P1_InstAddrPointer_PTR3), .B(_03297__PTR3), .S(_02435__PTR2), .Z(_02662__PTR131) );
  MUX2_X1 U9789 ( .A(P3_P1_InstAddrPointer_PTR4), .B(_03297__PTR4), .S(_02435__PTR2), .Z(_02662__PTR132) );
  MUX2_X1 U9790 ( .A(P3_P1_InstAddrPointer_PTR5), .B(_03297__PTR5), .S(_02435__PTR2), .Z(_02662__PTR133) );
  MUX2_X1 U9791 ( .A(P3_P1_InstAddrPointer_PTR6), .B(_03297__PTR6), .S(_02435__PTR2), .Z(_02662__PTR134) );
  MUX2_X1 U9792 ( .A(P3_P1_InstAddrPointer_PTR7), .B(_03297__PTR7), .S(_02435__PTR2), .Z(_02662__PTR135) );
  MUX2_X1 U9793 ( .A(P3_P1_InstAddrPointer_PTR8), .B(_03297__PTR8), .S(_02435__PTR2), .Z(_02662__PTR136) );
  MUX2_X1 U9794 ( .A(P3_P1_InstAddrPointer_PTR9), .B(_03297__PTR9), .S(_02435__PTR2), .Z(_02662__PTR137) );
  MUX2_X1 U9795 ( .A(P3_P1_InstAddrPointer_PTR10), .B(_03297__PTR10), .S(_02435__PTR2), .Z(_02662__PTR138) );
  MUX2_X1 U9796 ( .A(P3_P1_InstAddrPointer_PTR11), .B(_03297__PTR11), .S(_02435__PTR2), .Z(_02662__PTR139) );
  MUX2_X1 U9797 ( .A(P3_P1_InstAddrPointer_PTR12), .B(_03297__PTR12), .S(_02435__PTR2), .Z(_02662__PTR140) );
  MUX2_X1 U9798 ( .A(P3_P1_InstAddrPointer_PTR13), .B(_03297__PTR13), .S(_02435__PTR2), .Z(_02662__PTR141) );
  MUX2_X1 U9799 ( .A(P3_P1_InstAddrPointer_PTR14), .B(_03297__PTR14), .S(_02435__PTR2), .Z(_02662__PTR142) );
  MUX2_X1 U9800 ( .A(P3_P1_InstAddrPointer_PTR15), .B(_03297__PTR15), .S(_02435__PTR2), .Z(_02662__PTR143) );
  MUX2_X1 U9801 ( .A(P3_P1_InstAddrPointer_PTR16), .B(_03297__PTR16), .S(_02435__PTR2), .Z(_02662__PTR144) );
  MUX2_X1 U9802 ( .A(P3_P1_InstAddrPointer_PTR17), .B(_03297__PTR17), .S(_02435__PTR2), .Z(_02662__PTR145) );
  MUX2_X1 U9803 ( .A(P3_P1_InstAddrPointer_PTR18), .B(_03297__PTR18), .S(_02435__PTR2), .Z(_02662__PTR146) );
  MUX2_X1 U9804 ( .A(P3_P1_InstAddrPointer_PTR19), .B(_03297__PTR19), .S(_02435__PTR2), .Z(_02662__PTR147) );
  MUX2_X1 U9805 ( .A(P3_P1_InstAddrPointer_PTR20), .B(_03297__PTR20), .S(_02435__PTR2), .Z(_02662__PTR148) );
  MUX2_X1 U9806 ( .A(P3_P1_InstAddrPointer_PTR21), .B(_03297__PTR21), .S(_02435__PTR2), .Z(_02662__PTR149) );
  MUX2_X1 U9807 ( .A(P3_P1_InstAddrPointer_PTR22), .B(_03297__PTR22), .S(_02435__PTR2), .Z(_02662__PTR150) );
  MUX2_X1 U9808 ( .A(P3_P1_InstAddrPointer_PTR23), .B(_03297__PTR23), .S(_02435__PTR2), .Z(_02662__PTR151) );
  MUX2_X1 U9809 ( .A(P3_P1_InstAddrPointer_PTR24), .B(_03297__PTR24), .S(_02435__PTR2), .Z(_02662__PTR152) );
  MUX2_X1 U9810 ( .A(P3_P1_InstAddrPointer_PTR25), .B(_03297__PTR25), .S(_02435__PTR2), .Z(_02662__PTR153) );
  MUX2_X1 U9811 ( .A(P3_P1_InstAddrPointer_PTR26), .B(_03297__PTR26), .S(_02435__PTR2), .Z(_02662__PTR154) );
  MUX2_X1 U9812 ( .A(P3_P1_InstAddrPointer_PTR27), .B(_03297__PTR27), .S(_02435__PTR2), .Z(_02662__PTR155) );
  MUX2_X1 U9813 ( .A(P3_P1_InstAddrPointer_PTR28), .B(_03297__PTR28), .S(_02435__PTR2), .Z(_02662__PTR156) );
  MUX2_X1 U9814 ( .A(P3_P1_InstAddrPointer_PTR29), .B(_03297__PTR29), .S(_02435__PTR2), .Z(_02662__PTR157) );
  MUX2_X1 U9815 ( .A(P3_P1_InstAddrPointer_PTR30), .B(_03297__PTR30), .S(_02435__PTR2), .Z(_02662__PTR158) );
  MUX2_X1 U9816 ( .A(P3_P1_InstAddrPointer_PTR31), .B(_03297__PTR31), .S(_02435__PTR2), .Z(_02662__PTR159) );
  MUX2_X1 U9817 ( .A(P3_P1_InstAddrPointer_PTR0), .B(_03299__PTR0), .S(_02435__PTR2), .Z(_02662__PTR160) );
  MUX2_X1 U9818 ( .A(P3_P1_InstAddrPointer_PTR1), .B(_03300__PTR1), .S(_02435__PTR2), .Z(_02662__PTR161) );
  MUX2_X1 U9819 ( .A(P3_P1_InstAddrPointer_PTR2), .B(_03300__PTR2), .S(_02435__PTR2), .Z(_02662__PTR162) );
  MUX2_X1 U9820 ( .A(P3_P1_InstAddrPointer_PTR3), .B(_03300__PTR3), .S(_02435__PTR2), .Z(_02662__PTR163) );
  MUX2_X1 U9821 ( .A(P3_P1_InstAddrPointer_PTR4), .B(_03300__PTR4), .S(_02435__PTR2), .Z(_02662__PTR164) );
  MUX2_X1 U9822 ( .A(P3_P1_InstAddrPointer_PTR5), .B(_03300__PTR5), .S(_02435__PTR2), .Z(_02662__PTR165) );
  MUX2_X1 U9823 ( .A(P3_P1_InstAddrPointer_PTR6), .B(_03300__PTR6), .S(_02435__PTR2), .Z(_02662__PTR166) );
  MUX2_X1 U9824 ( .A(P3_P1_InstAddrPointer_PTR7), .B(_03300__PTR7), .S(_02435__PTR2), .Z(_02662__PTR167) );
  MUX2_X1 U9825 ( .A(P3_P1_InstAddrPointer_PTR8), .B(_03300__PTR8), .S(_02435__PTR2), .Z(_02662__PTR168) );
  MUX2_X1 U9826 ( .A(P3_P1_InstAddrPointer_PTR9), .B(_03300__PTR9), .S(_02435__PTR2), .Z(_02662__PTR169) );
  MUX2_X1 U9827 ( .A(P3_P1_InstAddrPointer_PTR10), .B(_03300__PTR10), .S(_02435__PTR2), .Z(_02662__PTR170) );
  MUX2_X1 U9828 ( .A(P3_P1_InstAddrPointer_PTR11), .B(_03300__PTR11), .S(_02435__PTR2), .Z(_02662__PTR171) );
  MUX2_X1 U9829 ( .A(P3_P1_InstAddrPointer_PTR12), .B(_03300__PTR12), .S(_02435__PTR2), .Z(_02662__PTR172) );
  MUX2_X1 U9830 ( .A(P3_P1_InstAddrPointer_PTR13), .B(_03300__PTR13), .S(_02435__PTR2), .Z(_02662__PTR173) );
  MUX2_X1 U9831 ( .A(P3_P1_InstAddrPointer_PTR14), .B(_03300__PTR14), .S(_02435__PTR2), .Z(_02662__PTR174) );
  MUX2_X1 U9832 ( .A(P3_P1_InstAddrPointer_PTR15), .B(_03300__PTR15), .S(_02435__PTR2), .Z(_02662__PTR175) );
  MUX2_X1 U9833 ( .A(P3_P1_InstAddrPointer_PTR16), .B(_03300__PTR16), .S(_02435__PTR2), .Z(_02662__PTR176) );
  MUX2_X1 U9834 ( .A(P3_P1_InstAddrPointer_PTR17), .B(_03300__PTR17), .S(_02435__PTR2), .Z(_02662__PTR177) );
  MUX2_X1 U9835 ( .A(P3_P1_InstAddrPointer_PTR18), .B(_03300__PTR18), .S(_02435__PTR2), .Z(_02662__PTR178) );
  MUX2_X1 U9836 ( .A(P3_P1_InstAddrPointer_PTR19), .B(_03300__PTR19), .S(_02435__PTR2), .Z(_02662__PTR179) );
  MUX2_X1 U9837 ( .A(P3_P1_InstAddrPointer_PTR20), .B(_03300__PTR20), .S(_02435__PTR2), .Z(_02662__PTR180) );
  MUX2_X1 U9838 ( .A(P3_P1_InstAddrPointer_PTR21), .B(_03300__PTR21), .S(_02435__PTR2), .Z(_02662__PTR181) );
  MUX2_X1 U9839 ( .A(P3_P1_InstAddrPointer_PTR22), .B(_03300__PTR22), .S(_02435__PTR2), .Z(_02662__PTR182) );
  MUX2_X1 U9840 ( .A(P3_P1_InstAddrPointer_PTR23), .B(_03300__PTR23), .S(_02435__PTR2), .Z(_02662__PTR183) );
  MUX2_X1 U9841 ( .A(P3_P1_InstAddrPointer_PTR24), .B(_03300__PTR24), .S(_02435__PTR2), .Z(_02662__PTR184) );
  MUX2_X1 U9842 ( .A(P3_P1_InstAddrPointer_PTR25), .B(_03300__PTR25), .S(_02435__PTR2), .Z(_02662__PTR185) );
  MUX2_X1 U9843 ( .A(P3_P1_InstAddrPointer_PTR26), .B(_03300__PTR26), .S(_02435__PTR2), .Z(_02662__PTR186) );
  MUX2_X1 U9844 ( .A(P3_P1_InstAddrPointer_PTR27), .B(_03300__PTR27), .S(_02435__PTR2), .Z(_02662__PTR187) );
  MUX2_X1 U9845 ( .A(P3_P1_InstAddrPointer_PTR28), .B(_03300__PTR28), .S(_02435__PTR2), .Z(_02662__PTR188) );
  MUX2_X1 U9846 ( .A(P3_P1_InstAddrPointer_PTR29), .B(_03300__PTR29), .S(_02435__PTR2), .Z(_02662__PTR189) );
  MUX2_X1 U9847 ( .A(P3_P1_InstAddrPointer_PTR30), .B(_03300__PTR30), .S(_02435__PTR2), .Z(_02662__PTR190) );
  MUX2_X1 U9848 ( .A(P3_P1_InstAddrPointer_PTR31), .B(_03300__PTR31), .S(_02435__PTR2), .Z(_02662__PTR191) );
  MUX2_X1 U9849 ( .A(P3_rEIP_PTR0), .B(_02465__PTR3), .S(_02585_), .Z(_02682__PTR32) );
  MUX2_X1 U9850 ( .A(P3_rEIP_PTR1), .B(_02465__PTR4), .S(_02585_), .Z(_02682__PTR33) );
  MUX2_X1 U9851 ( .A(P3_rEIP_PTR2), .B(_02465__PTR5), .S(_02585_), .Z(_02682__PTR34) );
  MUX2_X1 U9852 ( .A(P3_rEIP_PTR3), .B(_02465__PTR6), .S(_02585_), .Z(_02682__PTR35) );
  MUX2_X1 U9853 ( .A(P3_rEIP_PTR4), .B(_03290__PTR4), .S(_02585_), .Z(_02682__PTR36) );
  MUX2_X1 U9854 ( .A(P3_rEIP_PTR5), .B(_03289__PTR4), .S(_02585_), .Z(_02682__PTR37) );
  MUX2_X1 U9855 ( .A(P3_rEIP_PTR6), .B(1'b0), .S(_02585_), .Z(_02682__PTR38) );
  MUX2_X1 U9856 ( .A(P3_rEIP_PTR7), .B(1'b0), .S(_02585_), .Z(_02682__PTR39) );
  MUX2_X1 U9857 ( .A(P3_rEIP_PTR8), .B(1'b0), .S(_02585_), .Z(_02682__PTR40) );
  MUX2_X1 U9858 ( .A(P3_rEIP_PTR9), .B(1'b0), .S(_02585_), .Z(_02682__PTR41) );
  MUX2_X1 U9859 ( .A(P3_rEIP_PTR10), .B(1'b0), .S(_02585_), .Z(_02682__PTR42) );
  MUX2_X1 U9860 ( .A(P3_rEIP_PTR11), .B(1'b0), .S(_02585_), .Z(_02682__PTR43) );
  MUX2_X1 U9861 ( .A(P3_rEIP_PTR12), .B(1'b0), .S(_02585_), .Z(_02682__PTR44) );
  MUX2_X1 U9862 ( .A(P3_rEIP_PTR13), .B(1'b0), .S(_02585_), .Z(_02682__PTR45) );
  MUX2_X1 U9863 ( .A(P3_rEIP_PTR14), .B(1'b0), .S(_02585_), .Z(_02682__PTR46) );
  MUX2_X1 U9864 ( .A(P3_rEIP_PTR15), .B(1'b0), .S(_02585_), .Z(_02682__PTR47) );
  MUX2_X1 U9865 ( .A(P3_rEIP_PTR16), .B(1'b0), .S(_02585_), .Z(_02682__PTR48) );
  MUX2_X1 U9866 ( .A(P3_rEIP_PTR17), .B(1'b0), .S(_02585_), .Z(_02682__PTR49) );
  MUX2_X1 U9867 ( .A(P3_rEIP_PTR18), .B(1'b0), .S(_02585_), .Z(_02682__PTR50) );
  MUX2_X1 U9868 ( .A(P3_rEIP_PTR19), .B(1'b0), .S(_02585_), .Z(_02682__PTR51) );
  MUX2_X1 U9869 ( .A(P3_rEIP_PTR20), .B(1'b0), .S(_02585_), .Z(_02682__PTR52) );
  MUX2_X1 U9870 ( .A(P3_rEIP_PTR21), .B(1'b0), .S(_02585_), .Z(_02682__PTR53) );
  MUX2_X1 U9871 ( .A(P3_rEIP_PTR22), .B(1'b0), .S(_02585_), .Z(_02682__PTR54) );
  MUX2_X1 U9872 ( .A(P3_rEIP_PTR23), .B(1'b0), .S(_02585_), .Z(_02682__PTR55) );
  MUX2_X1 U9873 ( .A(P3_rEIP_PTR24), .B(1'b0), .S(_02585_), .Z(_02682__PTR56) );
  MUX2_X1 U9874 ( .A(P3_rEIP_PTR25), .B(1'b0), .S(_02585_), .Z(_02682__PTR57) );
  MUX2_X1 U9875 ( .A(P3_rEIP_PTR26), .B(1'b0), .S(_02585_), .Z(_02682__PTR58) );
  MUX2_X1 U9876 ( .A(P3_rEIP_PTR27), .B(1'b0), .S(_02585_), .Z(_02682__PTR59) );
  MUX2_X1 U9877 ( .A(P3_rEIP_PTR28), .B(1'b0), .S(_02585_), .Z(_02682__PTR60) );
  MUX2_X1 U9878 ( .A(P3_rEIP_PTR29), .B(1'b0), .S(_02585_), .Z(_02682__PTR61) );
  MUX2_X1 U9879 ( .A(P3_rEIP_PTR30), .B(1'b0), .S(_02585_), .Z(_02682__PTR62) );
  MUX2_X1 U9880 ( .A(P3_rEIP_PTR31), .B(1'b0), .S(_02585_), .Z(_02682__PTR63) );
  MUX2_X1 U9881 ( .A(P3_rEIP_PTR0), .B(_02612__PTR0), .S(_02585_), .Z(_02682__PTR64) );
  MUX2_X1 U9882 ( .A(P3_rEIP_PTR1), .B(_02612__PTR1), .S(_02585_), .Z(_02682__PTR65) );
  MUX2_X1 U9883 ( .A(P3_rEIP_PTR2), .B(_02612__PTR2), .S(_02585_), .Z(_02682__PTR66) );
  MUX2_X1 U9884 ( .A(P3_rEIP_PTR3), .B(_02612__PTR3), .S(_02585_), .Z(_02682__PTR67) );
  MUX2_X1 U9885 ( .A(P3_rEIP_PTR4), .B(_02612__PTR4), .S(_02585_), .Z(_02682__PTR68) );
  MUX2_X1 U9886 ( .A(P3_rEIP_PTR5), .B(_02612__PTR5), .S(_02585_), .Z(_02682__PTR69) );
  MUX2_X1 U9887 ( .A(P3_rEIP_PTR6), .B(_02612__PTR6), .S(_02585_), .Z(_02682__PTR70) );
  MUX2_X1 U9888 ( .A(P3_rEIP_PTR7), .B(_02612__PTR7), .S(_02585_), .Z(_02682__PTR71) );
  MUX2_X1 U9889 ( .A(P3_rEIP_PTR8), .B(_02612__PTR8), .S(_02585_), .Z(_02682__PTR72) );
  MUX2_X1 U9890 ( .A(P3_rEIP_PTR9), .B(_02612__PTR9), .S(_02585_), .Z(_02682__PTR73) );
  MUX2_X1 U9891 ( .A(P3_rEIP_PTR10), .B(_02612__PTR10), .S(_02585_), .Z(_02682__PTR74) );
  MUX2_X1 U9892 ( .A(P3_rEIP_PTR11), .B(_02612__PTR11), .S(_02585_), .Z(_02682__PTR75) );
  MUX2_X1 U9893 ( .A(P3_rEIP_PTR12), .B(_02612__PTR12), .S(_02585_), .Z(_02682__PTR76) );
  MUX2_X1 U9894 ( .A(P3_rEIP_PTR13), .B(_02612__PTR13), .S(_02585_), .Z(_02682__PTR77) );
  MUX2_X1 U9895 ( .A(P3_rEIP_PTR14), .B(_02612__PTR14), .S(_02585_), .Z(_02682__PTR78) );
  MUX2_X1 U9896 ( .A(P3_rEIP_PTR15), .B(_02612__PTR15), .S(_02585_), .Z(_02682__PTR79) );
  MUX2_X1 U9897 ( .A(P3_rEIP_PTR16), .B(_02612__PTR16), .S(_02585_), .Z(_02682__PTR80) );
  MUX2_X1 U9898 ( .A(P3_rEIP_PTR17), .B(_02612__PTR17), .S(_02585_), .Z(_02682__PTR81) );
  MUX2_X1 U9899 ( .A(P3_rEIP_PTR18), .B(_02612__PTR18), .S(_02585_), .Z(_02682__PTR82) );
  MUX2_X1 U9900 ( .A(P3_rEIP_PTR19), .B(_02612__PTR19), .S(_02585_), .Z(_02682__PTR83) );
  MUX2_X1 U9901 ( .A(P3_rEIP_PTR20), .B(_02612__PTR20), .S(_02585_), .Z(_02682__PTR84) );
  MUX2_X1 U9902 ( .A(P3_rEIP_PTR21), .B(_02612__PTR21), .S(_02585_), .Z(_02682__PTR85) );
  MUX2_X1 U9903 ( .A(P3_rEIP_PTR22), .B(_02612__PTR22), .S(_02585_), .Z(_02682__PTR86) );
  MUX2_X1 U9904 ( .A(P3_rEIP_PTR23), .B(_02612__PTR23), .S(_02585_), .Z(_02682__PTR87) );
  MUX2_X1 U9905 ( .A(P3_rEIP_PTR24), .B(_02612__PTR24), .S(_02585_), .Z(_02682__PTR88) );
  MUX2_X1 U9906 ( .A(P3_rEIP_PTR25), .B(_02612__PTR25), .S(_02585_), .Z(_02682__PTR89) );
  MUX2_X1 U9907 ( .A(P3_rEIP_PTR26), .B(_02612__PTR26), .S(_02585_), .Z(_02682__PTR90) );
  MUX2_X1 U9908 ( .A(P3_rEIP_PTR27), .B(_02612__PTR27), .S(_02585_), .Z(_02682__PTR91) );
  MUX2_X1 U9909 ( .A(P3_rEIP_PTR28), .B(_02612__PTR28), .S(_02585_), .Z(_02682__PTR92) );
  MUX2_X1 U9910 ( .A(P3_rEIP_PTR29), .B(_02612__PTR29), .S(_02585_), .Z(_02682__PTR93) );
  MUX2_X1 U9911 ( .A(P3_rEIP_PTR30), .B(_02612__PTR30), .S(_02585_), .Z(_02682__PTR94) );
  MUX2_X1 U9912 ( .A(P3_rEIP_PTR31), .B(_02612__PTR31), .S(_02585_), .Z(_02682__PTR95) );
  MUX2_X1 U9913 ( .A(P3_rEIP_PTR0), .B(_02594__PTR0), .S(_02585_), .Z(_02682__PTR96) );
  MUX2_X1 U9914 ( .A(P3_rEIP_PTR1), .B(_02594__PTR1), .S(_02585_), .Z(_02682__PTR97) );
  MUX2_X1 U9915 ( .A(P3_rEIP_PTR2), .B(_02594__PTR2), .S(_02585_), .Z(_02682__PTR98) );
  MUX2_X1 U9916 ( .A(P3_rEIP_PTR3), .B(_02594__PTR3), .S(_02585_), .Z(_02682__PTR99) );
  MUX2_X1 U9917 ( .A(P3_rEIP_PTR4), .B(_02594__PTR4), .S(_02585_), .Z(_02682__PTR100) );
  MUX2_X1 U9918 ( .A(P3_rEIP_PTR5), .B(_02594__PTR5), .S(_02585_), .Z(_02682__PTR101) );
  MUX2_X1 U9919 ( .A(P3_rEIP_PTR6), .B(_02594__PTR6), .S(_02585_), .Z(_02682__PTR102) );
  MUX2_X1 U9920 ( .A(P3_rEIP_PTR7), .B(_02594__PTR7), .S(_02585_), .Z(_02682__PTR103) );
  MUX2_X1 U9921 ( .A(P3_rEIP_PTR8), .B(_02594__PTR8), .S(_02585_), .Z(_02682__PTR104) );
  MUX2_X1 U9922 ( .A(P3_rEIP_PTR9), .B(_02594__PTR9), .S(_02585_), .Z(_02682__PTR105) );
  MUX2_X1 U9923 ( .A(P3_rEIP_PTR10), .B(_02594__PTR10), .S(_02585_), .Z(_02682__PTR106) );
  MUX2_X1 U9924 ( .A(P3_rEIP_PTR11), .B(_02594__PTR11), .S(_02585_), .Z(_02682__PTR107) );
  MUX2_X1 U9925 ( .A(P3_rEIP_PTR12), .B(_02594__PTR12), .S(_02585_), .Z(_02682__PTR108) );
  MUX2_X1 U9926 ( .A(P3_rEIP_PTR13), .B(_02594__PTR13), .S(_02585_), .Z(_02682__PTR109) );
  MUX2_X1 U9927 ( .A(P3_rEIP_PTR14), .B(_02594__PTR14), .S(_02585_), .Z(_02682__PTR110) );
  MUX2_X1 U9928 ( .A(P3_rEIP_PTR15), .B(_02594__PTR15), .S(_02585_), .Z(_02682__PTR111) );
  MUX2_X1 U9929 ( .A(P3_rEIP_PTR16), .B(_02594__PTR16), .S(_02585_), .Z(_02682__PTR112) );
  MUX2_X1 U9930 ( .A(P3_rEIP_PTR17), .B(_02594__PTR17), .S(_02585_), .Z(_02682__PTR113) );
  MUX2_X1 U9931 ( .A(P3_rEIP_PTR18), .B(_02594__PTR18), .S(_02585_), .Z(_02682__PTR114) );
  MUX2_X1 U9932 ( .A(P3_rEIP_PTR19), .B(_02594__PTR19), .S(_02585_), .Z(_02682__PTR115) );
  MUX2_X1 U9933 ( .A(P3_rEIP_PTR20), .B(_02594__PTR20), .S(_02585_), .Z(_02682__PTR116) );
  MUX2_X1 U9934 ( .A(P3_rEIP_PTR21), .B(_02594__PTR21), .S(_02585_), .Z(_02682__PTR117) );
  MUX2_X1 U9935 ( .A(P3_rEIP_PTR22), .B(_02594__PTR22), .S(_02585_), .Z(_02682__PTR118) );
  MUX2_X1 U9936 ( .A(P3_rEIP_PTR23), .B(_02594__PTR23), .S(_02585_), .Z(_02682__PTR119) );
  MUX2_X1 U9937 ( .A(P3_rEIP_PTR24), .B(_02594__PTR24), .S(_02585_), .Z(_02682__PTR120) );
  MUX2_X1 U9938 ( .A(P3_rEIP_PTR25), .B(_02594__PTR25), .S(_02585_), .Z(_02682__PTR121) );
  MUX2_X1 U9939 ( .A(P3_rEIP_PTR26), .B(_02594__PTR26), .S(_02585_), .Z(_02682__PTR122) );
  MUX2_X1 U9940 ( .A(P3_rEIP_PTR27), .B(_02594__PTR27), .S(_02585_), .Z(_02682__PTR123) );
  MUX2_X1 U9941 ( .A(P3_rEIP_PTR28), .B(_02594__PTR28), .S(_02585_), .Z(_02682__PTR124) );
  MUX2_X1 U9942 ( .A(P3_rEIP_PTR29), .B(_02594__PTR29), .S(_02585_), .Z(_02682__PTR125) );
  MUX2_X1 U9943 ( .A(P3_rEIP_PTR30), .B(_02594__PTR30), .S(_02585_), .Z(_02682__PTR126) );
  MUX2_X1 U9944 ( .A(P3_rEIP_PTR31), .B(_02594__PTR31), .S(_02585_), .Z(_02682__PTR127) );
  MUX2_X1 U9945 ( .A(P3_rEIP_PTR0), .B(P3_EBX_PTR0), .S(P3_StateBS16), .Z(_02589__PTR0) );
  MUX2_X1 U9946 ( .A(_02463__PTR7), .B(_02588__PTR1), .S(P3_StateBS16), .Z(_02589__PTR1) );
  MUX2_X1 U9947 ( .A(_03312__PTR1), .B(_02588__PTR2), .S(P3_StateBS16), .Z(_02589__PTR2) );
  MUX2_X1 U9948 ( .A(_03312__PTR2), .B(_02588__PTR3), .S(P3_StateBS16), .Z(_02589__PTR3) );
  MUX2_X1 U9949 ( .A(_03312__PTR3), .B(_02588__PTR4), .S(P3_StateBS16), .Z(_02589__PTR4) );
  MUX2_X1 U9950 ( .A(_03312__PTR4), .B(_02588__PTR5), .S(P3_StateBS16), .Z(_02589__PTR5) );
  MUX2_X1 U9951 ( .A(_03312__PTR5), .B(_02588__PTR6), .S(P3_StateBS16), .Z(_02589__PTR6) );
  MUX2_X1 U9952 ( .A(_03312__PTR6), .B(_02588__PTR7), .S(P3_StateBS16), .Z(_02589__PTR7) );
  MUX2_X1 U9953 ( .A(_03312__PTR7), .B(_02588__PTR8), .S(P3_StateBS16), .Z(_02589__PTR8) );
  MUX2_X1 U9954 ( .A(_03312__PTR8), .B(_02588__PTR9), .S(P3_StateBS16), .Z(_02589__PTR9) );
  MUX2_X1 U9955 ( .A(_03312__PTR9), .B(_02588__PTR10), .S(P3_StateBS16), .Z(_02589__PTR10) );
  MUX2_X1 U9956 ( .A(_03312__PTR10), .B(_02588__PTR11), .S(P3_StateBS16), .Z(_02589__PTR11) );
  MUX2_X1 U9957 ( .A(_03312__PTR11), .B(_02588__PTR12), .S(P3_StateBS16), .Z(_02589__PTR12) );
  MUX2_X1 U9958 ( .A(_03312__PTR12), .B(_02588__PTR13), .S(P3_StateBS16), .Z(_02589__PTR13) );
  MUX2_X1 U9959 ( .A(_03312__PTR13), .B(_02588__PTR14), .S(P3_StateBS16), .Z(_02589__PTR14) );
  MUX2_X1 U9960 ( .A(_03312__PTR14), .B(_02588__PTR15), .S(P3_StateBS16), .Z(_02589__PTR15) );
  MUX2_X1 U9961 ( .A(_03312__PTR15), .B(_02588__PTR16), .S(P3_StateBS16), .Z(_02589__PTR16) );
  MUX2_X1 U9962 ( .A(_03312__PTR16), .B(_02588__PTR17), .S(P3_StateBS16), .Z(_02589__PTR17) );
  MUX2_X1 U9963 ( .A(_03312__PTR17), .B(_02588__PTR18), .S(P3_StateBS16), .Z(_02589__PTR18) );
  MUX2_X1 U9964 ( .A(_03312__PTR18), .B(_02588__PTR19), .S(P3_StateBS16), .Z(_02589__PTR19) );
  MUX2_X1 U9965 ( .A(_03312__PTR19), .B(_02588__PTR20), .S(P3_StateBS16), .Z(_02589__PTR20) );
  MUX2_X1 U9966 ( .A(_03312__PTR20), .B(_02588__PTR21), .S(P3_StateBS16), .Z(_02589__PTR21) );
  MUX2_X1 U9967 ( .A(_03312__PTR21), .B(_02588__PTR22), .S(P3_StateBS16), .Z(_02589__PTR22) );
  MUX2_X1 U9968 ( .A(_03312__PTR22), .B(_02588__PTR23), .S(P3_StateBS16), .Z(_02589__PTR23) );
  MUX2_X1 U9969 ( .A(_03312__PTR23), .B(_02588__PTR24), .S(P3_StateBS16), .Z(_02589__PTR24) );
  MUX2_X1 U9970 ( .A(_03312__PTR24), .B(_02588__PTR25), .S(P3_StateBS16), .Z(_02589__PTR25) );
  MUX2_X1 U9971 ( .A(_03312__PTR25), .B(_02588__PTR26), .S(P3_StateBS16), .Z(_02589__PTR26) );
  MUX2_X1 U9972 ( .A(_03312__PTR26), .B(_02588__PTR27), .S(P3_StateBS16), .Z(_02589__PTR27) );
  MUX2_X1 U9973 ( .A(_03312__PTR27), .B(_02588__PTR28), .S(P3_StateBS16), .Z(_02589__PTR28) );
  MUX2_X1 U9974 ( .A(_03312__PTR28), .B(_02588__PTR29), .S(P3_StateBS16), .Z(_02589__PTR29) );
  MUX2_X1 U9975 ( .A(_03312__PTR29), .B(_02588__PTR30), .S(P3_StateBS16), .Z(_02589__PTR30) );
  MUX2_X1 U9976 ( .A(_03312__PTR30), .B(_02588__PTR31), .S(P3_StateBS16), .Z(_02589__PTR31) );
  MUX2_X1 U9977 ( .A(_03438__PTR1), .B(P3_EBX_PTR1), .S(_03223__PTR31), .Z(_02588__PTR1) );
  MUX2_X1 U9978 ( .A(_03438__PTR2), .B(P3_EBX_PTR2), .S(_03223__PTR31), .Z(_02588__PTR2) );
  MUX2_X1 U9979 ( .A(_03438__PTR3), .B(P3_EBX_PTR3), .S(_03223__PTR31), .Z(_02588__PTR3) );
  MUX2_X1 U9980 ( .A(_03438__PTR4), .B(P3_EBX_PTR4), .S(_03223__PTR31), .Z(_02588__PTR4) );
  MUX2_X1 U9981 ( .A(_03438__PTR5), .B(P3_EBX_PTR5), .S(_03223__PTR31), .Z(_02588__PTR5) );
  MUX2_X1 U9982 ( .A(_03438__PTR6), .B(P3_EBX_PTR6), .S(_03223__PTR31), .Z(_02588__PTR6) );
  MUX2_X1 U9983 ( .A(_03438__PTR7), .B(P3_EBX_PTR7), .S(_03223__PTR31), .Z(_02588__PTR7) );
  MUX2_X1 U9984 ( .A(_03438__PTR8), .B(P3_EBX_PTR8), .S(_03223__PTR31), .Z(_02588__PTR8) );
  MUX2_X1 U9985 ( .A(_03438__PTR9), .B(P3_EBX_PTR9), .S(_03223__PTR31), .Z(_02588__PTR9) );
  MUX2_X1 U9986 ( .A(_03438__PTR10), .B(P3_EBX_PTR10), .S(_03223__PTR31), .Z(_02588__PTR10) );
  MUX2_X1 U9987 ( .A(_03438__PTR11), .B(P3_EBX_PTR11), .S(_03223__PTR31), .Z(_02588__PTR11) );
  MUX2_X1 U9988 ( .A(_03438__PTR12), .B(P3_EBX_PTR12), .S(_03223__PTR31), .Z(_02588__PTR12) );
  MUX2_X1 U9989 ( .A(_03438__PTR13), .B(P3_EBX_PTR13), .S(_03223__PTR31), .Z(_02588__PTR13) );
  MUX2_X1 U9990 ( .A(_03438__PTR14), .B(P3_EBX_PTR14), .S(_03223__PTR31), .Z(_02588__PTR14) );
  MUX2_X1 U9991 ( .A(_03438__PTR15), .B(P3_EBX_PTR15), .S(_03223__PTR31), .Z(_02588__PTR15) );
  MUX2_X1 U9992 ( .A(_03438__PTR16), .B(P3_EBX_PTR16), .S(_03223__PTR31), .Z(_02588__PTR16) );
  MUX2_X1 U9993 ( .A(_03438__PTR17), .B(P3_EBX_PTR17), .S(_03223__PTR31), .Z(_02588__PTR17) );
  MUX2_X1 U9994 ( .A(_03438__PTR18), .B(P3_EBX_PTR18), .S(_03223__PTR31), .Z(_02588__PTR18) );
  MUX2_X1 U9995 ( .A(_03438__PTR19), .B(P3_EBX_PTR19), .S(_03223__PTR31), .Z(_02588__PTR19) );
  MUX2_X1 U9996 ( .A(_03438__PTR20), .B(P3_EBX_PTR20), .S(_03223__PTR31), .Z(_02588__PTR20) );
  MUX2_X1 U9997 ( .A(_03438__PTR21), .B(P3_EBX_PTR21), .S(_03223__PTR31), .Z(_02588__PTR21) );
  MUX2_X1 U9998 ( .A(_03438__PTR22), .B(P3_EBX_PTR22), .S(_03223__PTR31), .Z(_02588__PTR22) );
  MUX2_X1 U9999 ( .A(_03438__PTR23), .B(P3_EBX_PTR23), .S(_03223__PTR31), .Z(_02588__PTR23) );
  MUX2_X1 U10000 ( .A(_03438__PTR24), .B(P3_EBX_PTR24), .S(_03223__PTR31), .Z(_02588__PTR24) );
  MUX2_X1 U10001 ( .A(_03438__PTR25), .B(P3_EBX_PTR25), .S(_03223__PTR31), .Z(_02588__PTR25) );
  MUX2_X1 U10002 ( .A(_03438__PTR26), .B(P3_EBX_PTR26), .S(_03223__PTR31), .Z(_02588__PTR26) );
  MUX2_X1 U10003 ( .A(_03438__PTR27), .B(P3_EBX_PTR27), .S(_03223__PTR31), .Z(_02588__PTR27) );
  MUX2_X1 U10004 ( .A(_03438__PTR28), .B(P3_EBX_PTR28), .S(_03223__PTR31), .Z(_02588__PTR28) );
  MUX2_X1 U10005 ( .A(_03438__PTR29), .B(P3_EBX_PTR29), .S(_03223__PTR31), .Z(_02588__PTR29) );
  MUX2_X1 U10006 ( .A(_03438__PTR30), .B(P3_EBX_PTR30), .S(_03223__PTR31), .Z(_02588__PTR30) );
  MUX2_X1 U10007 ( .A(_03438__PTR31), .B(P3_EBX_PTR31), .S(_03223__PTR31), .Z(_02588__PTR31) );
  MUX2_X1 U10008 ( .A(P3_EBX_PTR0), .B(P3_P1_InstQueue_PTR0_PTR0), .S(_02435__PTR2), .Z(_02678__PTR64) );
  MUX2_X1 U10009 ( .A(P3_EBX_PTR1), .B(P3_P1_InstQueue_PTR0_PTR1), .S(_02435__PTR2), .Z(_02678__PTR65) );
  MUX2_X1 U10010 ( .A(P3_EBX_PTR2), .B(P3_P1_InstQueue_PTR0_PTR2), .S(_02435__PTR2), .Z(_02678__PTR66) );
  MUX2_X1 U10011 ( .A(P3_EBX_PTR3), .B(P3_P1_InstQueue_PTR0_PTR3), .S(_02435__PTR2), .Z(_02678__PTR67) );
  MUX2_X1 U10012 ( .A(P3_EBX_PTR4), .B(P3_P1_InstQueue_PTR0_PTR4), .S(_02435__PTR2), .Z(_02678__PTR68) );
  MUX2_X1 U10013 ( .A(P3_EBX_PTR5), .B(P3_P1_InstQueue_PTR0_PTR5), .S(_02435__PTR2), .Z(_02678__PTR69) );
  MUX2_X1 U10014 ( .A(P3_EBX_PTR6), .B(P3_P1_InstQueue_PTR0_PTR6), .S(_02435__PTR2), .Z(_02678__PTR70) );
  MUX2_X1 U10015 ( .A(P3_EBX_PTR7), .B(P3_P1_InstQueue_PTR0_PTR7), .S(_02435__PTR2), .Z(_02678__PTR71) );
  MUX2_X1 U10016 ( .A(P3_EBX_PTR8), .B(_02472__PTR0), .S(_02435__PTR2), .Z(_02678__PTR72) );
  MUX2_X1 U10017 ( .A(P3_EBX_PTR9), .B(_02472__PTR1), .S(_02435__PTR2), .Z(_02678__PTR73) );
  MUX2_X1 U10018 ( .A(P3_EBX_PTR10), .B(_02472__PTR2), .S(_02435__PTR2), .Z(_02678__PTR74) );
  MUX2_X1 U10019 ( .A(P3_EBX_PTR11), .B(_02472__PTR3), .S(_02435__PTR2), .Z(_02678__PTR75) );
  MUX2_X1 U10020 ( .A(P3_EBX_PTR12), .B(_02472__PTR4), .S(_02435__PTR2), .Z(_02678__PTR76) );
  MUX2_X1 U10021 ( .A(P3_EBX_PTR13), .B(_02472__PTR5), .S(_02435__PTR2), .Z(_02678__PTR77) );
  MUX2_X1 U10022 ( .A(P3_EBX_PTR14), .B(_02472__PTR6), .S(_02435__PTR2), .Z(_02678__PTR78) );
  MUX2_X1 U10023 ( .A(P3_EBX_PTR15), .B(_02472__PTR7), .S(_02435__PTR2), .Z(_02678__PTR79) );
  MUX2_X1 U10024 ( .A(P3_EBX_PTR16), .B(_02470__PTR0), .S(_02435__PTR2), .Z(_02678__PTR80) );
  MUX2_X1 U10025 ( .A(P3_EBX_PTR17), .B(_02470__PTR1), .S(_02435__PTR2), .Z(_02678__PTR81) );
  MUX2_X1 U10026 ( .A(P3_EBX_PTR18), .B(_02470__PTR2), .S(_02435__PTR2), .Z(_02678__PTR82) );
  MUX2_X1 U10027 ( .A(P3_EBX_PTR19), .B(_02470__PTR3), .S(_02435__PTR2), .Z(_02678__PTR83) );
  MUX2_X1 U10028 ( .A(P3_EBX_PTR20), .B(_02470__PTR4), .S(_02435__PTR2), .Z(_02678__PTR84) );
  MUX2_X1 U10029 ( .A(P3_EBX_PTR21), .B(_02470__PTR5), .S(_02435__PTR2), .Z(_02678__PTR85) );
  MUX2_X1 U10030 ( .A(P3_EBX_PTR22), .B(_02470__PTR6), .S(_02435__PTR2), .Z(_02678__PTR86) );
  MUX2_X1 U10031 ( .A(P3_EBX_PTR23), .B(_03305__PTR0), .S(_02435__PTR2), .Z(_02678__PTR87) );
  MUX2_X1 U10032 ( .A(P3_EBX_PTR24), .B(_03306__PTR1), .S(_02435__PTR2), .Z(_02678__PTR88) );
  MUX2_X1 U10033 ( .A(P3_EBX_PTR25), .B(_03306__PTR2), .S(_02435__PTR2), .Z(_02678__PTR89) );
  MUX2_X1 U10034 ( .A(P3_EBX_PTR26), .B(_03306__PTR3), .S(_02435__PTR2), .Z(_02678__PTR90) );
  MUX2_X1 U10035 ( .A(P3_EBX_PTR27), .B(_03306__PTR4), .S(_02435__PTR2), .Z(_02678__PTR91) );
  MUX2_X1 U10036 ( .A(P3_EBX_PTR28), .B(_03306__PTR5), .S(_02435__PTR2), .Z(_02678__PTR92) );
  MUX2_X1 U10037 ( .A(P3_EBX_PTR29), .B(_03306__PTR6), .S(_02435__PTR2), .Z(_02678__PTR93) );
  MUX2_X1 U10038 ( .A(P3_EBX_PTR30), .B(_03306__PTR7), .S(_02435__PTR2), .Z(_02678__PTR94) );
  MUX2_X1 U10039 ( .A(P3_EBX_PTR31), .B(_03304__PTR7), .S(_02435__PTR2), .Z(_02678__PTR95) );
  MUX2_X1 U10040 ( .A(P3_P1_InstQueueRd_Addr_PTR0), .B(_02465__PTR3), .S(_02435__PTR2), .Z(_02666__PTR25) );
  MUX2_X1 U10041 ( .A(P3_P1_InstQueueRd_Addr_PTR1), .B(_02465__PTR4), .S(_02435__PTR2), .Z(_02666__PTR26) );
  MUX2_X1 U10042 ( .A(P3_P1_InstQueueRd_Addr_PTR2), .B(_03310__PTR2), .S(_02435__PTR2), .Z(_02666__PTR27) );
  MUX2_X1 U10043 ( .A(P3_P1_InstQueueRd_Addr_PTR3), .B(_03310__PTR3), .S(_02435__PTR2), .Z(_02666__PTR28) );
  MUX2_X1 U10044 ( .A(P3_P1_InstQueueRd_Addr_PTR4), .B(1'b0), .S(_02435__PTR2), .Z(_02666__PTR29) );
  MUX2_X1 U10045 ( .A(P3_EAX_PTR0), .B(_02466__PTR0), .S(_02435__PTR2), .Z(_02674__PTR128) );
  MUX2_X1 U10046 ( .A(P3_EAX_PTR1), .B(_02466__PTR1), .S(_02435__PTR2), .Z(_02674__PTR129) );
  MUX2_X1 U10047 ( .A(P3_EAX_PTR2), .B(_02466__PTR2), .S(_02435__PTR2), .Z(_02674__PTR130) );
  MUX2_X1 U10048 ( .A(P3_EAX_PTR3), .B(_02466__PTR3), .S(_02435__PTR2), .Z(_02674__PTR131) );
  MUX2_X1 U10049 ( .A(P3_EAX_PTR4), .B(_02466__PTR4), .S(_02435__PTR2), .Z(_02674__PTR132) );
  MUX2_X1 U10050 ( .A(P3_EAX_PTR5), .B(_02466__PTR5), .S(_02435__PTR2), .Z(_02674__PTR133) );
  MUX2_X1 U10051 ( .A(P3_EAX_PTR6), .B(_02466__PTR6), .S(_02435__PTR2), .Z(_02674__PTR134) );
  MUX2_X1 U10052 ( .A(P3_EAX_PTR7), .B(_02466__PTR7), .S(_02435__PTR2), .Z(_02674__PTR135) );
  MUX2_X1 U10053 ( .A(P3_EAX_PTR8), .B(_02472__PTR0), .S(_02435__PTR2), .Z(_02674__PTR136) );
  MUX2_X1 U10054 ( .A(P3_EAX_PTR9), .B(_02472__PTR1), .S(_02435__PTR2), .Z(_02674__PTR137) );
  MUX2_X1 U10055 ( .A(P3_EAX_PTR10), .B(_02472__PTR2), .S(_02435__PTR2), .Z(_02674__PTR138) );
  MUX2_X1 U10056 ( .A(P3_EAX_PTR11), .B(_02472__PTR3), .S(_02435__PTR2), .Z(_02674__PTR139) );
  MUX2_X1 U10057 ( .A(P3_EAX_PTR12), .B(_02472__PTR4), .S(_02435__PTR2), .Z(_02674__PTR140) );
  MUX2_X1 U10058 ( .A(P3_EAX_PTR13), .B(_02472__PTR5), .S(_02435__PTR2), .Z(_02674__PTR141) );
  MUX2_X1 U10059 ( .A(P3_EAX_PTR14), .B(_02472__PTR6), .S(_02435__PTR2), .Z(_02674__PTR142) );
  MUX2_X1 U10060 ( .A(P3_EAX_PTR15), .B(_02472__PTR7), .S(_02435__PTR2), .Z(_02674__PTR143) );
  MUX2_X1 U10061 ( .A(P3_EAX_PTR16), .B(_02470__PTR0), .S(_02435__PTR2), .Z(_02674__PTR144) );
  MUX2_X1 U10062 ( .A(P3_EAX_PTR17), .B(_02470__PTR1), .S(_02435__PTR2), .Z(_02674__PTR145) );
  MUX2_X1 U10063 ( .A(P3_EAX_PTR18), .B(_02470__PTR2), .S(_02435__PTR2), .Z(_02674__PTR146) );
  MUX2_X1 U10064 ( .A(P3_EAX_PTR19), .B(_02470__PTR3), .S(_02435__PTR2), .Z(_02674__PTR147) );
  MUX2_X1 U10065 ( .A(P3_EAX_PTR20), .B(_02470__PTR4), .S(_02435__PTR2), .Z(_02674__PTR148) );
  MUX2_X1 U10066 ( .A(P3_EAX_PTR21), .B(_02470__PTR5), .S(_02435__PTR2), .Z(_02674__PTR149) );
  MUX2_X1 U10067 ( .A(P3_EAX_PTR22), .B(_02470__PTR6), .S(_02435__PTR2), .Z(_02674__PTR150) );
  MUX2_X1 U10068 ( .A(P3_EAX_PTR23), .B(_03305__PTR0), .S(_02435__PTR2), .Z(_02674__PTR151) );
  MUX2_X1 U10069 ( .A(P3_EAX_PTR24), .B(_03306__PTR1), .S(_02435__PTR2), .Z(_02674__PTR152) );
  MUX2_X1 U10070 ( .A(P3_EAX_PTR25), .B(_03306__PTR2), .S(_02435__PTR2), .Z(_02674__PTR153) );
  MUX2_X1 U10071 ( .A(P3_EAX_PTR26), .B(_03306__PTR3), .S(_02435__PTR2), .Z(_02674__PTR154) );
  MUX2_X1 U10072 ( .A(P3_EAX_PTR27), .B(_03306__PTR4), .S(_02435__PTR2), .Z(_02674__PTR155) );
  MUX2_X1 U10073 ( .A(P3_EAX_PTR28), .B(_03306__PTR5), .S(_02435__PTR2), .Z(_02674__PTR156) );
  MUX2_X1 U10074 ( .A(P3_EAX_PTR29), .B(_03306__PTR6), .S(_02435__PTR2), .Z(_02674__PTR157) );
  MUX2_X1 U10075 ( .A(P3_EAX_PTR30), .B(_03306__PTR7), .S(_02435__PTR2), .Z(_02674__PTR158) );
  MUX2_X1 U10076 ( .A(P3_EAX_PTR31), .B(_03304__PTR7), .S(_02435__PTR2), .Z(_02674__PTR159) );
  MUX2_X1 U10077 ( .A(P3_P1_PhyAddrPointer_PTR0), .B(_03299__PTR0), .S(_02435__PTR2), .Z(_02670__PTR32) );
  MUX2_X1 U10078 ( .A(P3_P1_PhyAddrPointer_PTR1), .B(_03300__PTR1), .S(_02435__PTR2), .Z(_02670__PTR33) );
  MUX2_X1 U10079 ( .A(P3_P1_PhyAddrPointer_PTR2), .B(_03300__PTR2), .S(_02435__PTR2), .Z(_02670__PTR34) );
  MUX2_X1 U10080 ( .A(P3_P1_PhyAddrPointer_PTR3), .B(_03300__PTR3), .S(_02435__PTR2), .Z(_02670__PTR35) );
  MUX2_X1 U10081 ( .A(P3_P1_PhyAddrPointer_PTR4), .B(_03300__PTR4), .S(_02435__PTR2), .Z(_02670__PTR36) );
  MUX2_X1 U10082 ( .A(P3_P1_PhyAddrPointer_PTR5), .B(_03300__PTR5), .S(_02435__PTR2), .Z(_02670__PTR37) );
  MUX2_X1 U10083 ( .A(P3_P1_PhyAddrPointer_PTR6), .B(_03300__PTR6), .S(_02435__PTR2), .Z(_02670__PTR38) );
  MUX2_X1 U10084 ( .A(P3_P1_PhyAddrPointer_PTR7), .B(_03300__PTR7), .S(_02435__PTR2), .Z(_02670__PTR39) );
  MUX2_X1 U10085 ( .A(P3_P1_PhyAddrPointer_PTR8), .B(_03300__PTR8), .S(_02435__PTR2), .Z(_02670__PTR40) );
  MUX2_X1 U10086 ( .A(P3_P1_PhyAddrPointer_PTR9), .B(_03300__PTR9), .S(_02435__PTR2), .Z(_02670__PTR41) );
  MUX2_X1 U10087 ( .A(P3_P1_PhyAddrPointer_PTR10), .B(_03300__PTR10), .S(_02435__PTR2), .Z(_02670__PTR42) );
  MUX2_X1 U10088 ( .A(P3_P1_PhyAddrPointer_PTR11), .B(_03300__PTR11), .S(_02435__PTR2), .Z(_02670__PTR43) );
  MUX2_X1 U10089 ( .A(P3_P1_PhyAddrPointer_PTR12), .B(_03300__PTR12), .S(_02435__PTR2), .Z(_02670__PTR44) );
  MUX2_X1 U10090 ( .A(P3_P1_PhyAddrPointer_PTR13), .B(_03300__PTR13), .S(_02435__PTR2), .Z(_02670__PTR45) );
  MUX2_X1 U10091 ( .A(P3_P1_PhyAddrPointer_PTR14), .B(_03300__PTR14), .S(_02435__PTR2), .Z(_02670__PTR46) );
  MUX2_X1 U10092 ( .A(P3_P1_PhyAddrPointer_PTR15), .B(_03300__PTR15), .S(_02435__PTR2), .Z(_02670__PTR47) );
  MUX2_X1 U10093 ( .A(P3_P1_PhyAddrPointer_PTR16), .B(_03300__PTR16), .S(_02435__PTR2), .Z(_02670__PTR48) );
  MUX2_X1 U10094 ( .A(P3_P1_PhyAddrPointer_PTR17), .B(_03300__PTR17), .S(_02435__PTR2), .Z(_02670__PTR49) );
  MUX2_X1 U10095 ( .A(P3_P1_PhyAddrPointer_PTR18), .B(_03300__PTR18), .S(_02435__PTR2), .Z(_02670__PTR50) );
  MUX2_X1 U10096 ( .A(P3_P1_PhyAddrPointer_PTR19), .B(_03300__PTR19), .S(_02435__PTR2), .Z(_02670__PTR51) );
  MUX2_X1 U10097 ( .A(P3_P1_PhyAddrPointer_PTR20), .B(_03300__PTR20), .S(_02435__PTR2), .Z(_02670__PTR52) );
  MUX2_X1 U10098 ( .A(P3_P1_PhyAddrPointer_PTR21), .B(_03300__PTR21), .S(_02435__PTR2), .Z(_02670__PTR53) );
  MUX2_X1 U10099 ( .A(P3_P1_PhyAddrPointer_PTR22), .B(_03300__PTR22), .S(_02435__PTR2), .Z(_02670__PTR54) );
  MUX2_X1 U10100 ( .A(P3_P1_PhyAddrPointer_PTR23), .B(_03300__PTR23), .S(_02435__PTR2), .Z(_02670__PTR55) );
  MUX2_X1 U10101 ( .A(P3_P1_PhyAddrPointer_PTR24), .B(_03300__PTR24), .S(_02435__PTR2), .Z(_02670__PTR56) );
  MUX2_X1 U10102 ( .A(P3_P1_PhyAddrPointer_PTR25), .B(_03300__PTR25), .S(_02435__PTR2), .Z(_02670__PTR57) );
  MUX2_X1 U10103 ( .A(P3_P1_PhyAddrPointer_PTR26), .B(_03300__PTR26), .S(_02435__PTR2), .Z(_02670__PTR58) );
  MUX2_X1 U10104 ( .A(P3_P1_PhyAddrPointer_PTR27), .B(_03300__PTR27), .S(_02435__PTR2), .Z(_02670__PTR59) );
  MUX2_X1 U10105 ( .A(P3_P1_PhyAddrPointer_PTR28), .B(_03300__PTR28), .S(_02435__PTR2), .Z(_02670__PTR60) );
  MUX2_X1 U10106 ( .A(P3_P1_PhyAddrPointer_PTR29), .B(_03300__PTR29), .S(_02435__PTR2), .Z(_02670__PTR61) );
  MUX2_X1 U10107 ( .A(P3_P1_PhyAddrPointer_PTR30), .B(_03300__PTR30), .S(_02435__PTR2), .Z(_02670__PTR62) );
  MUX2_X1 U10108 ( .A(P3_P1_PhyAddrPointer_PTR31), .B(_03300__PTR31), .S(_02435__PTR2), .Z(_02670__PTR63) );
  MUX2_X1 U10109 ( .A(P3_P1_InstAddrPointer_PTR1), .B(_02616__PTR1), .S(_02585_), .Z(_02662__PTR65) );
  MUX2_X1 U10110 ( .A(P3_P1_InstAddrPointer_PTR2), .B(_02616__PTR2), .S(_02585_), .Z(_02662__PTR66) );
  MUX2_X1 U10111 ( .A(P3_P1_InstAddrPointer_PTR3), .B(_02616__PTR3), .S(_02585_), .Z(_02662__PTR67) );
  MUX2_X1 U10112 ( .A(P3_P1_InstAddrPointer_PTR4), .B(_02616__PTR4), .S(_02585_), .Z(_02662__PTR68) );
  MUX2_X1 U10113 ( .A(P3_P1_InstAddrPointer_PTR5), .B(_02616__PTR5), .S(_02585_), .Z(_02662__PTR69) );
  MUX2_X1 U10114 ( .A(P3_P1_InstAddrPointer_PTR6), .B(_02616__PTR6), .S(_02585_), .Z(_02662__PTR70) );
  MUX2_X1 U10115 ( .A(P3_P1_InstAddrPointer_PTR7), .B(_02616__PTR7), .S(_02585_), .Z(_02662__PTR71) );
  MUX2_X1 U10116 ( .A(P3_P1_InstAddrPointer_PTR8), .B(_02616__PTR8), .S(_02585_), .Z(_02662__PTR72) );
  MUX2_X1 U10117 ( .A(P3_P1_InstAddrPointer_PTR9), .B(_02616__PTR9), .S(_02585_), .Z(_02662__PTR73) );
  MUX2_X1 U10118 ( .A(P3_P1_InstAddrPointer_PTR10), .B(_02616__PTR10), .S(_02585_), .Z(_02662__PTR74) );
  MUX2_X1 U10119 ( .A(P3_P1_InstAddrPointer_PTR11), .B(_02616__PTR11), .S(_02585_), .Z(_02662__PTR75) );
  MUX2_X1 U10120 ( .A(P3_P1_InstAddrPointer_PTR12), .B(_02616__PTR12), .S(_02585_), .Z(_02662__PTR76) );
  MUX2_X1 U10121 ( .A(P3_P1_InstAddrPointer_PTR13), .B(_02616__PTR13), .S(_02585_), .Z(_02662__PTR77) );
  MUX2_X1 U10122 ( .A(P3_P1_InstAddrPointer_PTR14), .B(_02616__PTR14), .S(_02585_), .Z(_02662__PTR78) );
  MUX2_X1 U10123 ( .A(P3_P1_InstAddrPointer_PTR15), .B(_02616__PTR15), .S(_02585_), .Z(_02662__PTR79) );
  MUX2_X1 U10124 ( .A(P3_P1_InstAddrPointer_PTR16), .B(_02616__PTR16), .S(_02585_), .Z(_02662__PTR80) );
  MUX2_X1 U10125 ( .A(P3_P1_InstAddrPointer_PTR17), .B(_02616__PTR17), .S(_02585_), .Z(_02662__PTR81) );
  MUX2_X1 U10126 ( .A(P3_P1_InstAddrPointer_PTR18), .B(_02616__PTR18), .S(_02585_), .Z(_02662__PTR82) );
  MUX2_X1 U10127 ( .A(P3_P1_InstAddrPointer_PTR19), .B(_02616__PTR19), .S(_02585_), .Z(_02662__PTR83) );
  MUX2_X1 U10128 ( .A(P3_P1_InstAddrPointer_PTR20), .B(_02616__PTR20), .S(_02585_), .Z(_02662__PTR84) );
  MUX2_X1 U10129 ( .A(P3_P1_InstAddrPointer_PTR21), .B(_02616__PTR21), .S(_02585_), .Z(_02662__PTR85) );
  MUX2_X1 U10130 ( .A(P3_P1_InstAddrPointer_PTR22), .B(_02616__PTR22), .S(_02585_), .Z(_02662__PTR86) );
  MUX2_X1 U10131 ( .A(P3_P1_InstAddrPointer_PTR23), .B(_02616__PTR23), .S(_02585_), .Z(_02662__PTR87) );
  MUX2_X1 U10132 ( .A(P3_P1_InstAddrPointer_PTR24), .B(_02616__PTR24), .S(_02585_), .Z(_02662__PTR88) );
  MUX2_X1 U10133 ( .A(P3_P1_InstAddrPointer_PTR25), .B(_02616__PTR25), .S(_02585_), .Z(_02662__PTR89) );
  MUX2_X1 U10134 ( .A(P3_P1_InstAddrPointer_PTR26), .B(_02616__PTR26), .S(_02585_), .Z(_02662__PTR90) );
  MUX2_X1 U10135 ( .A(P3_P1_InstAddrPointer_PTR27), .B(_02616__PTR27), .S(_02585_), .Z(_02662__PTR91) );
  MUX2_X1 U10136 ( .A(P3_P1_InstAddrPointer_PTR28), .B(_02616__PTR28), .S(_02585_), .Z(_02662__PTR92) );
  MUX2_X1 U10137 ( .A(P3_P1_InstAddrPointer_PTR29), .B(_02616__PTR29), .S(_02585_), .Z(_02662__PTR93) );
  MUX2_X1 U10138 ( .A(P3_P1_InstAddrPointer_PTR30), .B(_02616__PTR30), .S(_02585_), .Z(_02662__PTR94) );
  MUX2_X1 U10139 ( .A(P3_P1_InstAddrPointer_PTR31), .B(_02616__PTR31), .S(_02585_), .Z(_02662__PTR95) );
  MUX2_X1 U10140 ( .A(P3_P1_InstAddrPointer_PTR1), .B(_02598__PTR1), .S(_02585_), .Z(_02662__PTR97) );
  MUX2_X1 U10141 ( .A(P3_P1_InstAddrPointer_PTR2), .B(_02598__PTR2), .S(_02585_), .Z(_02662__PTR98) );
  MUX2_X1 U10142 ( .A(P3_P1_InstAddrPointer_PTR3), .B(_02598__PTR3), .S(_02585_), .Z(_02662__PTR99) );
  MUX2_X1 U10143 ( .A(P3_P1_InstAddrPointer_PTR4), .B(_02598__PTR4), .S(_02585_), .Z(_02662__PTR100) );
  MUX2_X1 U10144 ( .A(P3_P1_InstAddrPointer_PTR5), .B(_02598__PTR5), .S(_02585_), .Z(_02662__PTR101) );
  MUX2_X1 U10145 ( .A(P3_P1_InstAddrPointer_PTR6), .B(_02598__PTR6), .S(_02585_), .Z(_02662__PTR102) );
  MUX2_X1 U10146 ( .A(P3_P1_InstAddrPointer_PTR7), .B(_02598__PTR7), .S(_02585_), .Z(_02662__PTR103) );
  MUX2_X1 U10147 ( .A(P3_P1_InstAddrPointer_PTR8), .B(_02598__PTR8), .S(_02585_), .Z(_02662__PTR104) );
  MUX2_X1 U10148 ( .A(P3_P1_InstAddrPointer_PTR9), .B(_02598__PTR9), .S(_02585_), .Z(_02662__PTR105) );
  MUX2_X1 U10149 ( .A(P3_P1_InstAddrPointer_PTR10), .B(_02598__PTR10), .S(_02585_), .Z(_02662__PTR106) );
  MUX2_X1 U10150 ( .A(P3_P1_InstAddrPointer_PTR11), .B(_02598__PTR11), .S(_02585_), .Z(_02662__PTR107) );
  MUX2_X1 U10151 ( .A(P3_P1_InstAddrPointer_PTR12), .B(_02598__PTR12), .S(_02585_), .Z(_02662__PTR108) );
  MUX2_X1 U10152 ( .A(P3_P1_InstAddrPointer_PTR13), .B(_02598__PTR13), .S(_02585_), .Z(_02662__PTR109) );
  MUX2_X1 U10153 ( .A(P3_P1_InstAddrPointer_PTR14), .B(_02598__PTR14), .S(_02585_), .Z(_02662__PTR110) );
  MUX2_X1 U10154 ( .A(P3_P1_InstAddrPointer_PTR15), .B(_02598__PTR15), .S(_02585_), .Z(_02662__PTR111) );
  MUX2_X1 U10155 ( .A(P3_P1_InstAddrPointer_PTR16), .B(_02598__PTR16), .S(_02585_), .Z(_02662__PTR112) );
  MUX2_X1 U10156 ( .A(P3_P1_InstAddrPointer_PTR17), .B(_02598__PTR17), .S(_02585_), .Z(_02662__PTR113) );
  MUX2_X1 U10157 ( .A(P3_P1_InstAddrPointer_PTR18), .B(_02598__PTR18), .S(_02585_), .Z(_02662__PTR114) );
  MUX2_X1 U10158 ( .A(P3_P1_InstAddrPointer_PTR19), .B(_02598__PTR19), .S(_02585_), .Z(_02662__PTR115) );
  MUX2_X1 U10159 ( .A(P3_P1_InstAddrPointer_PTR20), .B(_02598__PTR20), .S(_02585_), .Z(_02662__PTR116) );
  MUX2_X1 U10160 ( .A(P3_P1_InstAddrPointer_PTR21), .B(_02598__PTR21), .S(_02585_), .Z(_02662__PTR117) );
  MUX2_X1 U10161 ( .A(P3_P1_InstAddrPointer_PTR22), .B(_02598__PTR22), .S(_02585_), .Z(_02662__PTR118) );
  MUX2_X1 U10162 ( .A(P3_P1_InstAddrPointer_PTR23), .B(_02598__PTR23), .S(_02585_), .Z(_02662__PTR119) );
  MUX2_X1 U10163 ( .A(P3_P1_InstAddrPointer_PTR24), .B(_02598__PTR24), .S(_02585_), .Z(_02662__PTR120) );
  MUX2_X1 U10164 ( .A(P3_P1_InstAddrPointer_PTR25), .B(_02598__PTR25), .S(_02585_), .Z(_02662__PTR121) );
  MUX2_X1 U10165 ( .A(P3_P1_InstAddrPointer_PTR26), .B(_02598__PTR26), .S(_02585_), .Z(_02662__PTR122) );
  MUX2_X1 U10166 ( .A(P3_P1_InstAddrPointer_PTR27), .B(_02598__PTR27), .S(_02585_), .Z(_02662__PTR123) );
  MUX2_X1 U10167 ( .A(P3_P1_InstAddrPointer_PTR28), .B(_02598__PTR28), .S(_02585_), .Z(_02662__PTR124) );
  MUX2_X1 U10168 ( .A(P3_P1_InstAddrPointer_PTR29), .B(_02598__PTR29), .S(_02585_), .Z(_02662__PTR125) );
  MUX2_X1 U10169 ( .A(P3_P1_InstAddrPointer_PTR30), .B(_02598__PTR30), .S(_02585_), .Z(_02662__PTR126) );
  MUX2_X1 U10170 ( .A(P3_P1_InstAddrPointer_PTR31), .B(_02598__PTR31), .S(_02585_), .Z(_02662__PTR127) );
  MUX2_X1 U10171 ( .A(P3_P1_InstAddrPointer_PTR0), .B(_02579__PTR0), .S(_02435__PTR3), .Z(_02662__PTR192) );
  MUX2_X1 U10172 ( .A(P3_P1_InstAddrPointer_PTR1), .B(_02579__PTR1), .S(_02435__PTR3), .Z(_02662__PTR193) );
  MUX2_X1 U10173 ( .A(P3_P1_InstAddrPointer_PTR2), .B(_02579__PTR2), .S(_02435__PTR3), .Z(_02662__PTR194) );
  MUX2_X1 U10174 ( .A(P3_P1_InstAddrPointer_PTR3), .B(_02579__PTR3), .S(_02435__PTR3), .Z(_02662__PTR195) );
  MUX2_X1 U10175 ( .A(P3_P1_InstAddrPointer_PTR4), .B(_02579__PTR4), .S(_02435__PTR3), .Z(_02662__PTR196) );
  MUX2_X1 U10176 ( .A(P3_P1_InstAddrPointer_PTR5), .B(_02579__PTR5), .S(_02435__PTR3), .Z(_02662__PTR197) );
  MUX2_X1 U10177 ( .A(P3_P1_InstAddrPointer_PTR6), .B(_02579__PTR6), .S(_02435__PTR3), .Z(_02662__PTR198) );
  MUX2_X1 U10178 ( .A(P3_P1_InstAddrPointer_PTR7), .B(_02579__PTR7), .S(_02435__PTR3), .Z(_02662__PTR199) );
  MUX2_X1 U10179 ( .A(P3_P1_InstAddrPointer_PTR8), .B(_02579__PTR8), .S(_02435__PTR3), .Z(_02662__PTR200) );
  MUX2_X1 U10180 ( .A(P3_P1_InstAddrPointer_PTR9), .B(_02579__PTR9), .S(_02435__PTR3), .Z(_02662__PTR201) );
  MUX2_X1 U10181 ( .A(P3_P1_InstAddrPointer_PTR10), .B(_02579__PTR10), .S(_02435__PTR3), .Z(_02662__PTR202) );
  MUX2_X1 U10182 ( .A(P3_P1_InstAddrPointer_PTR11), .B(_02579__PTR11), .S(_02435__PTR3), .Z(_02662__PTR203) );
  MUX2_X1 U10183 ( .A(P3_P1_InstAddrPointer_PTR12), .B(_02579__PTR12), .S(_02435__PTR3), .Z(_02662__PTR204) );
  MUX2_X1 U10184 ( .A(P3_P1_InstAddrPointer_PTR13), .B(_02579__PTR13), .S(_02435__PTR3), .Z(_02662__PTR205) );
  MUX2_X1 U10185 ( .A(P3_P1_InstAddrPointer_PTR14), .B(_02579__PTR14), .S(_02435__PTR3), .Z(_02662__PTR206) );
  MUX2_X1 U10186 ( .A(P3_P1_InstAddrPointer_PTR15), .B(_02579__PTR15), .S(_02435__PTR3), .Z(_02662__PTR207) );
  MUX2_X1 U10187 ( .A(P3_P1_InstAddrPointer_PTR16), .B(_02579__PTR16), .S(_02435__PTR3), .Z(_02662__PTR208) );
  MUX2_X1 U10188 ( .A(P3_P1_InstAddrPointer_PTR17), .B(_02579__PTR17), .S(_02435__PTR3), .Z(_02662__PTR209) );
  MUX2_X1 U10189 ( .A(P3_P1_InstAddrPointer_PTR18), .B(_02579__PTR18), .S(_02435__PTR3), .Z(_02662__PTR210) );
  MUX2_X1 U10190 ( .A(P3_P1_InstAddrPointer_PTR19), .B(_02579__PTR19), .S(_02435__PTR3), .Z(_02662__PTR211) );
  MUX2_X1 U10191 ( .A(P3_P1_InstAddrPointer_PTR20), .B(_02579__PTR20), .S(_02435__PTR3), .Z(_02662__PTR212) );
  MUX2_X1 U10192 ( .A(P3_P1_InstAddrPointer_PTR21), .B(_02579__PTR21), .S(_02435__PTR3), .Z(_02662__PTR213) );
  MUX2_X1 U10193 ( .A(P3_P1_InstAddrPointer_PTR22), .B(_02579__PTR22), .S(_02435__PTR3), .Z(_02662__PTR214) );
  MUX2_X1 U10194 ( .A(P3_P1_InstAddrPointer_PTR23), .B(_02579__PTR23), .S(_02435__PTR3), .Z(_02662__PTR215) );
  MUX2_X1 U10195 ( .A(P3_P1_InstAddrPointer_PTR24), .B(_02579__PTR24), .S(_02435__PTR3), .Z(_02662__PTR216) );
  MUX2_X1 U10196 ( .A(P3_P1_InstAddrPointer_PTR25), .B(_02579__PTR25), .S(_02435__PTR3), .Z(_02662__PTR217) );
  MUX2_X1 U10197 ( .A(P3_P1_InstAddrPointer_PTR26), .B(_02579__PTR26), .S(_02435__PTR3), .Z(_02662__PTR218) );
  MUX2_X1 U10198 ( .A(P3_P1_InstAddrPointer_PTR27), .B(_02579__PTR27), .S(_02435__PTR3), .Z(_02662__PTR219) );
  MUX2_X1 U10199 ( .A(P3_P1_InstAddrPointer_PTR28), .B(_02579__PTR28), .S(_02435__PTR3), .Z(_02662__PTR220) );
  MUX2_X1 U10200 ( .A(P3_P1_InstAddrPointer_PTR29), .B(_02579__PTR29), .S(_02435__PTR3), .Z(_02662__PTR221) );
  MUX2_X1 U10201 ( .A(P3_P1_InstAddrPointer_PTR30), .B(_02579__PTR30), .S(_02435__PTR3), .Z(_02662__PTR222) );
  MUX2_X1 U10202 ( .A(P3_P1_InstAddrPointer_PTR31), .B(_02579__PTR31), .S(_02435__PTR3), .Z(_02662__PTR223) );
  MUX2_X1 U10203 ( .A(P3_P1_PhyAddrPointer_PTR0), .B(_02579__PTR0), .S(_02435__PTR3), .Z(_02670__PTR64) );
  MUX2_X1 U10204 ( .A(P3_P1_PhyAddrPointer_PTR1), .B(_02579__PTR1), .S(_02435__PTR3), .Z(_02670__PTR65) );
  MUX2_X1 U10205 ( .A(P3_P1_PhyAddrPointer_PTR2), .B(_02579__PTR2), .S(_02435__PTR3), .Z(_02670__PTR66) );
  MUX2_X1 U10206 ( .A(P3_P1_PhyAddrPointer_PTR3), .B(_02579__PTR3), .S(_02435__PTR3), .Z(_02670__PTR67) );
  MUX2_X1 U10207 ( .A(P3_P1_PhyAddrPointer_PTR4), .B(_02579__PTR4), .S(_02435__PTR3), .Z(_02670__PTR68) );
  MUX2_X1 U10208 ( .A(P3_P1_PhyAddrPointer_PTR5), .B(_02579__PTR5), .S(_02435__PTR3), .Z(_02670__PTR69) );
  MUX2_X1 U10209 ( .A(P3_P1_PhyAddrPointer_PTR6), .B(_02579__PTR6), .S(_02435__PTR3), .Z(_02670__PTR70) );
  MUX2_X1 U10210 ( .A(P3_P1_PhyAddrPointer_PTR7), .B(_02579__PTR7), .S(_02435__PTR3), .Z(_02670__PTR71) );
  MUX2_X1 U10211 ( .A(P3_P1_PhyAddrPointer_PTR8), .B(_02579__PTR8), .S(_02435__PTR3), .Z(_02670__PTR72) );
  MUX2_X1 U10212 ( .A(P3_P1_PhyAddrPointer_PTR9), .B(_02579__PTR9), .S(_02435__PTR3), .Z(_02670__PTR73) );
  MUX2_X1 U10213 ( .A(P3_P1_PhyAddrPointer_PTR10), .B(_02579__PTR10), .S(_02435__PTR3), .Z(_02670__PTR74) );
  MUX2_X1 U10214 ( .A(P3_P1_PhyAddrPointer_PTR11), .B(_02579__PTR11), .S(_02435__PTR3), .Z(_02670__PTR75) );
  MUX2_X1 U10215 ( .A(P3_P1_PhyAddrPointer_PTR12), .B(_02579__PTR12), .S(_02435__PTR3), .Z(_02670__PTR76) );
  MUX2_X1 U10216 ( .A(P3_P1_PhyAddrPointer_PTR13), .B(_02579__PTR13), .S(_02435__PTR3), .Z(_02670__PTR77) );
  MUX2_X1 U10217 ( .A(P3_P1_PhyAddrPointer_PTR14), .B(_02579__PTR14), .S(_02435__PTR3), .Z(_02670__PTR78) );
  MUX2_X1 U10218 ( .A(P3_P1_PhyAddrPointer_PTR15), .B(_02579__PTR15), .S(_02435__PTR3), .Z(_02670__PTR79) );
  MUX2_X1 U10219 ( .A(P3_P1_PhyAddrPointer_PTR16), .B(_02579__PTR16), .S(_02435__PTR3), .Z(_02670__PTR80) );
  MUX2_X1 U10220 ( .A(P3_P1_PhyAddrPointer_PTR17), .B(_02579__PTR17), .S(_02435__PTR3), .Z(_02670__PTR81) );
  MUX2_X1 U10221 ( .A(P3_P1_PhyAddrPointer_PTR18), .B(_02579__PTR18), .S(_02435__PTR3), .Z(_02670__PTR82) );
  MUX2_X1 U10222 ( .A(P3_P1_PhyAddrPointer_PTR19), .B(_02579__PTR19), .S(_02435__PTR3), .Z(_02670__PTR83) );
  MUX2_X1 U10223 ( .A(P3_P1_PhyAddrPointer_PTR20), .B(_02579__PTR20), .S(_02435__PTR3), .Z(_02670__PTR84) );
  MUX2_X1 U10224 ( .A(P3_P1_PhyAddrPointer_PTR21), .B(_02579__PTR21), .S(_02435__PTR3), .Z(_02670__PTR85) );
  MUX2_X1 U10225 ( .A(P3_P1_PhyAddrPointer_PTR22), .B(_02579__PTR22), .S(_02435__PTR3), .Z(_02670__PTR86) );
  MUX2_X1 U10226 ( .A(P3_P1_PhyAddrPointer_PTR23), .B(_02579__PTR23), .S(_02435__PTR3), .Z(_02670__PTR87) );
  MUX2_X1 U10227 ( .A(P3_P1_PhyAddrPointer_PTR24), .B(_02579__PTR24), .S(_02435__PTR3), .Z(_02670__PTR88) );
  MUX2_X1 U10228 ( .A(P3_P1_PhyAddrPointer_PTR25), .B(_02579__PTR25), .S(_02435__PTR3), .Z(_02670__PTR89) );
  MUX2_X1 U10229 ( .A(P3_P1_PhyAddrPointer_PTR26), .B(_02579__PTR26), .S(_02435__PTR3), .Z(_02670__PTR90) );
  MUX2_X1 U10230 ( .A(P3_P1_PhyAddrPointer_PTR27), .B(_02579__PTR27), .S(_02435__PTR3), .Z(_02670__PTR91) );
  MUX2_X1 U10231 ( .A(P3_P1_PhyAddrPointer_PTR28), .B(_02579__PTR28), .S(_02435__PTR3), .Z(_02670__PTR92) );
  MUX2_X1 U10232 ( .A(P3_P1_PhyAddrPointer_PTR29), .B(_02579__PTR29), .S(_02435__PTR3), .Z(_02670__PTR93) );
  MUX2_X1 U10233 ( .A(P3_P1_PhyAddrPointer_PTR30), .B(_02579__PTR30), .S(_02435__PTR3), .Z(_02670__PTR94) );
  MUX2_X1 U10234 ( .A(P3_P1_PhyAddrPointer_PTR31), .B(_02579__PTR31), .S(_02435__PTR3), .Z(_02670__PTR95) );
  MUX2_X1 U10235 ( .A(_03429__PTR0), .B(_03293__PTR0), .S(_03214__PTR7), .Z(_02579__PTR0) );
  MUX2_X1 U10236 ( .A(_03429__PTR1), .B(_03294__PTR1), .S(_03214__PTR7), .Z(_02579__PTR1) );
  MUX2_X1 U10237 ( .A(_03429__PTR2), .B(_03294__PTR2), .S(_03214__PTR7), .Z(_02579__PTR2) );
  MUX2_X1 U10238 ( .A(_03429__PTR3), .B(_03294__PTR3), .S(_03214__PTR7), .Z(_02579__PTR3) );
  MUX2_X1 U10239 ( .A(_03429__PTR4), .B(_03294__PTR4), .S(_03214__PTR7), .Z(_02579__PTR4) );
  MUX2_X1 U10240 ( .A(_03429__PTR5), .B(_03294__PTR5), .S(_03214__PTR7), .Z(_02579__PTR5) );
  MUX2_X1 U10241 ( .A(_03429__PTR6), .B(_03294__PTR6), .S(_03214__PTR7), .Z(_02579__PTR6) );
  MUX2_X1 U10242 ( .A(_03429__PTR7), .B(_03294__PTR7), .S(_03214__PTR7), .Z(_02579__PTR7) );
  MUX2_X1 U10243 ( .A(_03429__PTR8), .B(_03294__PTR8), .S(_03214__PTR7), .Z(_02579__PTR8) );
  MUX2_X1 U10244 ( .A(_03429__PTR9), .B(_03294__PTR9), .S(_03214__PTR7), .Z(_02579__PTR9) );
  MUX2_X1 U10245 ( .A(_03429__PTR10), .B(_03294__PTR10), .S(_03214__PTR7), .Z(_02579__PTR10) );
  MUX2_X1 U10246 ( .A(_03429__PTR11), .B(_03294__PTR11), .S(_03214__PTR7), .Z(_02579__PTR11) );
  MUX2_X1 U10247 ( .A(_03429__PTR12), .B(_03294__PTR12), .S(_03214__PTR7), .Z(_02579__PTR12) );
  MUX2_X1 U10248 ( .A(_03429__PTR13), .B(_03294__PTR13), .S(_03214__PTR7), .Z(_02579__PTR13) );
  MUX2_X1 U10249 ( .A(_03429__PTR14), .B(_03294__PTR14), .S(_03214__PTR7), .Z(_02579__PTR14) );
  MUX2_X1 U10250 ( .A(_03429__PTR15), .B(_03294__PTR15), .S(_03214__PTR7), .Z(_02579__PTR15) );
  MUX2_X1 U10251 ( .A(_03429__PTR16), .B(_03294__PTR16), .S(_03214__PTR7), .Z(_02579__PTR16) );
  MUX2_X1 U10252 ( .A(_03429__PTR17), .B(_03294__PTR17), .S(_03214__PTR7), .Z(_02579__PTR17) );
  MUX2_X1 U10253 ( .A(_03429__PTR18), .B(_03294__PTR18), .S(_03214__PTR7), .Z(_02579__PTR18) );
  MUX2_X1 U10254 ( .A(_03429__PTR19), .B(_03294__PTR19), .S(_03214__PTR7), .Z(_02579__PTR19) );
  MUX2_X1 U10255 ( .A(_03429__PTR20), .B(_03294__PTR20), .S(_03214__PTR7), .Z(_02579__PTR20) );
  MUX2_X1 U10256 ( .A(_03429__PTR21), .B(_03294__PTR21), .S(_03214__PTR7), .Z(_02579__PTR21) );
  MUX2_X1 U10257 ( .A(_03429__PTR22), .B(_03294__PTR22), .S(_03214__PTR7), .Z(_02579__PTR22) );
  MUX2_X1 U10258 ( .A(_03429__PTR23), .B(_03294__PTR23), .S(_03214__PTR7), .Z(_02579__PTR23) );
  MUX2_X1 U10259 ( .A(_03429__PTR24), .B(_03294__PTR24), .S(_03214__PTR7), .Z(_02579__PTR24) );
  MUX2_X1 U10260 ( .A(_03429__PTR25), .B(_03294__PTR25), .S(_03214__PTR7), .Z(_02579__PTR25) );
  MUX2_X1 U10261 ( .A(_03429__PTR26), .B(_03294__PTR26), .S(_03214__PTR7), .Z(_02579__PTR26) );
  MUX2_X1 U10262 ( .A(_03429__PTR27), .B(_03294__PTR27), .S(_03214__PTR7), .Z(_02579__PTR27) );
  MUX2_X1 U10263 ( .A(_03429__PTR28), .B(_03294__PTR28), .S(_03214__PTR7), .Z(_02579__PTR28) );
  MUX2_X1 U10264 ( .A(_03429__PTR29), .B(_03294__PTR29), .S(_03214__PTR7), .Z(_02579__PTR29) );
  MUX2_X1 U10265 ( .A(_03429__PTR30), .B(_03294__PTR30), .S(_03214__PTR7), .Z(_02579__PTR30) );
  MUX2_X1 U10266 ( .A(_03429__PTR31), .B(_03294__PTR31), .S(_03214__PTR7), .Z(_02579__PTR31) );
  MUX2_X1 U10267 ( .A(P3_P1_PhyAddrPointer_PTR0), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR128) );
  MUX2_X1 U10268 ( .A(_02577__PTR1), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR129) );
  MUX2_X1 U10269 ( .A(_02577__PTR2), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR130) );
  MUX2_X1 U10270 ( .A(_02577__PTR3), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR131) );
  MUX2_X1 U10271 ( .A(_02577__PTR4), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR132) );
  MUX2_X1 U10272 ( .A(_02577__PTR5), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR133) );
  MUX2_X1 U10273 ( .A(_02577__PTR6), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR134) );
  MUX2_X1 U10274 ( .A(_02577__PTR7), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR135) );
  MUX2_X1 U10275 ( .A(_02577__PTR8), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR136) );
  MUX2_X1 U10276 ( .A(_02577__PTR9), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR137) );
  MUX2_X1 U10277 ( .A(_02577__PTR10), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR138) );
  MUX2_X1 U10278 ( .A(_02577__PTR11), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR139) );
  MUX2_X1 U10279 ( .A(_02577__PTR12), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR140) );
  MUX2_X1 U10280 ( .A(_02577__PTR13), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR141) );
  MUX2_X1 U10281 ( .A(_02577__PTR14), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR142) );
  MUX2_X1 U10282 ( .A(_02577__PTR15), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR143) );
  MUX2_X1 U10283 ( .A(_02577__PTR16), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR144) );
  MUX2_X1 U10284 ( .A(_02577__PTR17), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR145) );
  MUX2_X1 U10285 ( .A(_02577__PTR18), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR146) );
  MUX2_X1 U10286 ( .A(_02577__PTR19), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR147) );
  MUX2_X1 U10287 ( .A(_02577__PTR20), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR148) );
  MUX2_X1 U10288 ( .A(_02577__PTR21), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR149) );
  MUX2_X1 U10289 ( .A(_02577__PTR22), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR150) );
  MUX2_X1 U10290 ( .A(_02577__PTR23), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR151) );
  MUX2_X1 U10291 ( .A(_02577__PTR24), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR152) );
  MUX2_X1 U10292 ( .A(_02577__PTR25), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR153) );
  MUX2_X1 U10293 ( .A(_02577__PTR26), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR154) );
  MUX2_X1 U10294 ( .A(_02577__PTR27), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR155) );
  MUX2_X1 U10295 ( .A(_02577__PTR28), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR156) );
  MUX2_X1 U10296 ( .A(_02577__PTR29), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR157) );
  MUX2_X1 U10297 ( .A(_02577__PTR30), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR158) );
  MUX2_X1 U10298 ( .A(_02577__PTR31), .B(1'b0), .S(P3_StateBS16), .Z(_02477__PTR160) );
  MUX2_X1 U10299 ( .A(_02473__PTR129), .B(1'b0), .S(P3_StateBS16), .Z(_02473__PTR65) );
  MUX2_X1 U10300 ( .A(_02473__PTR130), .B(_03285__PTR0), .S(P3_StateBS16), .Z(_02473__PTR66) );
  MUX2_X1 U10301 ( .A(_02473__PTR131), .B(_03286__PTR1), .S(P3_StateBS16), .Z(_02473__PTR67) );
  MUX2_X1 U10302 ( .A(_02473__PTR132), .B(_03286__PTR2), .S(P3_StateBS16), .Z(_02473__PTR68) );
  MUX2_X1 U10303 ( .A(_02473__PTR133), .B(_03286__PTR3), .S(P3_StateBS16), .Z(_02473__PTR69) );
  MUX2_X1 U10304 ( .A(_02473__PTR134), .B(_03286__PTR4), .S(P3_StateBS16), .Z(_02473__PTR70) );
  MUX2_X1 U10305 ( .A(_02473__PTR135), .B(_03286__PTR5), .S(P3_StateBS16), .Z(_02473__PTR71) );
  MUX2_X1 U10306 ( .A(_02473__PTR136), .B(_03286__PTR6), .S(P3_StateBS16), .Z(_02473__PTR72) );
  MUX2_X1 U10307 ( .A(_02473__PTR137), .B(_03286__PTR7), .S(P3_StateBS16), .Z(_02473__PTR73) );
  MUX2_X1 U10308 ( .A(_02473__PTR138), .B(_03286__PTR8), .S(P3_StateBS16), .Z(_02473__PTR74) );
  MUX2_X1 U10309 ( .A(_02473__PTR139), .B(_03286__PTR9), .S(P3_StateBS16), .Z(_02473__PTR75) );
  MUX2_X1 U10310 ( .A(_02473__PTR140), .B(_03286__PTR10), .S(P3_StateBS16), .Z(_02473__PTR76) );
  MUX2_X1 U10311 ( .A(_02473__PTR141), .B(_03286__PTR11), .S(P3_StateBS16), .Z(_02473__PTR77) );
  MUX2_X1 U10312 ( .A(_02473__PTR142), .B(_03286__PTR12), .S(P3_StateBS16), .Z(_02473__PTR78) );
  MUX2_X1 U10313 ( .A(_02473__PTR143), .B(_03286__PTR13), .S(P3_StateBS16), .Z(_02473__PTR79) );
  MUX2_X1 U10314 ( .A(_02473__PTR144), .B(_03286__PTR14), .S(P3_StateBS16), .Z(_02473__PTR80) );
  MUX2_X1 U10315 ( .A(_02473__PTR145), .B(_03286__PTR15), .S(P3_StateBS16), .Z(_02473__PTR81) );
  MUX2_X1 U10316 ( .A(_02473__PTR146), .B(_03286__PTR16), .S(P3_StateBS16), .Z(_02473__PTR82) );
  MUX2_X1 U10317 ( .A(_02473__PTR147), .B(_03286__PTR17), .S(P3_StateBS16), .Z(_02473__PTR83) );
  MUX2_X1 U10318 ( .A(_02473__PTR148), .B(_03286__PTR18), .S(P3_StateBS16), .Z(_02473__PTR84) );
  MUX2_X1 U10319 ( .A(_02473__PTR149), .B(_03286__PTR19), .S(P3_StateBS16), .Z(_02473__PTR85) );
  MUX2_X1 U10320 ( .A(_02473__PTR150), .B(_03286__PTR20), .S(P3_StateBS16), .Z(_02473__PTR86) );
  MUX2_X1 U10321 ( .A(_02473__PTR151), .B(_03286__PTR21), .S(P3_StateBS16), .Z(_02473__PTR87) );
  MUX2_X1 U10322 ( .A(_02473__PTR152), .B(_03286__PTR22), .S(P3_StateBS16), .Z(_02473__PTR88) );
  MUX2_X1 U10323 ( .A(_02473__PTR153), .B(_03286__PTR23), .S(P3_StateBS16), .Z(_02473__PTR89) );
  MUX2_X1 U10324 ( .A(_02473__PTR154), .B(_03286__PTR24), .S(P3_StateBS16), .Z(_02473__PTR90) );
  MUX2_X1 U10325 ( .A(_02473__PTR155), .B(_03286__PTR25), .S(P3_StateBS16), .Z(_02473__PTR91) );
  MUX2_X1 U10326 ( .A(_02473__PTR156), .B(_03286__PTR26), .S(P3_StateBS16), .Z(_02473__PTR92) );
  MUX2_X1 U10327 ( .A(_02473__PTR157), .B(_03286__PTR27), .S(P3_StateBS16), .Z(_02473__PTR93) );
  MUX2_X1 U10328 ( .A(_02473__PTR158), .B(_03286__PTR28), .S(P3_StateBS16), .Z(_02473__PTR94) );
  MUX2_X1 U10329 ( .A(_02473__PTR159), .B(_03286__PTR29), .S(P3_StateBS16), .Z(_02473__PTR95) );
  MUX2_X1 U10330 ( .A(_02420__PTR1), .B(_03281__PTR1), .S(P3_StateBS16), .Z(_02511__PTR17) );
  MUX2_X1 U10331 ( .A(_02420__PTR2), .B(_03281__PTR2), .S(P3_StateBS16), .Z(_02511__PTR18) );
  MUX2_X1 U10332 ( .A(_02420__PTR3), .B(_03281__PTR3), .S(P3_StateBS16), .Z(_02511__PTR19) );
  MUX2_X1 U10333 ( .A(_02509__PTR32), .B(_02576__PTR0), .S(P3_StateBS16), .Z(_02509__PTR16) );
  MUX2_X1 U10334 ( .A(_02509__PTR33), .B(_02576__PTR1), .S(P3_StateBS16), .Z(_02509__PTR17) );
  MUX2_X1 U10335 ( .A(_02509__PTR34), .B(_02576__PTR2), .S(P3_StateBS16), .Z(_02509__PTR18) );
  MUX2_X1 U10336 ( .A(_02509__PTR35), .B(_02576__PTR3), .S(P3_StateBS16), .Z(_02509__PTR19) );
  MUX2_X1 U10337 ( .A(_02509__PTR36), .B(_02576__PTR4), .S(P3_StateBS16), .Z(_02509__PTR20) );
  MUX2_X1 U10338 ( .A(_02509__PTR37), .B(_02576__PTR5), .S(P3_StateBS16), .Z(_02509__PTR21) );
  MUX2_X1 U10339 ( .A(_02509__PTR38), .B(_02576__PTR6), .S(P3_StateBS16), .Z(_02509__PTR22) );
  MUX2_X1 U10340 ( .A(_02509__PTR39), .B(_02576__PTR7), .S(P3_StateBS16), .Z(_02509__PTR23) );
  MUX2_X1 U10341 ( .A(_02507__PTR32), .B(_02575__PTR0), .S(P3_StateBS16), .Z(_02507__PTR16) );
  MUX2_X1 U10342 ( .A(_02507__PTR33), .B(_02575__PTR1), .S(P3_StateBS16), .Z(_02507__PTR17) );
  MUX2_X1 U10343 ( .A(_02507__PTR34), .B(_02575__PTR2), .S(P3_StateBS16), .Z(_02507__PTR18) );
  MUX2_X1 U10344 ( .A(_02507__PTR35), .B(_02575__PTR3), .S(P3_StateBS16), .Z(_02507__PTR19) );
  MUX2_X1 U10345 ( .A(_02507__PTR36), .B(_02575__PTR4), .S(P3_StateBS16), .Z(_02507__PTR20) );
  MUX2_X1 U10346 ( .A(_02507__PTR37), .B(_02575__PTR5), .S(P3_StateBS16), .Z(_02507__PTR21) );
  MUX2_X1 U10347 ( .A(_02507__PTR38), .B(_02575__PTR6), .S(P3_StateBS16), .Z(_02507__PTR22) );
  MUX2_X1 U10348 ( .A(_02507__PTR39), .B(_02575__PTR7), .S(P3_StateBS16), .Z(_02507__PTR23) );
  MUX2_X1 U10349 ( .A(_02505__PTR32), .B(_02574__PTR0), .S(P3_StateBS16), .Z(_02505__PTR16) );
  MUX2_X1 U10350 ( .A(_02505__PTR33), .B(_02574__PTR1), .S(P3_StateBS16), .Z(_02505__PTR17) );
  MUX2_X1 U10351 ( .A(_02505__PTR34), .B(_02574__PTR2), .S(P3_StateBS16), .Z(_02505__PTR18) );
  MUX2_X1 U10352 ( .A(_02505__PTR35), .B(_02574__PTR3), .S(P3_StateBS16), .Z(_02505__PTR19) );
  MUX2_X1 U10353 ( .A(_02505__PTR36), .B(_02574__PTR4), .S(P3_StateBS16), .Z(_02505__PTR20) );
  MUX2_X1 U10354 ( .A(_02505__PTR37), .B(_02574__PTR5), .S(P3_StateBS16), .Z(_02505__PTR21) );
  MUX2_X1 U10355 ( .A(_02505__PTR38), .B(_02574__PTR6), .S(P3_StateBS16), .Z(_02505__PTR22) );
  MUX2_X1 U10356 ( .A(_02505__PTR39), .B(_02574__PTR7), .S(P3_StateBS16), .Z(_02505__PTR23) );
  MUX2_X1 U10357 ( .A(_02503__PTR32), .B(_02573__PTR0), .S(P3_StateBS16), .Z(_02503__PTR16) );
  MUX2_X1 U10358 ( .A(_02503__PTR33), .B(_02573__PTR1), .S(P3_StateBS16), .Z(_02503__PTR17) );
  MUX2_X1 U10359 ( .A(_02503__PTR34), .B(_02573__PTR2), .S(P3_StateBS16), .Z(_02503__PTR18) );
  MUX2_X1 U10360 ( .A(_02503__PTR35), .B(_02573__PTR3), .S(P3_StateBS16), .Z(_02503__PTR19) );
  MUX2_X1 U10361 ( .A(_02503__PTR36), .B(_02573__PTR4), .S(P3_StateBS16), .Z(_02503__PTR20) );
  MUX2_X1 U10362 ( .A(_02503__PTR37), .B(_02573__PTR5), .S(P3_StateBS16), .Z(_02503__PTR21) );
  MUX2_X1 U10363 ( .A(_02503__PTR38), .B(_02573__PTR6), .S(P3_StateBS16), .Z(_02503__PTR22) );
  MUX2_X1 U10364 ( .A(_02503__PTR39), .B(_02573__PTR7), .S(P3_StateBS16), .Z(_02503__PTR23) );
  MUX2_X1 U10365 ( .A(_02501__PTR32), .B(_02572__PTR0), .S(P3_StateBS16), .Z(_02501__PTR16) );
  MUX2_X1 U10366 ( .A(_02501__PTR33), .B(_02572__PTR1), .S(P3_StateBS16), .Z(_02501__PTR17) );
  MUX2_X1 U10367 ( .A(_02501__PTR34), .B(_02572__PTR2), .S(P3_StateBS16), .Z(_02501__PTR18) );
  MUX2_X1 U10368 ( .A(_02501__PTR35), .B(_02572__PTR3), .S(P3_StateBS16), .Z(_02501__PTR19) );
  MUX2_X1 U10369 ( .A(_02501__PTR36), .B(_02572__PTR4), .S(P3_StateBS16), .Z(_02501__PTR20) );
  MUX2_X1 U10370 ( .A(_02501__PTR37), .B(_02572__PTR5), .S(P3_StateBS16), .Z(_02501__PTR21) );
  MUX2_X1 U10371 ( .A(_02501__PTR38), .B(_02572__PTR6), .S(P3_StateBS16), .Z(_02501__PTR22) );
  MUX2_X1 U10372 ( .A(_02501__PTR39), .B(_02572__PTR7), .S(P3_StateBS16), .Z(_02501__PTR23) );
  MUX2_X1 U10373 ( .A(_02499__PTR32), .B(_02571__PTR0), .S(P3_StateBS16), .Z(_02499__PTR16) );
  MUX2_X1 U10374 ( .A(_02499__PTR33), .B(_02571__PTR1), .S(P3_StateBS16), .Z(_02499__PTR17) );
  MUX2_X1 U10375 ( .A(_02499__PTR34), .B(_02571__PTR2), .S(P3_StateBS16), .Z(_02499__PTR18) );
  MUX2_X1 U10376 ( .A(_02499__PTR35), .B(_02571__PTR3), .S(P3_StateBS16), .Z(_02499__PTR19) );
  MUX2_X1 U10377 ( .A(_02499__PTR36), .B(_02571__PTR4), .S(P3_StateBS16), .Z(_02499__PTR20) );
  MUX2_X1 U10378 ( .A(_02499__PTR37), .B(_02571__PTR5), .S(P3_StateBS16), .Z(_02499__PTR21) );
  MUX2_X1 U10379 ( .A(_02499__PTR38), .B(_02571__PTR6), .S(P3_StateBS16), .Z(_02499__PTR22) );
  MUX2_X1 U10380 ( .A(_02499__PTR39), .B(_02571__PTR7), .S(P3_StateBS16), .Z(_02499__PTR23) );
  MUX2_X1 U10381 ( .A(_02497__PTR32), .B(_02570__PTR0), .S(P3_StateBS16), .Z(_02497__PTR16) );
  MUX2_X1 U10382 ( .A(_02497__PTR33), .B(_02570__PTR1), .S(P3_StateBS16), .Z(_02497__PTR17) );
  MUX2_X1 U10383 ( .A(_02497__PTR34), .B(_02570__PTR2), .S(P3_StateBS16), .Z(_02497__PTR18) );
  MUX2_X1 U10384 ( .A(_02497__PTR35), .B(_02570__PTR3), .S(P3_StateBS16), .Z(_02497__PTR19) );
  MUX2_X1 U10385 ( .A(_02497__PTR36), .B(_02570__PTR4), .S(P3_StateBS16), .Z(_02497__PTR20) );
  MUX2_X1 U10386 ( .A(_02497__PTR37), .B(_02570__PTR5), .S(P3_StateBS16), .Z(_02497__PTR21) );
  MUX2_X1 U10387 ( .A(_02497__PTR38), .B(_02570__PTR6), .S(P3_StateBS16), .Z(_02497__PTR22) );
  MUX2_X1 U10388 ( .A(_02497__PTR39), .B(_02570__PTR7), .S(P3_StateBS16), .Z(_02497__PTR23) );
  MUX2_X1 U10389 ( .A(_02495__PTR32), .B(_02569__PTR0), .S(P3_StateBS16), .Z(_02495__PTR16) );
  MUX2_X1 U10390 ( .A(_02495__PTR33), .B(_02569__PTR1), .S(P3_StateBS16), .Z(_02495__PTR17) );
  MUX2_X1 U10391 ( .A(_02495__PTR34), .B(_02569__PTR2), .S(P3_StateBS16), .Z(_02495__PTR18) );
  MUX2_X1 U10392 ( .A(_02495__PTR35), .B(_02569__PTR3), .S(P3_StateBS16), .Z(_02495__PTR19) );
  MUX2_X1 U10393 ( .A(_02495__PTR36), .B(_02569__PTR4), .S(P3_StateBS16), .Z(_02495__PTR20) );
  MUX2_X1 U10394 ( .A(_02495__PTR37), .B(_02569__PTR5), .S(P3_StateBS16), .Z(_02495__PTR21) );
  MUX2_X1 U10395 ( .A(_02495__PTR38), .B(_02569__PTR6), .S(P3_StateBS16), .Z(_02495__PTR22) );
  MUX2_X1 U10396 ( .A(_02495__PTR39), .B(_02569__PTR7), .S(P3_StateBS16), .Z(_02495__PTR23) );
  MUX2_X1 U10397 ( .A(_02493__PTR32), .B(_02568__PTR0), .S(P3_StateBS16), .Z(_02493__PTR16) );
  MUX2_X1 U10398 ( .A(_02493__PTR33), .B(_02568__PTR1), .S(P3_StateBS16), .Z(_02493__PTR17) );
  MUX2_X1 U10399 ( .A(_02493__PTR34), .B(_02568__PTR2), .S(P3_StateBS16), .Z(_02493__PTR18) );
  MUX2_X1 U10400 ( .A(_02493__PTR35), .B(_02568__PTR3), .S(P3_StateBS16), .Z(_02493__PTR19) );
  MUX2_X1 U10401 ( .A(_02493__PTR36), .B(_02568__PTR4), .S(P3_StateBS16), .Z(_02493__PTR20) );
  MUX2_X1 U10402 ( .A(_02493__PTR37), .B(_02568__PTR5), .S(P3_StateBS16), .Z(_02493__PTR21) );
  MUX2_X1 U10403 ( .A(_02493__PTR38), .B(_02568__PTR6), .S(P3_StateBS16), .Z(_02493__PTR22) );
  MUX2_X1 U10404 ( .A(_02493__PTR39), .B(_02568__PTR7), .S(P3_StateBS16), .Z(_02493__PTR23) );
  MUX2_X1 U10405 ( .A(_02491__PTR32), .B(_02567__PTR0), .S(P3_StateBS16), .Z(_02491__PTR16) );
  MUX2_X1 U10406 ( .A(_02491__PTR33), .B(_02567__PTR1), .S(P3_StateBS16), .Z(_02491__PTR17) );
  MUX2_X1 U10407 ( .A(_02491__PTR34), .B(_02567__PTR2), .S(P3_StateBS16), .Z(_02491__PTR18) );
  MUX2_X1 U10408 ( .A(_02491__PTR35), .B(_02567__PTR3), .S(P3_StateBS16), .Z(_02491__PTR19) );
  MUX2_X1 U10409 ( .A(_02491__PTR36), .B(_02567__PTR4), .S(P3_StateBS16), .Z(_02491__PTR20) );
  MUX2_X1 U10410 ( .A(_02491__PTR37), .B(_02567__PTR5), .S(P3_StateBS16), .Z(_02491__PTR21) );
  MUX2_X1 U10411 ( .A(_02491__PTR38), .B(_02567__PTR6), .S(P3_StateBS16), .Z(_02491__PTR22) );
  MUX2_X1 U10412 ( .A(_02491__PTR39), .B(_02567__PTR7), .S(P3_StateBS16), .Z(_02491__PTR23) );
  MUX2_X1 U10413 ( .A(_02489__PTR32), .B(_02566__PTR0), .S(P3_StateBS16), .Z(_02489__PTR16) );
  MUX2_X1 U10414 ( .A(_02489__PTR33), .B(_02566__PTR1), .S(P3_StateBS16), .Z(_02489__PTR17) );
  MUX2_X1 U10415 ( .A(_02489__PTR34), .B(_02566__PTR2), .S(P3_StateBS16), .Z(_02489__PTR18) );
  MUX2_X1 U10416 ( .A(_02489__PTR35), .B(_02566__PTR3), .S(P3_StateBS16), .Z(_02489__PTR19) );
  MUX2_X1 U10417 ( .A(_02489__PTR36), .B(_02566__PTR4), .S(P3_StateBS16), .Z(_02489__PTR20) );
  MUX2_X1 U10418 ( .A(_02489__PTR37), .B(_02566__PTR5), .S(P3_StateBS16), .Z(_02489__PTR21) );
  MUX2_X1 U10419 ( .A(_02489__PTR38), .B(_02566__PTR6), .S(P3_StateBS16), .Z(_02489__PTR22) );
  MUX2_X1 U10420 ( .A(_02489__PTR39), .B(_02566__PTR7), .S(P3_StateBS16), .Z(_02489__PTR23) );
  MUX2_X1 U10421 ( .A(_02487__PTR32), .B(_02565__PTR0), .S(P3_StateBS16), .Z(_02487__PTR16) );
  MUX2_X1 U10422 ( .A(_02487__PTR33), .B(_02565__PTR1), .S(P3_StateBS16), .Z(_02487__PTR17) );
  MUX2_X1 U10423 ( .A(_02487__PTR34), .B(_02565__PTR2), .S(P3_StateBS16), .Z(_02487__PTR18) );
  MUX2_X1 U10424 ( .A(_02487__PTR35), .B(_02565__PTR3), .S(P3_StateBS16), .Z(_02487__PTR19) );
  MUX2_X1 U10425 ( .A(_02487__PTR36), .B(_02565__PTR4), .S(P3_StateBS16), .Z(_02487__PTR20) );
  MUX2_X1 U10426 ( .A(_02487__PTR37), .B(_02565__PTR5), .S(P3_StateBS16), .Z(_02487__PTR21) );
  MUX2_X1 U10427 ( .A(_02487__PTR38), .B(_02565__PTR6), .S(P3_StateBS16), .Z(_02487__PTR22) );
  MUX2_X1 U10428 ( .A(_02487__PTR39), .B(_02565__PTR7), .S(P3_StateBS16), .Z(_02487__PTR23) );
  MUX2_X1 U10429 ( .A(_02485__PTR32), .B(_02564__PTR0), .S(P3_StateBS16), .Z(_02485__PTR16) );
  MUX2_X1 U10430 ( .A(_02485__PTR33), .B(_02564__PTR1), .S(P3_StateBS16), .Z(_02485__PTR17) );
  MUX2_X1 U10431 ( .A(_02485__PTR34), .B(_02564__PTR2), .S(P3_StateBS16), .Z(_02485__PTR18) );
  MUX2_X1 U10432 ( .A(_02485__PTR35), .B(_02564__PTR3), .S(P3_StateBS16), .Z(_02485__PTR19) );
  MUX2_X1 U10433 ( .A(_02485__PTR36), .B(_02564__PTR4), .S(P3_StateBS16), .Z(_02485__PTR20) );
  MUX2_X1 U10434 ( .A(_02485__PTR37), .B(_02564__PTR5), .S(P3_StateBS16), .Z(_02485__PTR21) );
  MUX2_X1 U10435 ( .A(_02485__PTR38), .B(_02564__PTR6), .S(P3_StateBS16), .Z(_02485__PTR22) );
  MUX2_X1 U10436 ( .A(_02485__PTR39), .B(_02564__PTR7), .S(P3_StateBS16), .Z(_02485__PTR23) );
  MUX2_X1 U10437 ( .A(_02483__PTR32), .B(_02563__PTR0), .S(P3_StateBS16), .Z(_02483__PTR16) );
  MUX2_X1 U10438 ( .A(_02483__PTR33), .B(_02563__PTR1), .S(P3_StateBS16), .Z(_02483__PTR17) );
  MUX2_X1 U10439 ( .A(_02483__PTR34), .B(_02563__PTR2), .S(P3_StateBS16), .Z(_02483__PTR18) );
  MUX2_X1 U10440 ( .A(_02483__PTR35), .B(_02563__PTR3), .S(P3_StateBS16), .Z(_02483__PTR19) );
  MUX2_X1 U10441 ( .A(_02483__PTR36), .B(_02563__PTR4), .S(P3_StateBS16), .Z(_02483__PTR20) );
  MUX2_X1 U10442 ( .A(_02483__PTR37), .B(_02563__PTR5), .S(P3_StateBS16), .Z(_02483__PTR21) );
  MUX2_X1 U10443 ( .A(_02483__PTR38), .B(_02563__PTR6), .S(P3_StateBS16), .Z(_02483__PTR22) );
  MUX2_X1 U10444 ( .A(_02483__PTR39), .B(_02563__PTR7), .S(P3_StateBS16), .Z(_02483__PTR23) );
  MUX2_X1 U10445 ( .A(_02481__PTR32), .B(_02562__PTR0), .S(P3_StateBS16), .Z(_02481__PTR16) );
  MUX2_X1 U10446 ( .A(_02481__PTR33), .B(_02562__PTR1), .S(P3_StateBS16), .Z(_02481__PTR17) );
  MUX2_X1 U10447 ( .A(_02481__PTR34), .B(_02562__PTR2), .S(P3_StateBS16), .Z(_02481__PTR18) );
  MUX2_X1 U10448 ( .A(_02481__PTR35), .B(_02562__PTR3), .S(P3_StateBS16), .Z(_02481__PTR19) );
  MUX2_X1 U10449 ( .A(_02481__PTR36), .B(_02562__PTR4), .S(P3_StateBS16), .Z(_02481__PTR20) );
  MUX2_X1 U10450 ( .A(_02481__PTR37), .B(_02562__PTR5), .S(P3_StateBS16), .Z(_02481__PTR21) );
  MUX2_X1 U10451 ( .A(_02481__PTR38), .B(_02562__PTR6), .S(P3_StateBS16), .Z(_02481__PTR22) );
  MUX2_X1 U10452 ( .A(_02481__PTR39), .B(_02562__PTR7), .S(P3_StateBS16), .Z(_02481__PTR23) );
  MUX2_X1 U10453 ( .A(_02479__PTR32), .B(_02561__PTR0), .S(P3_StateBS16), .Z(_02479__PTR16) );
  MUX2_X1 U10454 ( .A(_02479__PTR33), .B(_02561__PTR1), .S(P3_StateBS16), .Z(_02479__PTR17) );
  MUX2_X1 U10455 ( .A(_02479__PTR34), .B(_02561__PTR2), .S(P3_StateBS16), .Z(_02479__PTR18) );
  MUX2_X1 U10456 ( .A(_02479__PTR35), .B(_02561__PTR3), .S(P3_StateBS16), .Z(_02479__PTR19) );
  MUX2_X1 U10457 ( .A(_02479__PTR36), .B(_02561__PTR4), .S(P3_StateBS16), .Z(_02479__PTR20) );
  MUX2_X1 U10458 ( .A(_02479__PTR37), .B(_02561__PTR5), .S(P3_StateBS16), .Z(_02479__PTR21) );
  MUX2_X1 U10459 ( .A(_02479__PTR38), .B(_02561__PTR6), .S(P3_StateBS16), .Z(_02479__PTR22) );
  MUX2_X1 U10460 ( .A(_02479__PTR39), .B(_02561__PTR7), .S(P3_StateBS16), .Z(_02479__PTR23) );
  MUX2_X1 U10461 ( .A(_03436__PTR1), .B(_02473__PTR129), .S(_03204__PTR31), .Z(_02577__PTR1) );
  MUX2_X1 U10462 ( .A(_03436__PTR2), .B(_02473__PTR130), .S(_03204__PTR31), .Z(_02577__PTR2) );
  MUX2_X1 U10463 ( .A(_03436__PTR3), .B(_02473__PTR131), .S(_03204__PTR31), .Z(_02577__PTR3) );
  MUX2_X1 U10464 ( .A(_03436__PTR4), .B(_02473__PTR132), .S(_03204__PTR31), .Z(_02577__PTR4) );
  MUX2_X1 U10465 ( .A(_03436__PTR5), .B(_02473__PTR133), .S(_03204__PTR31), .Z(_02577__PTR5) );
  MUX2_X1 U10466 ( .A(_03436__PTR6), .B(_02473__PTR134), .S(_03204__PTR31), .Z(_02577__PTR6) );
  MUX2_X1 U10467 ( .A(_03436__PTR7), .B(_02473__PTR135), .S(_03204__PTR31), .Z(_02577__PTR7) );
  MUX2_X1 U10468 ( .A(_03436__PTR8), .B(_02473__PTR136), .S(_03204__PTR31), .Z(_02577__PTR8) );
  MUX2_X1 U10469 ( .A(_03436__PTR9), .B(_02473__PTR137), .S(_03204__PTR31), .Z(_02577__PTR9) );
  MUX2_X1 U10470 ( .A(_03436__PTR10), .B(_02473__PTR138), .S(_03204__PTR31), .Z(_02577__PTR10) );
  MUX2_X1 U10471 ( .A(_03436__PTR11), .B(_02473__PTR139), .S(_03204__PTR31), .Z(_02577__PTR11) );
  MUX2_X1 U10472 ( .A(_03436__PTR12), .B(_02473__PTR140), .S(_03204__PTR31), .Z(_02577__PTR12) );
  MUX2_X1 U10473 ( .A(_03436__PTR13), .B(_02473__PTR141), .S(_03204__PTR31), .Z(_02577__PTR13) );
  MUX2_X1 U10474 ( .A(_03436__PTR14), .B(_02473__PTR142), .S(_03204__PTR31), .Z(_02577__PTR14) );
  MUX2_X1 U10475 ( .A(_03436__PTR15), .B(_02473__PTR143), .S(_03204__PTR31), .Z(_02577__PTR15) );
  MUX2_X1 U10476 ( .A(_03436__PTR16), .B(_02473__PTR144), .S(_03204__PTR31), .Z(_02577__PTR16) );
  MUX2_X1 U10477 ( .A(_03436__PTR17), .B(_02473__PTR145), .S(_03204__PTR31), .Z(_02577__PTR17) );
  MUX2_X1 U10478 ( .A(_03436__PTR18), .B(_02473__PTR146), .S(_03204__PTR31), .Z(_02577__PTR18) );
  MUX2_X1 U10479 ( .A(_03436__PTR19), .B(_02473__PTR147), .S(_03204__PTR31), .Z(_02577__PTR19) );
  MUX2_X1 U10480 ( .A(_03436__PTR20), .B(_02473__PTR148), .S(_03204__PTR31), .Z(_02577__PTR20) );
  MUX2_X1 U10481 ( .A(_03436__PTR21), .B(_02473__PTR149), .S(_03204__PTR31), .Z(_02577__PTR21) );
  MUX2_X1 U10482 ( .A(_03436__PTR22), .B(_02473__PTR150), .S(_03204__PTR31), .Z(_02577__PTR22) );
  MUX2_X1 U10483 ( .A(_03436__PTR23), .B(_02473__PTR151), .S(_03204__PTR31), .Z(_02577__PTR23) );
  MUX2_X1 U10484 ( .A(_03436__PTR24), .B(_02473__PTR152), .S(_03204__PTR31), .Z(_02577__PTR24) );
  MUX2_X1 U10485 ( .A(_03436__PTR25), .B(_02473__PTR153), .S(_03204__PTR31), .Z(_02577__PTR25) );
  MUX2_X1 U10486 ( .A(_03436__PTR26), .B(_02473__PTR154), .S(_03204__PTR31), .Z(_02577__PTR26) );
  MUX2_X1 U10487 ( .A(_03436__PTR27), .B(_02473__PTR155), .S(_03204__PTR31), .Z(_02577__PTR27) );
  MUX2_X1 U10488 ( .A(_03436__PTR28), .B(_02473__PTR156), .S(_03204__PTR31), .Z(_02577__PTR28) );
  MUX2_X1 U10489 ( .A(_03436__PTR29), .B(_02473__PTR157), .S(_03204__PTR31), .Z(_02577__PTR29) );
  MUX2_X1 U10490 ( .A(_03436__PTR30), .B(_02473__PTR158), .S(_03204__PTR31), .Z(_02577__PTR30) );
  MUX2_X1 U10491 ( .A(_03436__PTR31), .B(_02473__PTR159), .S(_03204__PTR31), .Z(_02577__PTR31) );
  MUX2_X1 U10492 ( .A(_02559__PTR0), .B(_03278__PTR0), .S(_02423__PTR0), .Z(_02576__PTR0) );
  MUX2_X1 U10493 ( .A(_02559__PTR1), .B(_03279__PTR1), .S(_02423__PTR0), .Z(_02576__PTR1) );
  MUX2_X1 U10494 ( .A(_02559__PTR2), .B(_03279__PTR2), .S(_02423__PTR0), .Z(_02576__PTR2) );
  MUX2_X1 U10495 ( .A(_02559__PTR3), .B(_03279__PTR3), .S(_02423__PTR0), .Z(_02576__PTR3) );
  MUX2_X1 U10496 ( .A(_02559__PTR4), .B(_03279__PTR4), .S(_02423__PTR0), .Z(_02576__PTR4) );
  MUX2_X1 U10497 ( .A(_02559__PTR5), .B(_03279__PTR5), .S(_02423__PTR0), .Z(_02576__PTR5) );
  MUX2_X1 U10498 ( .A(_02559__PTR6), .B(_03279__PTR6), .S(_02423__PTR0), .Z(_02576__PTR6) );
  MUX2_X1 U10499 ( .A(_02559__PTR7), .B(_03279__PTR7), .S(_02423__PTR0), .Z(_02576__PTR7) );
  MUX2_X1 U10500 ( .A(_02558__PTR0), .B(_03278__PTR0), .S(_02423__PTR1), .Z(_02575__PTR0) );
  MUX2_X1 U10501 ( .A(_02558__PTR1), .B(_03279__PTR1), .S(_02423__PTR1), .Z(_02575__PTR1) );
  MUX2_X1 U10502 ( .A(_02558__PTR2), .B(_03279__PTR2), .S(_02423__PTR1), .Z(_02575__PTR2) );
  MUX2_X1 U10503 ( .A(_02558__PTR3), .B(_03279__PTR3), .S(_02423__PTR1), .Z(_02575__PTR3) );
  MUX2_X1 U10504 ( .A(_02558__PTR4), .B(_03279__PTR4), .S(_02423__PTR1), .Z(_02575__PTR4) );
  MUX2_X1 U10505 ( .A(_02558__PTR5), .B(_03279__PTR5), .S(_02423__PTR1), .Z(_02575__PTR5) );
  MUX2_X1 U10506 ( .A(_02558__PTR6), .B(_03279__PTR6), .S(_02423__PTR1), .Z(_02575__PTR6) );
  MUX2_X1 U10507 ( .A(_02558__PTR7), .B(_03279__PTR7), .S(_02423__PTR1), .Z(_02575__PTR7) );
  MUX2_X1 U10508 ( .A(_02557__PTR0), .B(_03278__PTR0), .S(_02423__PTR2), .Z(_02574__PTR0) );
  MUX2_X1 U10509 ( .A(_02557__PTR1), .B(_03279__PTR1), .S(_02423__PTR2), .Z(_02574__PTR1) );
  MUX2_X1 U10510 ( .A(_02557__PTR2), .B(_03279__PTR2), .S(_02423__PTR2), .Z(_02574__PTR2) );
  MUX2_X1 U10511 ( .A(_02557__PTR3), .B(_03279__PTR3), .S(_02423__PTR2), .Z(_02574__PTR3) );
  MUX2_X1 U10512 ( .A(_02557__PTR4), .B(_03279__PTR4), .S(_02423__PTR2), .Z(_02574__PTR4) );
  MUX2_X1 U10513 ( .A(_02557__PTR5), .B(_03279__PTR5), .S(_02423__PTR2), .Z(_02574__PTR5) );
  MUX2_X1 U10514 ( .A(_02557__PTR6), .B(_03279__PTR6), .S(_02423__PTR2), .Z(_02574__PTR6) );
  MUX2_X1 U10515 ( .A(_02557__PTR7), .B(_03279__PTR7), .S(_02423__PTR2), .Z(_02574__PTR7) );
  MUX2_X1 U10516 ( .A(_02556__PTR0), .B(_03278__PTR0), .S(_02423__PTR3), .Z(_02573__PTR0) );
  MUX2_X1 U10517 ( .A(_02556__PTR1), .B(_03279__PTR1), .S(_02423__PTR3), .Z(_02573__PTR1) );
  MUX2_X1 U10518 ( .A(_02556__PTR2), .B(_03279__PTR2), .S(_02423__PTR3), .Z(_02573__PTR2) );
  MUX2_X1 U10519 ( .A(_02556__PTR3), .B(_03279__PTR3), .S(_02423__PTR3), .Z(_02573__PTR3) );
  MUX2_X1 U10520 ( .A(_02556__PTR4), .B(_03279__PTR4), .S(_02423__PTR3), .Z(_02573__PTR4) );
  MUX2_X1 U10521 ( .A(_02556__PTR5), .B(_03279__PTR5), .S(_02423__PTR3), .Z(_02573__PTR5) );
  MUX2_X1 U10522 ( .A(_02556__PTR6), .B(_03279__PTR6), .S(_02423__PTR3), .Z(_02573__PTR6) );
  MUX2_X1 U10523 ( .A(_02556__PTR7), .B(_03279__PTR7), .S(_02423__PTR3), .Z(_02573__PTR7) );
  MUX2_X1 U10524 ( .A(_02555__PTR0), .B(_03278__PTR0), .S(_02423__PTR4), .Z(_02572__PTR0) );
  MUX2_X1 U10525 ( .A(_02555__PTR1), .B(_03279__PTR1), .S(_02423__PTR4), .Z(_02572__PTR1) );
  MUX2_X1 U10526 ( .A(_02555__PTR2), .B(_03279__PTR2), .S(_02423__PTR4), .Z(_02572__PTR2) );
  MUX2_X1 U10527 ( .A(_02555__PTR3), .B(_03279__PTR3), .S(_02423__PTR4), .Z(_02572__PTR3) );
  MUX2_X1 U10528 ( .A(_02555__PTR4), .B(_03279__PTR4), .S(_02423__PTR4), .Z(_02572__PTR4) );
  MUX2_X1 U10529 ( .A(_02555__PTR5), .B(_03279__PTR5), .S(_02423__PTR4), .Z(_02572__PTR5) );
  MUX2_X1 U10530 ( .A(_02555__PTR6), .B(_03279__PTR6), .S(_02423__PTR4), .Z(_02572__PTR6) );
  MUX2_X1 U10531 ( .A(_02555__PTR7), .B(_03279__PTR7), .S(_02423__PTR4), .Z(_02572__PTR7) );
  MUX2_X1 U10532 ( .A(_02554__PTR0), .B(_03278__PTR0), .S(_02423__PTR5), .Z(_02571__PTR0) );
  MUX2_X1 U10533 ( .A(_02554__PTR1), .B(_03279__PTR1), .S(_02423__PTR5), .Z(_02571__PTR1) );
  MUX2_X1 U10534 ( .A(_02554__PTR2), .B(_03279__PTR2), .S(_02423__PTR5), .Z(_02571__PTR2) );
  MUX2_X1 U10535 ( .A(_02554__PTR3), .B(_03279__PTR3), .S(_02423__PTR5), .Z(_02571__PTR3) );
  MUX2_X1 U10536 ( .A(_02554__PTR4), .B(_03279__PTR4), .S(_02423__PTR5), .Z(_02571__PTR4) );
  MUX2_X1 U10537 ( .A(_02554__PTR5), .B(_03279__PTR5), .S(_02423__PTR5), .Z(_02571__PTR5) );
  MUX2_X1 U10538 ( .A(_02554__PTR6), .B(_03279__PTR6), .S(_02423__PTR5), .Z(_02571__PTR6) );
  MUX2_X1 U10539 ( .A(_02554__PTR7), .B(_03279__PTR7), .S(_02423__PTR5), .Z(_02571__PTR7) );
  MUX2_X1 U10540 ( .A(_02553__PTR0), .B(_03278__PTR0), .S(_02423__PTR6), .Z(_02570__PTR0) );
  MUX2_X1 U10541 ( .A(_02553__PTR1), .B(_03279__PTR1), .S(_02423__PTR6), .Z(_02570__PTR1) );
  MUX2_X1 U10542 ( .A(_02553__PTR2), .B(_03279__PTR2), .S(_02423__PTR6), .Z(_02570__PTR2) );
  MUX2_X1 U10543 ( .A(_02553__PTR3), .B(_03279__PTR3), .S(_02423__PTR6), .Z(_02570__PTR3) );
  MUX2_X1 U10544 ( .A(_02553__PTR4), .B(_03279__PTR4), .S(_02423__PTR6), .Z(_02570__PTR4) );
  MUX2_X1 U10545 ( .A(_02553__PTR5), .B(_03279__PTR5), .S(_02423__PTR6), .Z(_02570__PTR5) );
  MUX2_X1 U10546 ( .A(_02553__PTR6), .B(_03279__PTR6), .S(_02423__PTR6), .Z(_02570__PTR6) );
  MUX2_X1 U10547 ( .A(_02553__PTR7), .B(_03279__PTR7), .S(_02423__PTR6), .Z(_02570__PTR7) );
  MUX2_X1 U10548 ( .A(_02552__PTR0), .B(_03278__PTR0), .S(_02423__PTR7), .Z(_02569__PTR0) );
  MUX2_X1 U10549 ( .A(_02552__PTR1), .B(_03279__PTR1), .S(_02423__PTR7), .Z(_02569__PTR1) );
  MUX2_X1 U10550 ( .A(_02552__PTR2), .B(_03279__PTR2), .S(_02423__PTR7), .Z(_02569__PTR2) );
  MUX2_X1 U10551 ( .A(_02552__PTR3), .B(_03279__PTR3), .S(_02423__PTR7), .Z(_02569__PTR3) );
  MUX2_X1 U10552 ( .A(_02552__PTR4), .B(_03279__PTR4), .S(_02423__PTR7), .Z(_02569__PTR4) );
  MUX2_X1 U10553 ( .A(_02552__PTR5), .B(_03279__PTR5), .S(_02423__PTR7), .Z(_02569__PTR5) );
  MUX2_X1 U10554 ( .A(_02552__PTR6), .B(_03279__PTR6), .S(_02423__PTR7), .Z(_02569__PTR6) );
  MUX2_X1 U10555 ( .A(_02552__PTR7), .B(_03279__PTR7), .S(_02423__PTR7), .Z(_02569__PTR7) );
  MUX2_X1 U10556 ( .A(_02551__PTR0), .B(_03278__PTR0), .S(_02423__PTR8), .Z(_02568__PTR0) );
  MUX2_X1 U10557 ( .A(_02551__PTR1), .B(_03279__PTR1), .S(_02423__PTR8), .Z(_02568__PTR1) );
  MUX2_X1 U10558 ( .A(_02551__PTR2), .B(_03279__PTR2), .S(_02423__PTR8), .Z(_02568__PTR2) );
  MUX2_X1 U10559 ( .A(_02551__PTR3), .B(_03279__PTR3), .S(_02423__PTR8), .Z(_02568__PTR3) );
  MUX2_X1 U10560 ( .A(_02551__PTR4), .B(_03279__PTR4), .S(_02423__PTR8), .Z(_02568__PTR4) );
  MUX2_X1 U10561 ( .A(_02551__PTR5), .B(_03279__PTR5), .S(_02423__PTR8), .Z(_02568__PTR5) );
  MUX2_X1 U10562 ( .A(_02551__PTR6), .B(_03279__PTR6), .S(_02423__PTR8), .Z(_02568__PTR6) );
  MUX2_X1 U10563 ( .A(_02551__PTR7), .B(_03279__PTR7), .S(_02423__PTR8), .Z(_02568__PTR7) );
  MUX2_X1 U10564 ( .A(_02550__PTR0), .B(_03278__PTR0), .S(_02423__PTR9), .Z(_02567__PTR0) );
  MUX2_X1 U10565 ( .A(_02550__PTR1), .B(_03279__PTR1), .S(_02423__PTR9), .Z(_02567__PTR1) );
  MUX2_X1 U10566 ( .A(_02550__PTR2), .B(_03279__PTR2), .S(_02423__PTR9), .Z(_02567__PTR2) );
  MUX2_X1 U10567 ( .A(_02550__PTR3), .B(_03279__PTR3), .S(_02423__PTR9), .Z(_02567__PTR3) );
  MUX2_X1 U10568 ( .A(_02550__PTR4), .B(_03279__PTR4), .S(_02423__PTR9), .Z(_02567__PTR4) );
  MUX2_X1 U10569 ( .A(_02550__PTR5), .B(_03279__PTR5), .S(_02423__PTR9), .Z(_02567__PTR5) );
  MUX2_X1 U10570 ( .A(_02550__PTR6), .B(_03279__PTR6), .S(_02423__PTR9), .Z(_02567__PTR6) );
  MUX2_X1 U10571 ( .A(_02550__PTR7), .B(_03279__PTR7), .S(_02423__PTR9), .Z(_02567__PTR7) );
  MUX2_X1 U10572 ( .A(_02549__PTR0), .B(_03278__PTR0), .S(_02423__PTR10), .Z(_02566__PTR0) );
  MUX2_X1 U10573 ( .A(_02549__PTR1), .B(_03279__PTR1), .S(_02423__PTR10), .Z(_02566__PTR1) );
  MUX2_X1 U10574 ( .A(_02549__PTR2), .B(_03279__PTR2), .S(_02423__PTR10), .Z(_02566__PTR2) );
  MUX2_X1 U10575 ( .A(_02549__PTR3), .B(_03279__PTR3), .S(_02423__PTR10), .Z(_02566__PTR3) );
  MUX2_X1 U10576 ( .A(_02549__PTR4), .B(_03279__PTR4), .S(_02423__PTR10), .Z(_02566__PTR4) );
  MUX2_X1 U10577 ( .A(_02549__PTR5), .B(_03279__PTR5), .S(_02423__PTR10), .Z(_02566__PTR5) );
  MUX2_X1 U10578 ( .A(_02549__PTR6), .B(_03279__PTR6), .S(_02423__PTR10), .Z(_02566__PTR6) );
  MUX2_X1 U10579 ( .A(_02549__PTR7), .B(_03279__PTR7), .S(_02423__PTR10), .Z(_02566__PTR7) );
  MUX2_X1 U10580 ( .A(_02548__PTR0), .B(_03278__PTR0), .S(_02423__PTR11), .Z(_02565__PTR0) );
  MUX2_X1 U10581 ( .A(_02548__PTR1), .B(_03279__PTR1), .S(_02423__PTR11), .Z(_02565__PTR1) );
  MUX2_X1 U10582 ( .A(_02548__PTR2), .B(_03279__PTR2), .S(_02423__PTR11), .Z(_02565__PTR2) );
  MUX2_X1 U10583 ( .A(_02548__PTR3), .B(_03279__PTR3), .S(_02423__PTR11), .Z(_02565__PTR3) );
  MUX2_X1 U10584 ( .A(_02548__PTR4), .B(_03279__PTR4), .S(_02423__PTR11), .Z(_02565__PTR4) );
  MUX2_X1 U10585 ( .A(_02548__PTR5), .B(_03279__PTR5), .S(_02423__PTR11), .Z(_02565__PTR5) );
  MUX2_X1 U10586 ( .A(_02548__PTR6), .B(_03279__PTR6), .S(_02423__PTR11), .Z(_02565__PTR6) );
  MUX2_X1 U10587 ( .A(_02548__PTR7), .B(_03279__PTR7), .S(_02423__PTR11), .Z(_02565__PTR7) );
  MUX2_X1 U10588 ( .A(_02547__PTR0), .B(_03278__PTR0), .S(_02423__PTR12), .Z(_02564__PTR0) );
  MUX2_X1 U10589 ( .A(_02547__PTR1), .B(_03279__PTR1), .S(_02423__PTR12), .Z(_02564__PTR1) );
  MUX2_X1 U10590 ( .A(_02547__PTR2), .B(_03279__PTR2), .S(_02423__PTR12), .Z(_02564__PTR2) );
  MUX2_X1 U10591 ( .A(_02547__PTR3), .B(_03279__PTR3), .S(_02423__PTR12), .Z(_02564__PTR3) );
  MUX2_X1 U10592 ( .A(_02547__PTR4), .B(_03279__PTR4), .S(_02423__PTR12), .Z(_02564__PTR4) );
  MUX2_X1 U10593 ( .A(_02547__PTR5), .B(_03279__PTR5), .S(_02423__PTR12), .Z(_02564__PTR5) );
  MUX2_X1 U10594 ( .A(_02547__PTR6), .B(_03279__PTR6), .S(_02423__PTR12), .Z(_02564__PTR6) );
  MUX2_X1 U10595 ( .A(_02547__PTR7), .B(_03279__PTR7), .S(_02423__PTR12), .Z(_02564__PTR7) );
  MUX2_X1 U10596 ( .A(_02546__PTR0), .B(_03278__PTR0), .S(_02423__PTR13), .Z(_02563__PTR0) );
  MUX2_X1 U10597 ( .A(_02546__PTR1), .B(_03279__PTR1), .S(_02423__PTR13), .Z(_02563__PTR1) );
  MUX2_X1 U10598 ( .A(_02546__PTR2), .B(_03279__PTR2), .S(_02423__PTR13), .Z(_02563__PTR2) );
  MUX2_X1 U10599 ( .A(_02546__PTR3), .B(_03279__PTR3), .S(_02423__PTR13), .Z(_02563__PTR3) );
  MUX2_X1 U10600 ( .A(_02546__PTR4), .B(_03279__PTR4), .S(_02423__PTR13), .Z(_02563__PTR4) );
  MUX2_X1 U10601 ( .A(_02546__PTR5), .B(_03279__PTR5), .S(_02423__PTR13), .Z(_02563__PTR5) );
  MUX2_X1 U10602 ( .A(_02546__PTR6), .B(_03279__PTR6), .S(_02423__PTR13), .Z(_02563__PTR6) );
  MUX2_X1 U10603 ( .A(_02546__PTR7), .B(_03279__PTR7), .S(_02423__PTR13), .Z(_02563__PTR7) );
  MUX2_X1 U10604 ( .A(_02545__PTR0), .B(_03278__PTR0), .S(_02423__PTR14), .Z(_02562__PTR0) );
  MUX2_X1 U10605 ( .A(_02545__PTR1), .B(_03279__PTR1), .S(_02423__PTR14), .Z(_02562__PTR1) );
  MUX2_X1 U10606 ( .A(_02545__PTR2), .B(_03279__PTR2), .S(_02423__PTR14), .Z(_02562__PTR2) );
  MUX2_X1 U10607 ( .A(_02545__PTR3), .B(_03279__PTR3), .S(_02423__PTR14), .Z(_02562__PTR3) );
  MUX2_X1 U10608 ( .A(_02545__PTR4), .B(_03279__PTR4), .S(_02423__PTR14), .Z(_02562__PTR4) );
  MUX2_X1 U10609 ( .A(_02545__PTR5), .B(_03279__PTR5), .S(_02423__PTR14), .Z(_02562__PTR5) );
  MUX2_X1 U10610 ( .A(_02545__PTR6), .B(_03279__PTR6), .S(_02423__PTR14), .Z(_02562__PTR6) );
  MUX2_X1 U10611 ( .A(_02545__PTR7), .B(_03279__PTR7), .S(_02423__PTR14), .Z(_02562__PTR7) );
  MUX2_X1 U10612 ( .A(_02544__PTR0), .B(_03278__PTR0), .S(_02423__PTR15), .Z(_02561__PTR0) );
  MUX2_X1 U10613 ( .A(_02544__PTR1), .B(_03279__PTR1), .S(_02423__PTR15), .Z(_02561__PTR1) );
  MUX2_X1 U10614 ( .A(_02544__PTR2), .B(_03279__PTR2), .S(_02423__PTR15), .Z(_02561__PTR2) );
  MUX2_X1 U10615 ( .A(_02544__PTR3), .B(_03279__PTR3), .S(_02423__PTR15), .Z(_02561__PTR3) );
  MUX2_X1 U10616 ( .A(_02544__PTR4), .B(_03279__PTR4), .S(_02423__PTR15), .Z(_02561__PTR4) );
  MUX2_X1 U10617 ( .A(_02544__PTR5), .B(_03279__PTR5), .S(_02423__PTR15), .Z(_02561__PTR5) );
  MUX2_X1 U10618 ( .A(_02544__PTR6), .B(_03279__PTR6), .S(_02423__PTR15), .Z(_02561__PTR6) );
  MUX2_X1 U10619 ( .A(_02544__PTR7), .B(_03279__PTR7), .S(_02423__PTR15), .Z(_02561__PTR7) );
  MUX2_X1 U10620 ( .A(_02509__PTR32), .B(_03273__PTR0), .S(_02421__PTR0), .Z(_02559__PTR0) );
  MUX2_X1 U10621 ( .A(_02509__PTR33), .B(_03274__PTR1), .S(_02421__PTR0), .Z(_02559__PTR1) );
  MUX2_X1 U10622 ( .A(_02509__PTR34), .B(_03274__PTR2), .S(_02421__PTR0), .Z(_02559__PTR2) );
  MUX2_X1 U10623 ( .A(_02509__PTR35), .B(_03274__PTR3), .S(_02421__PTR0), .Z(_02559__PTR3) );
  MUX2_X1 U10624 ( .A(_02509__PTR36), .B(_03274__PTR4), .S(_02421__PTR0), .Z(_02559__PTR4) );
  MUX2_X1 U10625 ( .A(_02509__PTR37), .B(_03274__PTR5), .S(_02421__PTR0), .Z(_02559__PTR5) );
  MUX2_X1 U10626 ( .A(_02509__PTR38), .B(_03274__PTR6), .S(_02421__PTR0), .Z(_02559__PTR6) );
  MUX2_X1 U10627 ( .A(_02509__PTR39), .B(_03274__PTR7), .S(_02421__PTR0), .Z(_02559__PTR7) );
  MUX2_X1 U10628 ( .A(_02507__PTR32), .B(_03273__PTR0), .S(_02421__PTR1), .Z(_02558__PTR0) );
  MUX2_X1 U10629 ( .A(_02507__PTR33), .B(_03274__PTR1), .S(_02421__PTR1), .Z(_02558__PTR1) );
  MUX2_X1 U10630 ( .A(_02507__PTR34), .B(_03274__PTR2), .S(_02421__PTR1), .Z(_02558__PTR2) );
  MUX2_X1 U10631 ( .A(_02507__PTR35), .B(_03274__PTR3), .S(_02421__PTR1), .Z(_02558__PTR3) );
  MUX2_X1 U10632 ( .A(_02507__PTR36), .B(_03274__PTR4), .S(_02421__PTR1), .Z(_02558__PTR4) );
  MUX2_X1 U10633 ( .A(_02507__PTR37), .B(_03274__PTR5), .S(_02421__PTR1), .Z(_02558__PTR5) );
  MUX2_X1 U10634 ( .A(_02507__PTR38), .B(_03274__PTR6), .S(_02421__PTR1), .Z(_02558__PTR6) );
  MUX2_X1 U10635 ( .A(_02507__PTR39), .B(_03274__PTR7), .S(_02421__PTR1), .Z(_02558__PTR7) );
  MUX2_X1 U10636 ( .A(_02505__PTR32), .B(_03273__PTR0), .S(_02421__PTR2), .Z(_02557__PTR0) );
  MUX2_X1 U10637 ( .A(_02505__PTR33), .B(_03274__PTR1), .S(_02421__PTR2), .Z(_02557__PTR1) );
  MUX2_X1 U10638 ( .A(_02505__PTR34), .B(_03274__PTR2), .S(_02421__PTR2), .Z(_02557__PTR2) );
  MUX2_X1 U10639 ( .A(_02505__PTR35), .B(_03274__PTR3), .S(_02421__PTR2), .Z(_02557__PTR3) );
  MUX2_X1 U10640 ( .A(_02505__PTR36), .B(_03274__PTR4), .S(_02421__PTR2), .Z(_02557__PTR4) );
  MUX2_X1 U10641 ( .A(_02505__PTR37), .B(_03274__PTR5), .S(_02421__PTR2), .Z(_02557__PTR5) );
  MUX2_X1 U10642 ( .A(_02505__PTR38), .B(_03274__PTR6), .S(_02421__PTR2), .Z(_02557__PTR6) );
  MUX2_X1 U10643 ( .A(_02505__PTR39), .B(_03274__PTR7), .S(_02421__PTR2), .Z(_02557__PTR7) );
  MUX2_X1 U10644 ( .A(_02503__PTR32), .B(_03273__PTR0), .S(_02421__PTR3), .Z(_02556__PTR0) );
  MUX2_X1 U10645 ( .A(_02503__PTR33), .B(_03274__PTR1), .S(_02421__PTR3), .Z(_02556__PTR1) );
  MUX2_X1 U10646 ( .A(_02503__PTR34), .B(_03274__PTR2), .S(_02421__PTR3), .Z(_02556__PTR2) );
  MUX2_X1 U10647 ( .A(_02503__PTR35), .B(_03274__PTR3), .S(_02421__PTR3), .Z(_02556__PTR3) );
  MUX2_X1 U10648 ( .A(_02503__PTR36), .B(_03274__PTR4), .S(_02421__PTR3), .Z(_02556__PTR4) );
  MUX2_X1 U10649 ( .A(_02503__PTR37), .B(_03274__PTR5), .S(_02421__PTR3), .Z(_02556__PTR5) );
  MUX2_X1 U10650 ( .A(_02503__PTR38), .B(_03274__PTR6), .S(_02421__PTR3), .Z(_02556__PTR6) );
  MUX2_X1 U10651 ( .A(_02503__PTR39), .B(_03274__PTR7), .S(_02421__PTR3), .Z(_02556__PTR7) );
  MUX2_X1 U10652 ( .A(_02501__PTR32), .B(_03273__PTR0), .S(_02421__PTR4), .Z(_02555__PTR0) );
  MUX2_X1 U10653 ( .A(_02501__PTR33), .B(_03274__PTR1), .S(_02421__PTR4), .Z(_02555__PTR1) );
  MUX2_X1 U10654 ( .A(_02501__PTR34), .B(_03274__PTR2), .S(_02421__PTR4), .Z(_02555__PTR2) );
  MUX2_X1 U10655 ( .A(_02501__PTR35), .B(_03274__PTR3), .S(_02421__PTR4), .Z(_02555__PTR3) );
  MUX2_X1 U10656 ( .A(_02501__PTR36), .B(_03274__PTR4), .S(_02421__PTR4), .Z(_02555__PTR4) );
  MUX2_X1 U10657 ( .A(_02501__PTR37), .B(_03274__PTR5), .S(_02421__PTR4), .Z(_02555__PTR5) );
  MUX2_X1 U10658 ( .A(_02501__PTR38), .B(_03274__PTR6), .S(_02421__PTR4), .Z(_02555__PTR6) );
  MUX2_X1 U10659 ( .A(_02501__PTR39), .B(_03274__PTR7), .S(_02421__PTR4), .Z(_02555__PTR7) );
  MUX2_X1 U10660 ( .A(_02499__PTR32), .B(_03273__PTR0), .S(_02421__PTR5), .Z(_02554__PTR0) );
  MUX2_X1 U10661 ( .A(_02499__PTR33), .B(_03274__PTR1), .S(_02421__PTR5), .Z(_02554__PTR1) );
  MUX2_X1 U10662 ( .A(_02499__PTR34), .B(_03274__PTR2), .S(_02421__PTR5), .Z(_02554__PTR2) );
  MUX2_X1 U10663 ( .A(_02499__PTR35), .B(_03274__PTR3), .S(_02421__PTR5), .Z(_02554__PTR3) );
  MUX2_X1 U10664 ( .A(_02499__PTR36), .B(_03274__PTR4), .S(_02421__PTR5), .Z(_02554__PTR4) );
  MUX2_X1 U10665 ( .A(_02499__PTR37), .B(_03274__PTR5), .S(_02421__PTR5), .Z(_02554__PTR5) );
  MUX2_X1 U10666 ( .A(_02499__PTR38), .B(_03274__PTR6), .S(_02421__PTR5), .Z(_02554__PTR6) );
  MUX2_X1 U10667 ( .A(_02499__PTR39), .B(_03274__PTR7), .S(_02421__PTR5), .Z(_02554__PTR7) );
  MUX2_X1 U10668 ( .A(_02497__PTR32), .B(_03273__PTR0), .S(_02421__PTR6), .Z(_02553__PTR0) );
  MUX2_X1 U10669 ( .A(_02497__PTR33), .B(_03274__PTR1), .S(_02421__PTR6), .Z(_02553__PTR1) );
  MUX2_X1 U10670 ( .A(_02497__PTR34), .B(_03274__PTR2), .S(_02421__PTR6), .Z(_02553__PTR2) );
  MUX2_X1 U10671 ( .A(_02497__PTR35), .B(_03274__PTR3), .S(_02421__PTR6), .Z(_02553__PTR3) );
  MUX2_X1 U10672 ( .A(_02497__PTR36), .B(_03274__PTR4), .S(_02421__PTR6), .Z(_02553__PTR4) );
  MUX2_X1 U10673 ( .A(_02497__PTR37), .B(_03274__PTR5), .S(_02421__PTR6), .Z(_02553__PTR5) );
  MUX2_X1 U10674 ( .A(_02497__PTR38), .B(_03274__PTR6), .S(_02421__PTR6), .Z(_02553__PTR6) );
  MUX2_X1 U10675 ( .A(_02497__PTR39), .B(_03274__PTR7), .S(_02421__PTR6), .Z(_02553__PTR7) );
  MUX2_X1 U10676 ( .A(_02495__PTR32), .B(_03273__PTR0), .S(_02421__PTR7), .Z(_02552__PTR0) );
  MUX2_X1 U10677 ( .A(_02495__PTR33), .B(_03274__PTR1), .S(_02421__PTR7), .Z(_02552__PTR1) );
  MUX2_X1 U10678 ( .A(_02495__PTR34), .B(_03274__PTR2), .S(_02421__PTR7), .Z(_02552__PTR2) );
  MUX2_X1 U10679 ( .A(_02495__PTR35), .B(_03274__PTR3), .S(_02421__PTR7), .Z(_02552__PTR3) );
  MUX2_X1 U10680 ( .A(_02495__PTR36), .B(_03274__PTR4), .S(_02421__PTR7), .Z(_02552__PTR4) );
  MUX2_X1 U10681 ( .A(_02495__PTR37), .B(_03274__PTR5), .S(_02421__PTR7), .Z(_02552__PTR5) );
  MUX2_X1 U10682 ( .A(_02495__PTR38), .B(_03274__PTR6), .S(_02421__PTR7), .Z(_02552__PTR6) );
  MUX2_X1 U10683 ( .A(_02495__PTR39), .B(_03274__PTR7), .S(_02421__PTR7), .Z(_02552__PTR7) );
  MUX2_X1 U10684 ( .A(_02493__PTR32), .B(_03273__PTR0), .S(_02421__PTR8), .Z(_02551__PTR0) );
  MUX2_X1 U10685 ( .A(_02493__PTR33), .B(_03274__PTR1), .S(_02421__PTR8), .Z(_02551__PTR1) );
  MUX2_X1 U10686 ( .A(_02493__PTR34), .B(_03274__PTR2), .S(_02421__PTR8), .Z(_02551__PTR2) );
  MUX2_X1 U10687 ( .A(_02493__PTR35), .B(_03274__PTR3), .S(_02421__PTR8), .Z(_02551__PTR3) );
  MUX2_X1 U10688 ( .A(_02493__PTR36), .B(_03274__PTR4), .S(_02421__PTR8), .Z(_02551__PTR4) );
  MUX2_X1 U10689 ( .A(_02493__PTR37), .B(_03274__PTR5), .S(_02421__PTR8), .Z(_02551__PTR5) );
  MUX2_X1 U10690 ( .A(_02493__PTR38), .B(_03274__PTR6), .S(_02421__PTR8), .Z(_02551__PTR6) );
  MUX2_X1 U10691 ( .A(_02493__PTR39), .B(_03274__PTR7), .S(_02421__PTR8), .Z(_02551__PTR7) );
  MUX2_X1 U10692 ( .A(_02491__PTR32), .B(_03273__PTR0), .S(_02421__PTR9), .Z(_02550__PTR0) );
  MUX2_X1 U10693 ( .A(_02491__PTR33), .B(_03274__PTR1), .S(_02421__PTR9), .Z(_02550__PTR1) );
  MUX2_X1 U10694 ( .A(_02491__PTR34), .B(_03274__PTR2), .S(_02421__PTR9), .Z(_02550__PTR2) );
  MUX2_X1 U10695 ( .A(_02491__PTR35), .B(_03274__PTR3), .S(_02421__PTR9), .Z(_02550__PTR3) );
  MUX2_X1 U10696 ( .A(_02491__PTR36), .B(_03274__PTR4), .S(_02421__PTR9), .Z(_02550__PTR4) );
  MUX2_X1 U10697 ( .A(_02491__PTR37), .B(_03274__PTR5), .S(_02421__PTR9), .Z(_02550__PTR5) );
  MUX2_X1 U10698 ( .A(_02491__PTR38), .B(_03274__PTR6), .S(_02421__PTR9), .Z(_02550__PTR6) );
  MUX2_X1 U10699 ( .A(_02491__PTR39), .B(_03274__PTR7), .S(_02421__PTR9), .Z(_02550__PTR7) );
  MUX2_X1 U10700 ( .A(_02489__PTR32), .B(_03273__PTR0), .S(_02421__PTR10), .Z(_02549__PTR0) );
  MUX2_X1 U10701 ( .A(_02489__PTR33), .B(_03274__PTR1), .S(_02421__PTR10), .Z(_02549__PTR1) );
  MUX2_X1 U10702 ( .A(_02489__PTR34), .B(_03274__PTR2), .S(_02421__PTR10), .Z(_02549__PTR2) );
  MUX2_X1 U10703 ( .A(_02489__PTR35), .B(_03274__PTR3), .S(_02421__PTR10), .Z(_02549__PTR3) );
  MUX2_X1 U10704 ( .A(_02489__PTR36), .B(_03274__PTR4), .S(_02421__PTR10), .Z(_02549__PTR4) );
  MUX2_X1 U10705 ( .A(_02489__PTR37), .B(_03274__PTR5), .S(_02421__PTR10), .Z(_02549__PTR5) );
  MUX2_X1 U10706 ( .A(_02489__PTR38), .B(_03274__PTR6), .S(_02421__PTR10), .Z(_02549__PTR6) );
  MUX2_X1 U10707 ( .A(_02489__PTR39), .B(_03274__PTR7), .S(_02421__PTR10), .Z(_02549__PTR7) );
  MUX2_X1 U10708 ( .A(_02487__PTR32), .B(_03273__PTR0), .S(_02421__PTR11), .Z(_02548__PTR0) );
  MUX2_X1 U10709 ( .A(_02487__PTR33), .B(_03274__PTR1), .S(_02421__PTR11), .Z(_02548__PTR1) );
  MUX2_X1 U10710 ( .A(_02487__PTR34), .B(_03274__PTR2), .S(_02421__PTR11), .Z(_02548__PTR2) );
  MUX2_X1 U10711 ( .A(_02487__PTR35), .B(_03274__PTR3), .S(_02421__PTR11), .Z(_02548__PTR3) );
  MUX2_X1 U10712 ( .A(_02487__PTR36), .B(_03274__PTR4), .S(_02421__PTR11), .Z(_02548__PTR4) );
  MUX2_X1 U10713 ( .A(_02487__PTR37), .B(_03274__PTR5), .S(_02421__PTR11), .Z(_02548__PTR5) );
  MUX2_X1 U10714 ( .A(_02487__PTR38), .B(_03274__PTR6), .S(_02421__PTR11), .Z(_02548__PTR6) );
  MUX2_X1 U10715 ( .A(_02487__PTR39), .B(_03274__PTR7), .S(_02421__PTR11), .Z(_02548__PTR7) );
  MUX2_X1 U10716 ( .A(_02485__PTR32), .B(_03273__PTR0), .S(_02421__PTR12), .Z(_02547__PTR0) );
  MUX2_X1 U10717 ( .A(_02485__PTR33), .B(_03274__PTR1), .S(_02421__PTR12), .Z(_02547__PTR1) );
  MUX2_X1 U10718 ( .A(_02485__PTR34), .B(_03274__PTR2), .S(_02421__PTR12), .Z(_02547__PTR2) );
  MUX2_X1 U10719 ( .A(_02485__PTR35), .B(_03274__PTR3), .S(_02421__PTR12), .Z(_02547__PTR3) );
  MUX2_X1 U10720 ( .A(_02485__PTR36), .B(_03274__PTR4), .S(_02421__PTR12), .Z(_02547__PTR4) );
  MUX2_X1 U10721 ( .A(_02485__PTR37), .B(_03274__PTR5), .S(_02421__PTR12), .Z(_02547__PTR5) );
  MUX2_X1 U10722 ( .A(_02485__PTR38), .B(_03274__PTR6), .S(_02421__PTR12), .Z(_02547__PTR6) );
  MUX2_X1 U10723 ( .A(_02485__PTR39), .B(_03274__PTR7), .S(_02421__PTR12), .Z(_02547__PTR7) );
  MUX2_X1 U10724 ( .A(_02483__PTR32), .B(_03273__PTR0), .S(_02421__PTR13), .Z(_02546__PTR0) );
  MUX2_X1 U10725 ( .A(_02483__PTR33), .B(_03274__PTR1), .S(_02421__PTR13), .Z(_02546__PTR1) );
  MUX2_X1 U10726 ( .A(_02483__PTR34), .B(_03274__PTR2), .S(_02421__PTR13), .Z(_02546__PTR2) );
  MUX2_X1 U10727 ( .A(_02483__PTR35), .B(_03274__PTR3), .S(_02421__PTR13), .Z(_02546__PTR3) );
  MUX2_X1 U10728 ( .A(_02483__PTR36), .B(_03274__PTR4), .S(_02421__PTR13), .Z(_02546__PTR4) );
  MUX2_X1 U10729 ( .A(_02483__PTR37), .B(_03274__PTR5), .S(_02421__PTR13), .Z(_02546__PTR5) );
  MUX2_X1 U10730 ( .A(_02483__PTR38), .B(_03274__PTR6), .S(_02421__PTR13), .Z(_02546__PTR6) );
  MUX2_X1 U10731 ( .A(_02483__PTR39), .B(_03274__PTR7), .S(_02421__PTR13), .Z(_02546__PTR7) );
  MUX2_X1 U10732 ( .A(_02481__PTR32), .B(_03273__PTR0), .S(_02421__PTR14), .Z(_02545__PTR0) );
  MUX2_X1 U10733 ( .A(_02481__PTR33), .B(_03274__PTR1), .S(_02421__PTR14), .Z(_02545__PTR1) );
  MUX2_X1 U10734 ( .A(_02481__PTR34), .B(_03274__PTR2), .S(_02421__PTR14), .Z(_02545__PTR2) );
  MUX2_X1 U10735 ( .A(_02481__PTR35), .B(_03274__PTR3), .S(_02421__PTR14), .Z(_02545__PTR3) );
  MUX2_X1 U10736 ( .A(_02481__PTR36), .B(_03274__PTR4), .S(_02421__PTR14), .Z(_02545__PTR4) );
  MUX2_X1 U10737 ( .A(_02481__PTR37), .B(_03274__PTR5), .S(_02421__PTR14), .Z(_02545__PTR5) );
  MUX2_X1 U10738 ( .A(_02481__PTR38), .B(_03274__PTR6), .S(_02421__PTR14), .Z(_02545__PTR6) );
  MUX2_X1 U10739 ( .A(_02481__PTR39), .B(_03274__PTR7), .S(_02421__PTR14), .Z(_02545__PTR7) );
  MUX2_X1 U10740 ( .A(_02479__PTR32), .B(_03273__PTR0), .S(_02421__PTR15), .Z(_02544__PTR0) );
  MUX2_X1 U10741 ( .A(_02479__PTR33), .B(_03274__PTR1), .S(_02421__PTR15), .Z(_02544__PTR1) );
  MUX2_X1 U10742 ( .A(_02479__PTR34), .B(_03274__PTR2), .S(_02421__PTR15), .Z(_02544__PTR2) );
  MUX2_X1 U10743 ( .A(_02479__PTR35), .B(_03274__PTR3), .S(_02421__PTR15), .Z(_02544__PTR3) );
  MUX2_X1 U10744 ( .A(_02479__PTR36), .B(_03274__PTR4), .S(_02421__PTR15), .Z(_02544__PTR4) );
  MUX2_X1 U10745 ( .A(_02479__PTR37), .B(_03274__PTR5), .S(_02421__PTR15), .Z(_02544__PTR5) );
  MUX2_X1 U10746 ( .A(_02479__PTR38), .B(_03274__PTR6), .S(_02421__PTR15), .Z(_02544__PTR6) );
  MUX2_X1 U10747 ( .A(_02479__PTR39), .B(_03274__PTR7), .S(_02421__PTR15), .Z(_02544__PTR7) );
  MUX2_X1 U10748 ( .A(_02543__PTR0), .B(buf2_PTR0), .S(_02419__PTR0), .Z(_02509__PTR32) );
  MUX2_X1 U10749 ( .A(_02543__PTR1), .B(buf2_PTR1), .S(_02419__PTR0), .Z(_02509__PTR33) );
  MUX2_X1 U10750 ( .A(_02543__PTR2), .B(buf2_PTR2), .S(_02419__PTR0), .Z(_02509__PTR34) );
  MUX2_X1 U10751 ( .A(_02543__PTR3), .B(buf2_PTR3), .S(_02419__PTR0), .Z(_02509__PTR35) );
  MUX2_X1 U10752 ( .A(_02543__PTR4), .B(buf2_PTR4), .S(_02419__PTR0), .Z(_02509__PTR36) );
  MUX2_X1 U10753 ( .A(_02543__PTR5), .B(buf2_PTR5), .S(_02419__PTR0), .Z(_02509__PTR37) );
  MUX2_X1 U10754 ( .A(_02543__PTR6), .B(buf2_PTR6), .S(_02419__PTR0), .Z(_02509__PTR38) );
  MUX2_X1 U10755 ( .A(_02543__PTR7), .B(buf2_PTR7), .S(_02419__PTR0), .Z(_02509__PTR39) );
  MUX2_X1 U10756 ( .A(_02542__PTR0), .B(buf2_PTR0), .S(_02419__PTR1), .Z(_02507__PTR32) );
  MUX2_X1 U10757 ( .A(_02542__PTR1), .B(buf2_PTR1), .S(_02419__PTR1), .Z(_02507__PTR33) );
  MUX2_X1 U10758 ( .A(_02542__PTR2), .B(buf2_PTR2), .S(_02419__PTR1), .Z(_02507__PTR34) );
  MUX2_X1 U10759 ( .A(_02542__PTR3), .B(buf2_PTR3), .S(_02419__PTR1), .Z(_02507__PTR35) );
  MUX2_X1 U10760 ( .A(_02542__PTR4), .B(buf2_PTR4), .S(_02419__PTR1), .Z(_02507__PTR36) );
  MUX2_X1 U10761 ( .A(_02542__PTR5), .B(buf2_PTR5), .S(_02419__PTR1), .Z(_02507__PTR37) );
  MUX2_X1 U10762 ( .A(_02542__PTR6), .B(buf2_PTR6), .S(_02419__PTR1), .Z(_02507__PTR38) );
  MUX2_X1 U10763 ( .A(_02542__PTR7), .B(buf2_PTR7), .S(_02419__PTR1), .Z(_02507__PTR39) );
  MUX2_X1 U10764 ( .A(_02541__PTR0), .B(buf2_PTR0), .S(_02419__PTR2), .Z(_02505__PTR32) );
  MUX2_X1 U10765 ( .A(_02541__PTR1), .B(buf2_PTR1), .S(_02419__PTR2), .Z(_02505__PTR33) );
  MUX2_X1 U10766 ( .A(_02541__PTR2), .B(buf2_PTR2), .S(_02419__PTR2), .Z(_02505__PTR34) );
  MUX2_X1 U10767 ( .A(_02541__PTR3), .B(buf2_PTR3), .S(_02419__PTR2), .Z(_02505__PTR35) );
  MUX2_X1 U10768 ( .A(_02541__PTR4), .B(buf2_PTR4), .S(_02419__PTR2), .Z(_02505__PTR36) );
  MUX2_X1 U10769 ( .A(_02541__PTR5), .B(buf2_PTR5), .S(_02419__PTR2), .Z(_02505__PTR37) );
  MUX2_X1 U10770 ( .A(_02541__PTR6), .B(buf2_PTR6), .S(_02419__PTR2), .Z(_02505__PTR38) );
  MUX2_X1 U10771 ( .A(_02541__PTR7), .B(buf2_PTR7), .S(_02419__PTR2), .Z(_02505__PTR39) );
  MUX2_X1 U10772 ( .A(_02540__PTR0), .B(buf2_PTR0), .S(_02419__PTR3), .Z(_02503__PTR32) );
  MUX2_X1 U10773 ( .A(_02540__PTR1), .B(buf2_PTR1), .S(_02419__PTR3), .Z(_02503__PTR33) );
  MUX2_X1 U10774 ( .A(_02540__PTR2), .B(buf2_PTR2), .S(_02419__PTR3), .Z(_02503__PTR34) );
  MUX2_X1 U10775 ( .A(_02540__PTR3), .B(buf2_PTR3), .S(_02419__PTR3), .Z(_02503__PTR35) );
  MUX2_X1 U10776 ( .A(_02540__PTR4), .B(buf2_PTR4), .S(_02419__PTR3), .Z(_02503__PTR36) );
  MUX2_X1 U10777 ( .A(_02540__PTR5), .B(buf2_PTR5), .S(_02419__PTR3), .Z(_02503__PTR37) );
  MUX2_X1 U10778 ( .A(_02540__PTR6), .B(buf2_PTR6), .S(_02419__PTR3), .Z(_02503__PTR38) );
  MUX2_X1 U10779 ( .A(_02540__PTR7), .B(buf2_PTR7), .S(_02419__PTR3), .Z(_02503__PTR39) );
  MUX2_X1 U10780 ( .A(_02539__PTR0), .B(buf2_PTR0), .S(_02419__PTR4), .Z(_02501__PTR32) );
  MUX2_X1 U10781 ( .A(_02539__PTR1), .B(buf2_PTR1), .S(_02419__PTR4), .Z(_02501__PTR33) );
  MUX2_X1 U10782 ( .A(_02539__PTR2), .B(buf2_PTR2), .S(_02419__PTR4), .Z(_02501__PTR34) );
  MUX2_X1 U10783 ( .A(_02539__PTR3), .B(buf2_PTR3), .S(_02419__PTR4), .Z(_02501__PTR35) );
  MUX2_X1 U10784 ( .A(_02539__PTR4), .B(buf2_PTR4), .S(_02419__PTR4), .Z(_02501__PTR36) );
  MUX2_X1 U10785 ( .A(_02539__PTR5), .B(buf2_PTR5), .S(_02419__PTR4), .Z(_02501__PTR37) );
  MUX2_X1 U10786 ( .A(_02539__PTR6), .B(buf2_PTR6), .S(_02419__PTR4), .Z(_02501__PTR38) );
  MUX2_X1 U10787 ( .A(_02539__PTR7), .B(buf2_PTR7), .S(_02419__PTR4), .Z(_02501__PTR39) );
  MUX2_X1 U10788 ( .A(_02538__PTR0), .B(buf2_PTR0), .S(_02419__PTR5), .Z(_02499__PTR32) );
  MUX2_X1 U10789 ( .A(_02538__PTR1), .B(buf2_PTR1), .S(_02419__PTR5), .Z(_02499__PTR33) );
  MUX2_X1 U10790 ( .A(_02538__PTR2), .B(buf2_PTR2), .S(_02419__PTR5), .Z(_02499__PTR34) );
  MUX2_X1 U10791 ( .A(_02538__PTR3), .B(buf2_PTR3), .S(_02419__PTR5), .Z(_02499__PTR35) );
  MUX2_X1 U10792 ( .A(_02538__PTR4), .B(buf2_PTR4), .S(_02419__PTR5), .Z(_02499__PTR36) );
  MUX2_X1 U10793 ( .A(_02538__PTR5), .B(buf2_PTR5), .S(_02419__PTR5), .Z(_02499__PTR37) );
  MUX2_X1 U10794 ( .A(_02538__PTR6), .B(buf2_PTR6), .S(_02419__PTR5), .Z(_02499__PTR38) );
  MUX2_X1 U10795 ( .A(_02538__PTR7), .B(buf2_PTR7), .S(_02419__PTR5), .Z(_02499__PTR39) );
  MUX2_X1 U10796 ( .A(_02537__PTR0), .B(buf2_PTR0), .S(_02419__PTR6), .Z(_02497__PTR32) );
  MUX2_X1 U10797 ( .A(_02537__PTR1), .B(buf2_PTR1), .S(_02419__PTR6), .Z(_02497__PTR33) );
  MUX2_X1 U10798 ( .A(_02537__PTR2), .B(buf2_PTR2), .S(_02419__PTR6), .Z(_02497__PTR34) );
  MUX2_X1 U10799 ( .A(_02537__PTR3), .B(buf2_PTR3), .S(_02419__PTR6), .Z(_02497__PTR35) );
  MUX2_X1 U10800 ( .A(_02537__PTR4), .B(buf2_PTR4), .S(_02419__PTR6), .Z(_02497__PTR36) );
  MUX2_X1 U10801 ( .A(_02537__PTR5), .B(buf2_PTR5), .S(_02419__PTR6), .Z(_02497__PTR37) );
  MUX2_X1 U10802 ( .A(_02537__PTR6), .B(buf2_PTR6), .S(_02419__PTR6), .Z(_02497__PTR38) );
  MUX2_X1 U10803 ( .A(_02537__PTR7), .B(buf2_PTR7), .S(_02419__PTR6), .Z(_02497__PTR39) );
  MUX2_X1 U10804 ( .A(_02536__PTR0), .B(buf2_PTR0), .S(_02419__PTR7), .Z(_02495__PTR32) );
  MUX2_X1 U10805 ( .A(_02536__PTR1), .B(buf2_PTR1), .S(_02419__PTR7), .Z(_02495__PTR33) );
  MUX2_X1 U10806 ( .A(_02536__PTR2), .B(buf2_PTR2), .S(_02419__PTR7), .Z(_02495__PTR34) );
  MUX2_X1 U10807 ( .A(_02536__PTR3), .B(buf2_PTR3), .S(_02419__PTR7), .Z(_02495__PTR35) );
  MUX2_X1 U10808 ( .A(_02536__PTR4), .B(buf2_PTR4), .S(_02419__PTR7), .Z(_02495__PTR36) );
  MUX2_X1 U10809 ( .A(_02536__PTR5), .B(buf2_PTR5), .S(_02419__PTR7), .Z(_02495__PTR37) );
  MUX2_X1 U10810 ( .A(_02536__PTR6), .B(buf2_PTR6), .S(_02419__PTR7), .Z(_02495__PTR38) );
  MUX2_X1 U10811 ( .A(_02536__PTR7), .B(buf2_PTR7), .S(_02419__PTR7), .Z(_02495__PTR39) );
  MUX2_X1 U10812 ( .A(_02535__PTR0), .B(buf2_PTR0), .S(_02419__PTR8), .Z(_02493__PTR32) );
  MUX2_X1 U10813 ( .A(_02535__PTR1), .B(buf2_PTR1), .S(_02419__PTR8), .Z(_02493__PTR33) );
  MUX2_X1 U10814 ( .A(_02535__PTR2), .B(buf2_PTR2), .S(_02419__PTR8), .Z(_02493__PTR34) );
  MUX2_X1 U10815 ( .A(_02535__PTR3), .B(buf2_PTR3), .S(_02419__PTR8), .Z(_02493__PTR35) );
  MUX2_X1 U10816 ( .A(_02535__PTR4), .B(buf2_PTR4), .S(_02419__PTR8), .Z(_02493__PTR36) );
  MUX2_X1 U10817 ( .A(_02535__PTR5), .B(buf2_PTR5), .S(_02419__PTR8), .Z(_02493__PTR37) );
  MUX2_X1 U10818 ( .A(_02535__PTR6), .B(buf2_PTR6), .S(_02419__PTR8), .Z(_02493__PTR38) );
  MUX2_X1 U10819 ( .A(_02535__PTR7), .B(buf2_PTR7), .S(_02419__PTR8), .Z(_02493__PTR39) );
  MUX2_X1 U10820 ( .A(_02534__PTR0), .B(buf2_PTR0), .S(_02419__PTR9), .Z(_02491__PTR32) );
  MUX2_X1 U10821 ( .A(_02534__PTR1), .B(buf2_PTR1), .S(_02419__PTR9), .Z(_02491__PTR33) );
  MUX2_X1 U10822 ( .A(_02534__PTR2), .B(buf2_PTR2), .S(_02419__PTR9), .Z(_02491__PTR34) );
  MUX2_X1 U10823 ( .A(_02534__PTR3), .B(buf2_PTR3), .S(_02419__PTR9), .Z(_02491__PTR35) );
  MUX2_X1 U10824 ( .A(_02534__PTR4), .B(buf2_PTR4), .S(_02419__PTR9), .Z(_02491__PTR36) );
  MUX2_X1 U10825 ( .A(_02534__PTR5), .B(buf2_PTR5), .S(_02419__PTR9), .Z(_02491__PTR37) );
  MUX2_X1 U10826 ( .A(_02534__PTR6), .B(buf2_PTR6), .S(_02419__PTR9), .Z(_02491__PTR38) );
  MUX2_X1 U10827 ( .A(_02534__PTR7), .B(buf2_PTR7), .S(_02419__PTR9), .Z(_02491__PTR39) );
  MUX2_X1 U10828 ( .A(_02533__PTR0), .B(buf2_PTR0), .S(_02419__PTR10), .Z(_02489__PTR32) );
  MUX2_X1 U10829 ( .A(_02533__PTR1), .B(buf2_PTR1), .S(_02419__PTR10), .Z(_02489__PTR33) );
  MUX2_X1 U10830 ( .A(_02533__PTR2), .B(buf2_PTR2), .S(_02419__PTR10), .Z(_02489__PTR34) );
  MUX2_X1 U10831 ( .A(_02533__PTR3), .B(buf2_PTR3), .S(_02419__PTR10), .Z(_02489__PTR35) );
  MUX2_X1 U10832 ( .A(_02533__PTR4), .B(buf2_PTR4), .S(_02419__PTR10), .Z(_02489__PTR36) );
  MUX2_X1 U10833 ( .A(_02533__PTR5), .B(buf2_PTR5), .S(_02419__PTR10), .Z(_02489__PTR37) );
  MUX2_X1 U10834 ( .A(_02533__PTR6), .B(buf2_PTR6), .S(_02419__PTR10), .Z(_02489__PTR38) );
  MUX2_X1 U10835 ( .A(_02533__PTR7), .B(buf2_PTR7), .S(_02419__PTR10), .Z(_02489__PTR39) );
  MUX2_X1 U10836 ( .A(_02532__PTR0), .B(buf2_PTR0), .S(_02419__PTR11), .Z(_02487__PTR32) );
  MUX2_X1 U10837 ( .A(_02532__PTR1), .B(buf2_PTR1), .S(_02419__PTR11), .Z(_02487__PTR33) );
  MUX2_X1 U10838 ( .A(_02532__PTR2), .B(buf2_PTR2), .S(_02419__PTR11), .Z(_02487__PTR34) );
  MUX2_X1 U10839 ( .A(_02532__PTR3), .B(buf2_PTR3), .S(_02419__PTR11), .Z(_02487__PTR35) );
  MUX2_X1 U10840 ( .A(_02532__PTR4), .B(buf2_PTR4), .S(_02419__PTR11), .Z(_02487__PTR36) );
  MUX2_X1 U10841 ( .A(_02532__PTR5), .B(buf2_PTR5), .S(_02419__PTR11), .Z(_02487__PTR37) );
  MUX2_X1 U10842 ( .A(_02532__PTR6), .B(buf2_PTR6), .S(_02419__PTR11), .Z(_02487__PTR38) );
  MUX2_X1 U10843 ( .A(_02532__PTR7), .B(buf2_PTR7), .S(_02419__PTR11), .Z(_02487__PTR39) );
  MUX2_X1 U10844 ( .A(_02531__PTR0), .B(buf2_PTR0), .S(_02419__PTR12), .Z(_02485__PTR32) );
  MUX2_X1 U10845 ( .A(_02531__PTR1), .B(buf2_PTR1), .S(_02419__PTR12), .Z(_02485__PTR33) );
  MUX2_X1 U10846 ( .A(_02531__PTR2), .B(buf2_PTR2), .S(_02419__PTR12), .Z(_02485__PTR34) );
  MUX2_X1 U10847 ( .A(_02531__PTR3), .B(buf2_PTR3), .S(_02419__PTR12), .Z(_02485__PTR35) );
  MUX2_X1 U10848 ( .A(_02531__PTR4), .B(buf2_PTR4), .S(_02419__PTR12), .Z(_02485__PTR36) );
  MUX2_X1 U10849 ( .A(_02531__PTR5), .B(buf2_PTR5), .S(_02419__PTR12), .Z(_02485__PTR37) );
  MUX2_X1 U10850 ( .A(_02531__PTR6), .B(buf2_PTR6), .S(_02419__PTR12), .Z(_02485__PTR38) );
  MUX2_X1 U10851 ( .A(_02531__PTR7), .B(buf2_PTR7), .S(_02419__PTR12), .Z(_02485__PTR39) );
  MUX2_X1 U10852 ( .A(_02530__PTR0), .B(buf2_PTR0), .S(_02419__PTR13), .Z(_02483__PTR32) );
  MUX2_X1 U10853 ( .A(_02530__PTR1), .B(buf2_PTR1), .S(_02419__PTR13), .Z(_02483__PTR33) );
  MUX2_X1 U10854 ( .A(_02530__PTR2), .B(buf2_PTR2), .S(_02419__PTR13), .Z(_02483__PTR34) );
  MUX2_X1 U10855 ( .A(_02530__PTR3), .B(buf2_PTR3), .S(_02419__PTR13), .Z(_02483__PTR35) );
  MUX2_X1 U10856 ( .A(_02530__PTR4), .B(buf2_PTR4), .S(_02419__PTR13), .Z(_02483__PTR36) );
  MUX2_X1 U10857 ( .A(_02530__PTR5), .B(buf2_PTR5), .S(_02419__PTR13), .Z(_02483__PTR37) );
  MUX2_X1 U10858 ( .A(_02530__PTR6), .B(buf2_PTR6), .S(_02419__PTR13), .Z(_02483__PTR38) );
  MUX2_X1 U10859 ( .A(_02530__PTR7), .B(buf2_PTR7), .S(_02419__PTR13), .Z(_02483__PTR39) );
  MUX2_X1 U10860 ( .A(_02529__PTR0), .B(buf2_PTR0), .S(_02419__PTR14), .Z(_02481__PTR32) );
  MUX2_X1 U10861 ( .A(_02529__PTR1), .B(buf2_PTR1), .S(_02419__PTR14), .Z(_02481__PTR33) );
  MUX2_X1 U10862 ( .A(_02529__PTR2), .B(buf2_PTR2), .S(_02419__PTR14), .Z(_02481__PTR34) );
  MUX2_X1 U10863 ( .A(_02529__PTR3), .B(buf2_PTR3), .S(_02419__PTR14), .Z(_02481__PTR35) );
  MUX2_X1 U10864 ( .A(_02529__PTR4), .B(buf2_PTR4), .S(_02419__PTR14), .Z(_02481__PTR36) );
  MUX2_X1 U10865 ( .A(_02529__PTR5), .B(buf2_PTR5), .S(_02419__PTR14), .Z(_02481__PTR37) );
  MUX2_X1 U10866 ( .A(_02529__PTR6), .B(buf2_PTR6), .S(_02419__PTR14), .Z(_02481__PTR38) );
  MUX2_X1 U10867 ( .A(_02529__PTR7), .B(buf2_PTR7), .S(_02419__PTR14), .Z(_02481__PTR39) );
  MUX2_X1 U10868 ( .A(_02528__PTR0), .B(buf2_PTR0), .S(_02419__PTR15), .Z(_02479__PTR32) );
  MUX2_X1 U10869 ( .A(_02528__PTR1), .B(buf2_PTR1), .S(_02419__PTR15), .Z(_02479__PTR33) );
  MUX2_X1 U10870 ( .A(_02528__PTR2), .B(buf2_PTR2), .S(_02419__PTR15), .Z(_02479__PTR34) );
  MUX2_X1 U10871 ( .A(_02528__PTR3), .B(buf2_PTR3), .S(_02419__PTR15), .Z(_02479__PTR35) );
  MUX2_X1 U10872 ( .A(_02528__PTR4), .B(buf2_PTR4), .S(_02419__PTR15), .Z(_02479__PTR36) );
  MUX2_X1 U10873 ( .A(_02528__PTR5), .B(buf2_PTR5), .S(_02419__PTR15), .Z(_02479__PTR37) );
  MUX2_X1 U10874 ( .A(_02528__PTR6), .B(buf2_PTR6), .S(_02419__PTR15), .Z(_02479__PTR38) );
  MUX2_X1 U10875 ( .A(_02528__PTR7), .B(buf2_PTR7), .S(_02419__PTR15), .Z(_02479__PTR39) );
  MUX2_X1 U10876 ( .A(P3_P1_InstQueue_PTR0_PTR0), .B(buf2_PTR0), .S(_02417__PTR0), .Z(_02543__PTR0) );
  MUX2_X1 U10877 ( .A(P3_P1_InstQueue_PTR0_PTR1), .B(buf2_PTR1), .S(_02417__PTR0), .Z(_02543__PTR1) );
  MUX2_X1 U10878 ( .A(P3_P1_InstQueue_PTR0_PTR2), .B(buf2_PTR2), .S(_02417__PTR0), .Z(_02543__PTR2) );
  MUX2_X1 U10879 ( .A(P3_P1_InstQueue_PTR0_PTR3), .B(buf2_PTR3), .S(_02417__PTR0), .Z(_02543__PTR3) );
  MUX2_X1 U10880 ( .A(P3_P1_InstQueue_PTR0_PTR4), .B(buf2_PTR4), .S(_02417__PTR0), .Z(_02543__PTR4) );
  MUX2_X1 U10881 ( .A(P3_P1_InstQueue_PTR0_PTR5), .B(buf2_PTR5), .S(_02417__PTR0), .Z(_02543__PTR5) );
  MUX2_X1 U10882 ( .A(P3_P1_InstQueue_PTR0_PTR6), .B(buf2_PTR6), .S(_02417__PTR0), .Z(_02543__PTR6) );
  MUX2_X1 U10883 ( .A(P3_P1_InstQueue_PTR0_PTR7), .B(buf2_PTR7), .S(_02417__PTR0), .Z(_02543__PTR7) );
  MUX2_X1 U10884 ( .A(P3_P1_InstQueue_PTR1_PTR0), .B(buf2_PTR0), .S(_02417__PTR1), .Z(_02542__PTR0) );
  MUX2_X1 U10885 ( .A(P3_P1_InstQueue_PTR1_PTR1), .B(buf2_PTR1), .S(_02417__PTR1), .Z(_02542__PTR1) );
  MUX2_X1 U10886 ( .A(P3_P1_InstQueue_PTR1_PTR2), .B(buf2_PTR2), .S(_02417__PTR1), .Z(_02542__PTR2) );
  MUX2_X1 U10887 ( .A(P3_P1_InstQueue_PTR1_PTR3), .B(buf2_PTR3), .S(_02417__PTR1), .Z(_02542__PTR3) );
  MUX2_X1 U10888 ( .A(P3_P1_InstQueue_PTR1_PTR4), .B(buf2_PTR4), .S(_02417__PTR1), .Z(_02542__PTR4) );
  MUX2_X1 U10889 ( .A(P3_P1_InstQueue_PTR1_PTR5), .B(buf2_PTR5), .S(_02417__PTR1), .Z(_02542__PTR5) );
  MUX2_X1 U10890 ( .A(P3_P1_InstQueue_PTR1_PTR6), .B(buf2_PTR6), .S(_02417__PTR1), .Z(_02542__PTR6) );
  MUX2_X1 U10891 ( .A(P3_P1_InstQueue_PTR1_PTR7), .B(buf2_PTR7), .S(_02417__PTR1), .Z(_02542__PTR7) );
  MUX2_X1 U10892 ( .A(P3_P1_InstQueue_PTR2_PTR0), .B(buf2_PTR0), .S(_02417__PTR2), .Z(_02541__PTR0) );
  MUX2_X1 U10893 ( .A(P3_P1_InstQueue_PTR2_PTR1), .B(buf2_PTR1), .S(_02417__PTR2), .Z(_02541__PTR1) );
  MUX2_X1 U10894 ( .A(P3_P1_InstQueue_PTR2_PTR2), .B(buf2_PTR2), .S(_02417__PTR2), .Z(_02541__PTR2) );
  MUX2_X1 U10895 ( .A(P3_P1_InstQueue_PTR2_PTR3), .B(buf2_PTR3), .S(_02417__PTR2), .Z(_02541__PTR3) );
  MUX2_X1 U10896 ( .A(P3_P1_InstQueue_PTR2_PTR4), .B(buf2_PTR4), .S(_02417__PTR2), .Z(_02541__PTR4) );
  MUX2_X1 U10897 ( .A(P3_P1_InstQueue_PTR2_PTR5), .B(buf2_PTR5), .S(_02417__PTR2), .Z(_02541__PTR5) );
  MUX2_X1 U10898 ( .A(P3_P1_InstQueue_PTR2_PTR6), .B(buf2_PTR6), .S(_02417__PTR2), .Z(_02541__PTR6) );
  MUX2_X1 U10899 ( .A(P3_P1_InstQueue_PTR2_PTR7), .B(buf2_PTR7), .S(_02417__PTR2), .Z(_02541__PTR7) );
  MUX2_X1 U10900 ( .A(P3_P1_InstQueue_PTR3_PTR0), .B(buf2_PTR0), .S(_02417__PTR3), .Z(_02540__PTR0) );
  MUX2_X1 U10901 ( .A(P3_P1_InstQueue_PTR3_PTR1), .B(buf2_PTR1), .S(_02417__PTR3), .Z(_02540__PTR1) );
  MUX2_X1 U10902 ( .A(P3_P1_InstQueue_PTR3_PTR2), .B(buf2_PTR2), .S(_02417__PTR3), .Z(_02540__PTR2) );
  MUX2_X1 U10903 ( .A(P3_P1_InstQueue_PTR3_PTR3), .B(buf2_PTR3), .S(_02417__PTR3), .Z(_02540__PTR3) );
  MUX2_X1 U10904 ( .A(P3_P1_InstQueue_PTR3_PTR4), .B(buf2_PTR4), .S(_02417__PTR3), .Z(_02540__PTR4) );
  MUX2_X1 U10905 ( .A(P3_P1_InstQueue_PTR3_PTR5), .B(buf2_PTR5), .S(_02417__PTR3), .Z(_02540__PTR5) );
  MUX2_X1 U10906 ( .A(P3_P1_InstQueue_PTR3_PTR6), .B(buf2_PTR6), .S(_02417__PTR3), .Z(_02540__PTR6) );
  MUX2_X1 U10907 ( .A(P3_P1_InstQueue_PTR3_PTR7), .B(buf2_PTR7), .S(_02417__PTR3), .Z(_02540__PTR7) );
  MUX2_X1 U10908 ( .A(P3_P1_InstQueue_PTR4_PTR0), .B(buf2_PTR0), .S(_02417__PTR4), .Z(_02539__PTR0) );
  MUX2_X1 U10909 ( .A(P3_P1_InstQueue_PTR4_PTR1), .B(buf2_PTR1), .S(_02417__PTR4), .Z(_02539__PTR1) );
  MUX2_X1 U10910 ( .A(P3_P1_InstQueue_PTR4_PTR2), .B(buf2_PTR2), .S(_02417__PTR4), .Z(_02539__PTR2) );
  MUX2_X1 U10911 ( .A(P3_P1_InstQueue_PTR4_PTR3), .B(buf2_PTR3), .S(_02417__PTR4), .Z(_02539__PTR3) );
  MUX2_X1 U10912 ( .A(P3_P1_InstQueue_PTR4_PTR4), .B(buf2_PTR4), .S(_02417__PTR4), .Z(_02539__PTR4) );
  MUX2_X1 U10913 ( .A(P3_P1_InstQueue_PTR4_PTR5), .B(buf2_PTR5), .S(_02417__PTR4), .Z(_02539__PTR5) );
  MUX2_X1 U10914 ( .A(P3_P1_InstQueue_PTR4_PTR6), .B(buf2_PTR6), .S(_02417__PTR4), .Z(_02539__PTR6) );
  MUX2_X1 U10915 ( .A(P3_P1_InstQueue_PTR4_PTR7), .B(buf2_PTR7), .S(_02417__PTR4), .Z(_02539__PTR7) );
  MUX2_X1 U10916 ( .A(P3_P1_InstQueue_PTR5_PTR0), .B(buf2_PTR0), .S(_02417__PTR5), .Z(_02538__PTR0) );
  MUX2_X1 U10917 ( .A(P3_P1_InstQueue_PTR5_PTR1), .B(buf2_PTR1), .S(_02417__PTR5), .Z(_02538__PTR1) );
  MUX2_X1 U10918 ( .A(P3_P1_InstQueue_PTR5_PTR2), .B(buf2_PTR2), .S(_02417__PTR5), .Z(_02538__PTR2) );
  MUX2_X1 U10919 ( .A(P3_P1_InstQueue_PTR5_PTR3), .B(buf2_PTR3), .S(_02417__PTR5), .Z(_02538__PTR3) );
  MUX2_X1 U10920 ( .A(P3_P1_InstQueue_PTR5_PTR4), .B(buf2_PTR4), .S(_02417__PTR5), .Z(_02538__PTR4) );
  MUX2_X1 U10921 ( .A(P3_P1_InstQueue_PTR5_PTR5), .B(buf2_PTR5), .S(_02417__PTR5), .Z(_02538__PTR5) );
  MUX2_X1 U10922 ( .A(P3_P1_InstQueue_PTR5_PTR6), .B(buf2_PTR6), .S(_02417__PTR5), .Z(_02538__PTR6) );
  MUX2_X1 U10923 ( .A(P3_P1_InstQueue_PTR5_PTR7), .B(buf2_PTR7), .S(_02417__PTR5), .Z(_02538__PTR7) );
  MUX2_X1 U10924 ( .A(P3_P1_InstQueue_PTR6_PTR0), .B(buf2_PTR0), .S(_02417__PTR6), .Z(_02537__PTR0) );
  MUX2_X1 U10925 ( .A(P3_P1_InstQueue_PTR6_PTR1), .B(buf2_PTR1), .S(_02417__PTR6), .Z(_02537__PTR1) );
  MUX2_X1 U10926 ( .A(P3_P1_InstQueue_PTR6_PTR2), .B(buf2_PTR2), .S(_02417__PTR6), .Z(_02537__PTR2) );
  MUX2_X1 U10927 ( .A(P3_P1_InstQueue_PTR6_PTR3), .B(buf2_PTR3), .S(_02417__PTR6), .Z(_02537__PTR3) );
  MUX2_X1 U10928 ( .A(P3_P1_InstQueue_PTR6_PTR4), .B(buf2_PTR4), .S(_02417__PTR6), .Z(_02537__PTR4) );
  MUX2_X1 U10929 ( .A(P3_P1_InstQueue_PTR6_PTR5), .B(buf2_PTR5), .S(_02417__PTR6), .Z(_02537__PTR5) );
  MUX2_X1 U10930 ( .A(P3_P1_InstQueue_PTR6_PTR6), .B(buf2_PTR6), .S(_02417__PTR6), .Z(_02537__PTR6) );
  MUX2_X1 U10931 ( .A(P3_P1_InstQueue_PTR6_PTR7), .B(buf2_PTR7), .S(_02417__PTR6), .Z(_02537__PTR7) );
  MUX2_X1 U10932 ( .A(P3_P1_InstQueue_PTR7_PTR0), .B(buf2_PTR0), .S(_02417__PTR7), .Z(_02536__PTR0) );
  MUX2_X1 U10933 ( .A(P3_P1_InstQueue_PTR7_PTR1), .B(buf2_PTR1), .S(_02417__PTR7), .Z(_02536__PTR1) );
  MUX2_X1 U10934 ( .A(P3_P1_InstQueue_PTR7_PTR2), .B(buf2_PTR2), .S(_02417__PTR7), .Z(_02536__PTR2) );
  MUX2_X1 U10935 ( .A(P3_P1_InstQueue_PTR7_PTR3), .B(buf2_PTR3), .S(_02417__PTR7), .Z(_02536__PTR3) );
  MUX2_X1 U10936 ( .A(P3_P1_InstQueue_PTR7_PTR4), .B(buf2_PTR4), .S(_02417__PTR7), .Z(_02536__PTR4) );
  MUX2_X1 U10937 ( .A(P3_P1_InstQueue_PTR7_PTR5), .B(buf2_PTR5), .S(_02417__PTR7), .Z(_02536__PTR5) );
  MUX2_X1 U10938 ( .A(P3_P1_InstQueue_PTR7_PTR6), .B(buf2_PTR6), .S(_02417__PTR7), .Z(_02536__PTR6) );
  MUX2_X1 U10939 ( .A(P3_P1_InstQueue_PTR7_PTR7), .B(buf2_PTR7), .S(_02417__PTR7), .Z(_02536__PTR7) );
  MUX2_X1 U10940 ( .A(P3_P1_InstQueue_PTR8_PTR0), .B(buf2_PTR0), .S(_02417__PTR8), .Z(_02535__PTR0) );
  MUX2_X1 U10941 ( .A(P3_P1_InstQueue_PTR8_PTR1), .B(buf2_PTR1), .S(_02417__PTR8), .Z(_02535__PTR1) );
  MUX2_X1 U10942 ( .A(P3_P1_InstQueue_PTR8_PTR2), .B(buf2_PTR2), .S(_02417__PTR8), .Z(_02535__PTR2) );
  MUX2_X1 U10943 ( .A(P3_P1_InstQueue_PTR8_PTR3), .B(buf2_PTR3), .S(_02417__PTR8), .Z(_02535__PTR3) );
  MUX2_X1 U10944 ( .A(P3_P1_InstQueue_PTR8_PTR4), .B(buf2_PTR4), .S(_02417__PTR8), .Z(_02535__PTR4) );
  MUX2_X1 U10945 ( .A(P3_P1_InstQueue_PTR8_PTR5), .B(buf2_PTR5), .S(_02417__PTR8), .Z(_02535__PTR5) );
  MUX2_X1 U10946 ( .A(P3_P1_InstQueue_PTR8_PTR6), .B(buf2_PTR6), .S(_02417__PTR8), .Z(_02535__PTR6) );
  MUX2_X1 U10947 ( .A(P3_P1_InstQueue_PTR8_PTR7), .B(buf2_PTR7), .S(_02417__PTR8), .Z(_02535__PTR7) );
  MUX2_X1 U10948 ( .A(P3_P1_InstQueue_PTR9_PTR0), .B(buf2_PTR0), .S(_02417__PTR9), .Z(_02534__PTR0) );
  MUX2_X1 U10949 ( .A(P3_P1_InstQueue_PTR9_PTR1), .B(buf2_PTR1), .S(_02417__PTR9), .Z(_02534__PTR1) );
  MUX2_X1 U10950 ( .A(P3_P1_InstQueue_PTR9_PTR2), .B(buf2_PTR2), .S(_02417__PTR9), .Z(_02534__PTR2) );
  MUX2_X1 U10951 ( .A(P3_P1_InstQueue_PTR9_PTR3), .B(buf2_PTR3), .S(_02417__PTR9), .Z(_02534__PTR3) );
  MUX2_X1 U10952 ( .A(P3_P1_InstQueue_PTR9_PTR4), .B(buf2_PTR4), .S(_02417__PTR9), .Z(_02534__PTR4) );
  MUX2_X1 U10953 ( .A(P3_P1_InstQueue_PTR9_PTR5), .B(buf2_PTR5), .S(_02417__PTR9), .Z(_02534__PTR5) );
  MUX2_X1 U10954 ( .A(P3_P1_InstQueue_PTR9_PTR6), .B(buf2_PTR6), .S(_02417__PTR9), .Z(_02534__PTR6) );
  MUX2_X1 U10955 ( .A(P3_P1_InstQueue_PTR9_PTR7), .B(buf2_PTR7), .S(_02417__PTR9), .Z(_02534__PTR7) );
  MUX2_X1 U10956 ( .A(P3_P1_InstQueue_PTR10_PTR0), .B(buf2_PTR0), .S(_02417__PTR10), .Z(_02533__PTR0) );
  MUX2_X1 U10957 ( .A(P3_P1_InstQueue_PTR10_PTR1), .B(buf2_PTR1), .S(_02417__PTR10), .Z(_02533__PTR1) );
  MUX2_X1 U10958 ( .A(P3_P1_InstQueue_PTR10_PTR2), .B(buf2_PTR2), .S(_02417__PTR10), .Z(_02533__PTR2) );
  MUX2_X1 U10959 ( .A(P3_P1_InstQueue_PTR10_PTR3), .B(buf2_PTR3), .S(_02417__PTR10), .Z(_02533__PTR3) );
  MUX2_X1 U10960 ( .A(P3_P1_InstQueue_PTR10_PTR4), .B(buf2_PTR4), .S(_02417__PTR10), .Z(_02533__PTR4) );
  MUX2_X1 U10961 ( .A(P3_P1_InstQueue_PTR10_PTR5), .B(buf2_PTR5), .S(_02417__PTR10), .Z(_02533__PTR5) );
  MUX2_X1 U10962 ( .A(P3_P1_InstQueue_PTR10_PTR6), .B(buf2_PTR6), .S(_02417__PTR10), .Z(_02533__PTR6) );
  MUX2_X1 U10963 ( .A(P3_P1_InstQueue_PTR10_PTR7), .B(buf2_PTR7), .S(_02417__PTR10), .Z(_02533__PTR7) );
  MUX2_X1 U10964 ( .A(P3_P1_InstQueue_PTR11_PTR0), .B(buf2_PTR0), .S(_02417__PTR11), .Z(_02532__PTR0) );
  MUX2_X1 U10965 ( .A(P3_P1_InstQueue_PTR11_PTR1), .B(buf2_PTR1), .S(_02417__PTR11), .Z(_02532__PTR1) );
  MUX2_X1 U10966 ( .A(P3_P1_InstQueue_PTR11_PTR2), .B(buf2_PTR2), .S(_02417__PTR11), .Z(_02532__PTR2) );
  MUX2_X1 U10967 ( .A(P3_P1_InstQueue_PTR11_PTR3), .B(buf2_PTR3), .S(_02417__PTR11), .Z(_02532__PTR3) );
  MUX2_X1 U10968 ( .A(P3_P1_InstQueue_PTR11_PTR4), .B(buf2_PTR4), .S(_02417__PTR11), .Z(_02532__PTR4) );
  MUX2_X1 U10969 ( .A(P3_P1_InstQueue_PTR11_PTR5), .B(buf2_PTR5), .S(_02417__PTR11), .Z(_02532__PTR5) );
  MUX2_X1 U10970 ( .A(P3_P1_InstQueue_PTR11_PTR6), .B(buf2_PTR6), .S(_02417__PTR11), .Z(_02532__PTR6) );
  MUX2_X1 U10971 ( .A(P3_P1_InstQueue_PTR11_PTR7), .B(buf2_PTR7), .S(_02417__PTR11), .Z(_02532__PTR7) );
  MUX2_X1 U10972 ( .A(P3_P1_InstQueue_PTR12_PTR0), .B(buf2_PTR0), .S(_02417__PTR12), .Z(_02531__PTR0) );
  MUX2_X1 U10973 ( .A(P3_P1_InstQueue_PTR12_PTR1), .B(buf2_PTR1), .S(_02417__PTR12), .Z(_02531__PTR1) );
  MUX2_X1 U10974 ( .A(P3_P1_InstQueue_PTR12_PTR2), .B(buf2_PTR2), .S(_02417__PTR12), .Z(_02531__PTR2) );
  MUX2_X1 U10975 ( .A(P3_P1_InstQueue_PTR12_PTR3), .B(buf2_PTR3), .S(_02417__PTR12), .Z(_02531__PTR3) );
  MUX2_X1 U10976 ( .A(P3_P1_InstQueue_PTR12_PTR4), .B(buf2_PTR4), .S(_02417__PTR12), .Z(_02531__PTR4) );
  MUX2_X1 U10977 ( .A(P3_P1_InstQueue_PTR12_PTR5), .B(buf2_PTR5), .S(_02417__PTR12), .Z(_02531__PTR5) );
  MUX2_X1 U10978 ( .A(P3_P1_InstQueue_PTR12_PTR6), .B(buf2_PTR6), .S(_02417__PTR12), .Z(_02531__PTR6) );
  MUX2_X1 U10979 ( .A(P3_P1_InstQueue_PTR12_PTR7), .B(buf2_PTR7), .S(_02417__PTR12), .Z(_02531__PTR7) );
  MUX2_X1 U10980 ( .A(P3_P1_InstQueue_PTR13_PTR0), .B(buf2_PTR0), .S(_02417__PTR13), .Z(_02530__PTR0) );
  MUX2_X1 U10981 ( .A(P3_P1_InstQueue_PTR13_PTR1), .B(buf2_PTR1), .S(_02417__PTR13), .Z(_02530__PTR1) );
  MUX2_X1 U10982 ( .A(P3_P1_InstQueue_PTR13_PTR2), .B(buf2_PTR2), .S(_02417__PTR13), .Z(_02530__PTR2) );
  MUX2_X1 U10983 ( .A(P3_P1_InstQueue_PTR13_PTR3), .B(buf2_PTR3), .S(_02417__PTR13), .Z(_02530__PTR3) );
  MUX2_X1 U10984 ( .A(P3_P1_InstQueue_PTR13_PTR4), .B(buf2_PTR4), .S(_02417__PTR13), .Z(_02530__PTR4) );
  MUX2_X1 U10985 ( .A(P3_P1_InstQueue_PTR13_PTR5), .B(buf2_PTR5), .S(_02417__PTR13), .Z(_02530__PTR5) );
  MUX2_X1 U10986 ( .A(P3_P1_InstQueue_PTR13_PTR6), .B(buf2_PTR6), .S(_02417__PTR13), .Z(_02530__PTR6) );
  MUX2_X1 U10987 ( .A(P3_P1_InstQueue_PTR13_PTR7), .B(buf2_PTR7), .S(_02417__PTR13), .Z(_02530__PTR7) );
  MUX2_X1 U10988 ( .A(P3_P1_InstQueue_PTR14_PTR0), .B(buf2_PTR0), .S(_02417__PTR14), .Z(_02529__PTR0) );
  MUX2_X1 U10989 ( .A(P3_P1_InstQueue_PTR14_PTR1), .B(buf2_PTR1), .S(_02417__PTR14), .Z(_02529__PTR1) );
  MUX2_X1 U10990 ( .A(P3_P1_InstQueue_PTR14_PTR2), .B(buf2_PTR2), .S(_02417__PTR14), .Z(_02529__PTR2) );
  MUX2_X1 U10991 ( .A(P3_P1_InstQueue_PTR14_PTR3), .B(buf2_PTR3), .S(_02417__PTR14), .Z(_02529__PTR3) );
  MUX2_X1 U10992 ( .A(P3_P1_InstQueue_PTR14_PTR4), .B(buf2_PTR4), .S(_02417__PTR14), .Z(_02529__PTR4) );
  MUX2_X1 U10993 ( .A(P3_P1_InstQueue_PTR14_PTR5), .B(buf2_PTR5), .S(_02417__PTR14), .Z(_02529__PTR5) );
  MUX2_X1 U10994 ( .A(P3_P1_InstQueue_PTR14_PTR6), .B(buf2_PTR6), .S(_02417__PTR14), .Z(_02529__PTR6) );
  MUX2_X1 U10995 ( .A(P3_P1_InstQueue_PTR14_PTR7), .B(buf2_PTR7), .S(_02417__PTR14), .Z(_02529__PTR7) );
  MUX2_X1 U10996 ( .A(P3_P1_InstQueue_PTR15_PTR0), .B(buf2_PTR0), .S(_02417__PTR15), .Z(_02528__PTR0) );
  MUX2_X1 U10997 ( .A(P3_P1_InstQueue_PTR15_PTR1), .B(buf2_PTR1), .S(_02417__PTR15), .Z(_02528__PTR1) );
  MUX2_X1 U10998 ( .A(P3_P1_InstQueue_PTR15_PTR2), .B(buf2_PTR2), .S(_02417__PTR15), .Z(_02528__PTR2) );
  MUX2_X1 U10999 ( .A(P3_P1_InstQueue_PTR15_PTR3), .B(buf2_PTR3), .S(_02417__PTR15), .Z(_02528__PTR3) );
  MUX2_X1 U11000 ( .A(P3_P1_InstQueue_PTR15_PTR4), .B(buf2_PTR4), .S(_02417__PTR15), .Z(_02528__PTR4) );
  MUX2_X1 U11001 ( .A(P3_P1_InstQueue_PTR15_PTR5), .B(buf2_PTR5), .S(_02417__PTR15), .Z(_02528__PTR5) );
  MUX2_X1 U11002 ( .A(P3_P1_InstQueue_PTR15_PTR6), .B(buf2_PTR6), .S(_02417__PTR15), .Z(_02528__PTR6) );
  MUX2_X1 U11003 ( .A(P3_P1_InstQueue_PTR15_PTR7), .B(buf2_PTR7), .S(_02417__PTR15), .Z(_02528__PTR7) );
  MUX2_X1 U11004 ( .A(_02527__PTR0), .B(1'b0), .S(_02522_), .Z(_02458__PTR28) );
  MUX2_X1 U11005 ( .A(_02527__PTR1), .B(1'b1), .S(_02522_), .Z(_02458__PTR29) );
  MUX2_X1 U11006 ( .A(_02527__PTR2), .B(1'b1), .S(_02522_), .Z(_02458__PTR30) );
  MUX2_X1 U11007 ( .A(_02526__PTR0), .B(1'b1), .S(_02523_), .Z(_02527__PTR0) );
  MUX2_X1 U11008 ( .A(_02526__PTR1), .B(1'b0), .S(_02523_), .Z(_02527__PTR1) );
  MUX2_X1 U11009 ( .A(_02526__PTR2), .B(1'b1), .S(_02523_), .Z(_02527__PTR2) );
  INV_X1 U11010 ( .A(_01765__PTR4), .ZN(_02526__PTR0) );
  MUX2_X1 U11011 ( .A(_02525__PTR2), .B(1'b1), .S(_01765__PTR4), .Z(_02526__PTR1) );
  MUX2_X1 U11012 ( .A(_02525__PTR2), .B(1'b0), .S(_01765__PTR4), .Z(_02526__PTR2) );
  INV_X1 U11013 ( .A(_02524_), .ZN(_02525__PTR2) );
  MUX2_X1 U11014 ( .A(P3_EAX_PTR16), .B(_02623__PTR16), .S(_02585_), .Z(_02674__PTR80) );
  MUX2_X1 U11015 ( .A(P3_EAX_PTR17), .B(_02623__PTR17), .S(_02585_), .Z(_02674__PTR81) );
  MUX2_X1 U11016 ( .A(P3_EAX_PTR18), .B(_02623__PTR18), .S(_02585_), .Z(_02674__PTR82) );
  MUX2_X1 U11017 ( .A(P3_EAX_PTR19), .B(_02623__PTR19), .S(_02585_), .Z(_02674__PTR83) );
  MUX2_X1 U11018 ( .A(P3_EAX_PTR20), .B(_02623__PTR20), .S(_02585_), .Z(_02674__PTR84) );
  MUX2_X1 U11019 ( .A(P3_EAX_PTR21), .B(_02623__PTR21), .S(_02585_), .Z(_02674__PTR85) );
  MUX2_X1 U11020 ( .A(P3_EAX_PTR22), .B(_02623__PTR22), .S(_02585_), .Z(_02674__PTR86) );
  MUX2_X1 U11021 ( .A(P3_EAX_PTR23), .B(_02623__PTR23), .S(_02585_), .Z(_02674__PTR87) );
  MUX2_X1 U11022 ( .A(P3_EAX_PTR24), .B(_02623__PTR24), .S(_02585_), .Z(_02674__PTR88) );
  MUX2_X1 U11023 ( .A(P3_EAX_PTR25), .B(_02623__PTR25), .S(_02585_), .Z(_02674__PTR89) );
  MUX2_X1 U11024 ( .A(P3_EAX_PTR26), .B(_02623__PTR26), .S(_02585_), .Z(_02674__PTR90) );
  MUX2_X1 U11025 ( .A(P3_EAX_PTR27), .B(_02623__PTR27), .S(_02585_), .Z(_02674__PTR91) );
  MUX2_X1 U11026 ( .A(P3_EAX_PTR28), .B(_02623__PTR28), .S(_02585_), .Z(_02674__PTR92) );
  MUX2_X1 U11027 ( .A(P3_EAX_PTR29), .B(_02623__PTR29), .S(_02585_), .Z(_02674__PTR93) );
  MUX2_X1 U11028 ( .A(P3_EAX_PTR30), .B(_02623__PTR30), .S(_02585_), .Z(_02674__PTR94) );
  MUX2_X1 U11029 ( .A(P3_EAX_PTR31), .B(_02623__PTR31), .S(_02585_), .Z(_02674__PTR95) );
  MUX2_X1 U11030 ( .A(P3_EAX_PTR0), .B(_02595__PTR0), .S(_02585_), .Z(_02674__PTR96) );
  MUX2_X1 U11031 ( .A(P3_EAX_PTR1), .B(_02595__PTR1), .S(_02585_), .Z(_02674__PTR97) );
  MUX2_X1 U11032 ( .A(P3_EAX_PTR2), .B(_02595__PTR2), .S(_02585_), .Z(_02674__PTR98) );
  MUX2_X1 U11033 ( .A(P3_EAX_PTR3), .B(_02595__PTR3), .S(_02585_), .Z(_02674__PTR99) );
  MUX2_X1 U11034 ( .A(P3_EAX_PTR4), .B(_02595__PTR4), .S(_02585_), .Z(_02674__PTR100) );
  MUX2_X1 U11035 ( .A(P3_EAX_PTR5), .B(_02595__PTR5), .S(_02585_), .Z(_02674__PTR101) );
  MUX2_X1 U11036 ( .A(P3_EAX_PTR6), .B(_02595__PTR6), .S(_02585_), .Z(_02674__PTR102) );
  MUX2_X1 U11037 ( .A(P3_EAX_PTR7), .B(_02595__PTR7), .S(_02585_), .Z(_02674__PTR103) );
  MUX2_X1 U11038 ( .A(P3_EAX_PTR8), .B(_02595__PTR8), .S(_02585_), .Z(_02674__PTR104) );
  MUX2_X1 U11039 ( .A(P3_EAX_PTR9), .B(_02595__PTR9), .S(_02585_), .Z(_02674__PTR105) );
  MUX2_X1 U11040 ( .A(P3_EAX_PTR10), .B(_02595__PTR10), .S(_02585_), .Z(_02674__PTR106) );
  MUX2_X1 U11041 ( .A(P3_EAX_PTR11), .B(_02595__PTR11), .S(_02585_), .Z(_02674__PTR107) );
  MUX2_X1 U11042 ( .A(P3_EAX_PTR12), .B(_02595__PTR12), .S(_02585_), .Z(_02674__PTR108) );
  MUX2_X1 U11043 ( .A(P3_EAX_PTR13), .B(_02595__PTR13), .S(_02585_), .Z(_02674__PTR109) );
  MUX2_X1 U11044 ( .A(P3_EAX_PTR14), .B(_02595__PTR14), .S(_02585_), .Z(_02674__PTR110) );
  MUX2_X1 U11045 ( .A(P3_EAX_PTR15), .B(_02595__PTR15), .S(_02585_), .Z(_02674__PTR111) );
  MUX2_X1 U11046 ( .A(P3_EAX_PTR16), .B(_02595__PTR16), .S(_02585_), .Z(_02674__PTR112) );
  MUX2_X1 U11047 ( .A(P3_EAX_PTR17), .B(_02595__PTR17), .S(_02585_), .Z(_02674__PTR113) );
  MUX2_X1 U11048 ( .A(P3_EAX_PTR18), .B(_02595__PTR18), .S(_02585_), .Z(_02674__PTR114) );
  MUX2_X1 U11049 ( .A(P3_EAX_PTR19), .B(_02595__PTR19), .S(_02585_), .Z(_02674__PTR115) );
  MUX2_X1 U11050 ( .A(P3_EAX_PTR20), .B(_02595__PTR20), .S(_02585_), .Z(_02674__PTR116) );
  MUX2_X1 U11051 ( .A(P3_EAX_PTR21), .B(_02595__PTR21), .S(_02585_), .Z(_02674__PTR117) );
  MUX2_X1 U11052 ( .A(P3_EAX_PTR22), .B(_02595__PTR22), .S(_02585_), .Z(_02674__PTR118) );
  MUX2_X1 U11053 ( .A(P3_EAX_PTR23), .B(_02595__PTR23), .S(_02585_), .Z(_02674__PTR119) );
  MUX2_X1 U11054 ( .A(P3_EAX_PTR24), .B(_02595__PTR24), .S(_02585_), .Z(_02674__PTR120) );
  MUX2_X1 U11055 ( .A(P3_EAX_PTR25), .B(_02595__PTR25), .S(_02585_), .Z(_02674__PTR121) );
  MUX2_X1 U11056 ( .A(P3_EAX_PTR26), .B(_02595__PTR26), .S(_02585_), .Z(_02674__PTR122) );
  MUX2_X1 U11057 ( .A(P3_EAX_PTR27), .B(_02595__PTR27), .S(_02585_), .Z(_02674__PTR123) );
  MUX2_X1 U11058 ( .A(P3_EAX_PTR28), .B(_02595__PTR28), .S(_02585_), .Z(_02674__PTR124) );
  MUX2_X1 U11059 ( .A(P3_EAX_PTR29), .B(_02595__PTR29), .S(_02585_), .Z(_02674__PTR125) );
  MUX2_X1 U11060 ( .A(P3_EAX_PTR30), .B(_02595__PTR30), .S(_02585_), .Z(_02674__PTR126) );
  MUX2_X1 U11061 ( .A(P3_EAX_PTR31), .B(_02595__PTR31), .S(_02585_), .Z(_02674__PTR127) );
  INV_X1 U11062 ( .A(_02458__PTR21), .ZN(_02458__PTR20) );
  MUX2_X1 U11063 ( .A(_02520__PTR2), .B(1'b0), .S(_02458__PTR21), .Z(_02458__PTR22) );
  INV_X1 U11064 ( .A(_02590_), .ZN(_02520__PTR2) );
  MUX2_X1 U11065 ( .A(_02661__PTR1), .B(1'b0), .S(_02627_), .Z(_02458__PTR16) );
  MUX2_X1 U11066 ( .A(_02661__PTR1), .B(1'b1), .S(_02627_), .Z(_02458__PTR17) );
  MUX2_X1 U11067 ( .A(_02661__PTR2), .B(1'b1), .S(_02627_), .Z(_02458__PTR18) );
  MUX2_X1 U11068 ( .A(na), .B(1'b1), .S(_02638_), .Z(_02661__PTR1) );
  MUX2_X1 U11069 ( .A(_02003_), .B(1'b1), .S(_02638_), .Z(_02661__PTR2) );
  MUX2_X1 U11070 ( .A(_02622__PTR0), .B(1'b0), .S(_01765__PTR4), .Z(_02458__PTR12) );
  MUX2_X1 U11071 ( .A(_02622__PTR1), .B(1'b1), .S(_01765__PTR4), .Z(_02458__PTR13) );
  MUX2_X1 U11072 ( .A(_02622__PTR2), .B(1'b0), .S(_01765__PTR4), .Z(_02458__PTR14) );
  MUX2_X1 U11073 ( .A(_02621__PTR0), .B(1'b0), .S(_02581_), .Z(_02622__PTR0) );
  MUX2_X1 U11074 ( .A(_02621__PTR1), .B(1'b0), .S(_02581_), .Z(_02622__PTR1) );
  MUX2_X1 U11075 ( .A(_02621__PTR2), .B(1'b0), .S(_02581_), .Z(_02622__PTR2) );
  MUX2_X1 U11076 ( .A(_02620__PTR0), .B(1'b1), .S(_02584_), .Z(_02621__PTR0) );
  MUX2_X1 U11077 ( .A(_02620__PTR1), .B(1'b1), .S(_02584_), .Z(_02621__PTR1) );
  MUX2_X1 U11078 ( .A(_02620__PTR2), .B(1'b1), .S(_02584_), .Z(_02621__PTR2) );
  INV_X1 U11079 ( .A(_02587_), .ZN(_02620__PTR0) );
  MUX2_X1 U11080 ( .A(_02619__PTR1), .B(1'b1), .S(_02587_), .Z(_02620__PTR1) );
  MUX2_X1 U11081 ( .A(_02619__PTR2), .B(1'b1), .S(_02587_), .Z(_02620__PTR2) );
  MUX2_X1 U11082 ( .A(_02618__PTR1), .B(1'b0), .S(_02591_), .Z(_02619__PTR1) );
  MUX2_X1 U11083 ( .A(_02600_), .B(1'b0), .S(_02591_), .Z(_02619__PTR2) );
  INV_X1 U11084 ( .A(_02600_), .ZN(_02618__PTR1) );
  INV_X1 U11085 ( .A(P3_CodeFetch), .ZN(_02424__PTR6) );
  INV_X1 U11086 ( .A(P3_ReadRequest), .ZN(_02428__PTR6) );
  INV_X1 U11087 ( .A(P3_RequestPending), .ZN(_02458__PTR4) );
  MUX2_X1 U11088 ( .A(hold), .B(1'b0), .S(P3_RequestPending), .Z(_02458__PTR6) );
  MUX2_X1 U11089 ( .A(1'b0), .B(_02126__PTR0), .S(_02929_), .Z(_02125__PTR0) );
  MUX2_X1 U11090 ( .A(1'b0), .B(_02126__PTR1), .S(_02929_), .Z(_02125__PTR1) );
  MUX2_X1 U11091 ( .A(1'b0), .B(_02126__PTR2), .S(_02929_), .Z(_02125__PTR2) );
  MUX2_X1 U11092 ( .A(1'b0), .B(_02126__PTR3), .S(_02929_), .Z(_02125__PTR3) );
  INV_X1 U11093 ( .A(_02750__PTR4), .ZN(_02752_) );
  INV_X1 U11094 ( .A(_02741__PTR5), .ZN(_02061_) );
  INV_X1 U11095 ( .A(_02729__PTR5), .ZN(_02730_) );
  INV_X1 U11096 ( .A(_02726__PTR5), .ZN(_02727_) );
  INV_X1 U11097 ( .A(_02719__PTR5), .ZN(_02721_) );
  INV_X1 U11098 ( .A(_02995__PTR4), .ZN(_02997_) );
  INV_X1 U11099 ( .A(_02986__PTR5), .ZN(_02350_) );
  INV_X1 U11100 ( .A(_02974__PTR5), .ZN(_02975_) );
  INV_X1 U11101 ( .A(_02971__PTR5), .ZN(_02972_) );
  INV_X1 U11102 ( .A(_02964__PTR5), .ZN(_02966_) );
  INV_X1 U11103 ( .A(_03240__PTR4), .ZN(_03242_) );
  INV_X1 U11104 ( .A(_03231__PTR5), .ZN(_02639_) );
  INV_X1 U11105 ( .A(_03219__PTR5), .ZN(_03220_) );
  INV_X1 U11106 ( .A(_03216__PTR5), .ZN(_03217_) );
  INV_X1 U11107 ( .A(_03209__PTR5), .ZN(_03211_) );
  INV_X1 U11108 ( .A(P3_Datao_PTR31), .ZN(_05728__PTR31) );
  INV_X1 U11109 ( .A(P2_Datao_PTR31), .ZN(_05724__PTR31) );
  INV_X1 U11110 ( .A(P1_Datao_PTR31), .ZN(_05720__PTR31) );
  INV_X1 U11111 ( .A(P2_Address_PTR0), .ZN(_05712__PTR0) );
  INV_X1 U11112 ( .A(P2_Address_PTR1), .ZN(_05712__PTR1) );
  INV_X1 U11113 ( .A(P2_Address_PTR2), .ZN(_05712__PTR2) );
  INV_X1 U11114 ( .A(P2_Address_PTR3), .ZN(_05712__PTR3) );
  INV_X1 U11115 ( .A(P2_Address_PTR4), .ZN(_05712__PTR4) );
  INV_X1 U11116 ( .A(P2_Address_PTR5), .ZN(_05712__PTR5) );
  INV_X1 U11117 ( .A(P2_Address_PTR6), .ZN(_05712__PTR6) );
  INV_X1 U11118 ( .A(P2_Address_PTR7), .ZN(_05712__PTR7) );
  INV_X1 U11119 ( .A(P2_Address_PTR8), .ZN(_05712__PTR8) );
  INV_X1 U11120 ( .A(P2_Address_PTR9), .ZN(_05712__PTR9) );
  INV_X1 U11121 ( .A(P2_Address_PTR10), .ZN(_05712__PTR10) );
  INV_X1 U11122 ( .A(P2_Address_PTR11), .ZN(_05712__PTR11) );
  INV_X1 U11123 ( .A(P2_Address_PTR12), .ZN(_05712__PTR12) );
  INV_X1 U11124 ( .A(P2_Address_PTR13), .ZN(_05712__PTR13) );
  INV_X1 U11125 ( .A(P2_Address_PTR14), .ZN(_05712__PTR14) );
  INV_X1 U11126 ( .A(P2_Address_PTR15), .ZN(_05712__PTR15) );
  INV_X1 U11127 ( .A(P2_Address_PTR16), .ZN(_05712__PTR16) );
  INV_X1 U11128 ( .A(P2_Address_PTR17), .ZN(_05712__PTR17) );
  INV_X1 U11129 ( .A(P2_Address_PTR18), .ZN(_05712__PTR18) );
  INV_X1 U11130 ( .A(P2_Address_PTR19), .ZN(_05712__PTR19) );
  INV_X1 U11131 ( .A(P2_Address_PTR20), .ZN(_05712__PTR20) );
  INV_X1 U11132 ( .A(P2_Address_PTR21), .ZN(_05712__PTR21) );
  INV_X1 U11133 ( .A(P2_Address_PTR22), .ZN(_05712__PTR22) );
  INV_X1 U11134 ( .A(P2_Address_PTR23), .ZN(_05712__PTR23) );
  INV_X1 U11135 ( .A(P2_Address_PTR24), .ZN(_05712__PTR24) );
  INV_X1 U11136 ( .A(P2_Address_PTR25), .ZN(_05712__PTR25) );
  INV_X1 U11137 ( .A(P2_Address_PTR26), .ZN(_05712__PTR26) );
  INV_X1 U11138 ( .A(P2_Address_PTR27), .ZN(_05712__PTR27) );
  INV_X1 U11139 ( .A(P2_Address_PTR28), .ZN(_05712__PTR28) );
  INV_X1 U11140 ( .A(P2_Address_PTR29), .ZN(_05712__PTR29) );
  INV_X1 U11141 ( .A(P1_Address_PTR0), .ZN(_05717__PTR0) );
  INV_X1 U11142 ( .A(P1_Address_PTR1), .ZN(_05717__PTR1) );
  INV_X1 U11143 ( .A(P1_Address_PTR2), .ZN(_05717__PTR2) );
  INV_X1 U11144 ( .A(P1_Address_PTR3), .ZN(_05717__PTR3) );
  INV_X1 U11145 ( .A(P1_Address_PTR4), .ZN(_05717__PTR4) );
  INV_X1 U11146 ( .A(P1_Address_PTR5), .ZN(_05717__PTR5) );
  INV_X1 U11147 ( .A(P1_Address_PTR6), .ZN(_05717__PTR6) );
  INV_X1 U11148 ( .A(P1_Address_PTR7), .ZN(_05717__PTR7) );
  INV_X1 U11149 ( .A(P1_Address_PTR8), .ZN(_05717__PTR8) );
  INV_X1 U11150 ( .A(P1_Address_PTR9), .ZN(_05717__PTR9) );
  INV_X1 U11151 ( .A(P1_Address_PTR10), .ZN(_05717__PTR10) );
  INV_X1 U11152 ( .A(P1_Address_PTR11), .ZN(_05717__PTR11) );
  INV_X1 U11153 ( .A(P1_Address_PTR12), .ZN(_05717__PTR12) );
  INV_X1 U11154 ( .A(P1_Address_PTR13), .ZN(_05717__PTR13) );
  INV_X1 U11155 ( .A(P1_Address_PTR14), .ZN(_05717__PTR14) );
  INV_X1 U11156 ( .A(P1_Address_PTR15), .ZN(_05717__PTR15) );
  INV_X1 U11157 ( .A(P1_Address_PTR16), .ZN(_05717__PTR16) );
  INV_X1 U11158 ( .A(P1_Address_PTR17), .ZN(_05717__PTR17) );
  INV_X1 U11159 ( .A(P1_Address_PTR18), .ZN(_05717__PTR18) );
  INV_X1 U11160 ( .A(P1_Address_PTR19), .ZN(_05717__PTR19) );
  INV_X1 U11161 ( .A(P1_Address_PTR20), .ZN(_05717__PTR20) );
  INV_X1 U11162 ( .A(P1_Address_PTR21), .ZN(_05717__PTR21) );
  INV_X1 U11163 ( .A(P1_Address_PTR22), .ZN(_05717__PTR22) );
  INV_X1 U11164 ( .A(P1_Address_PTR23), .ZN(_05717__PTR23) );
  INV_X1 U11165 ( .A(P1_Address_PTR24), .ZN(_05717__PTR24) );
  INV_X1 U11166 ( .A(P1_Address_PTR25), .ZN(_05717__PTR25) );
  INV_X1 U11167 ( .A(P1_Address_PTR26), .ZN(_05717__PTR26) );
  INV_X1 U11168 ( .A(P1_Address_PTR27), .ZN(_05717__PTR27) );
  INV_X1 U11169 ( .A(P1_Address_PTR28), .ZN(_05717__PTR28) );
  INV_X1 U11170 ( .A(P1_Address_PTR29), .ZN(_05717__PTR29) );
  INV_X1 U11171 ( .A(_01932__PTR56), .ZN(_02746__PTR0) );
  INV_X1 U11172 ( .A(_01932__PTR57), .ZN(_02746__PTR1) );
  INV_X1 U11173 ( .A(_01932__PTR58), .ZN(_02746__PTR2) );
  INV_X1 U11174 ( .A(_01932__PTR59), .ZN(_02746__PTR3) );
  INV_X1 U11175 ( .A(_01932__PTR60), .ZN(_02943__PTR4) );
  INV_X1 U11176 ( .A(P1_P1_InstAddrPointer_PTR31), .ZN(_02743__PTR31) );
  INV_X1 U11177 ( .A(_01932__PTR42), .ZN(_02739__PTR2) );
  INV_X1 U11178 ( .A(_01932__PTR43), .ZN(_02739__PTR3) );
  INV_X1 U11179 ( .A(_01932__PTR44), .ZN(_02941__PTR4) );
  INV_X1 U11180 ( .A(P1_P1_InstQueueWr_Addr_PTR1), .ZN(_02735__PTR1) );
  INV_X1 U11181 ( .A(P1_P1_InstQueueWr_Addr_PTR2), .ZN(_02735__PTR2) );
  INV_X1 U11182 ( .A(P1_P1_InstQueueWr_Addr_PTR3), .ZN(_02735__PTR3) );
  INV_X1 U11183 ( .A(P1_P1_InstQueueWr_Addr_PTR4), .ZN(_02735__PTR4) );
  INV_X1 U11184 ( .A(P1_EBX_PTR31), .ZN(_02732__PTR31) );
  INV_X1 U11185 ( .A(P1_P1_InstQueueRd_Addr_PTR3), .ZN(_02930__PTR3) );
  INV_X1 U11186 ( .A(P1_P1_InstQueueRd_Addr_PTR4), .ZN(_02751__PTR4) );
  INV_X1 U11187 ( .A(_01885__PTR7), .ZN(_02723__PTR7) );
  INV_X1 U11188 ( .A(_02725__PTR4), .ZN(_02936__PTR4) );
  INV_X1 U11189 ( .A(_02725__PTR5), .ZN(_02936__PTR5) );
  INV_X1 U11190 ( .A(_02725__PTR6), .ZN(_02936__PTR6) );
  INV_X1 U11191 ( .A(_02935__PTR7), .ZN(_02936__PTR7) );
  INV_X1 U11192 ( .A(_01885__PTR2), .ZN(_02723__PTR2) );
  INV_X1 U11193 ( .A(_01885__PTR3), .ZN(_02723__PTR3) );
  INV_X1 U11194 ( .A(_01885__PTR4), .ZN(_02723__PTR4) );
  INV_X1 U11195 ( .A(_01885__PTR5), .ZN(_02723__PTR5) );
  INV_X1 U11196 ( .A(_01885__PTR6), .ZN(_02723__PTR6) );
  INV_X1 U11197 ( .A(_02717__PTR1), .ZN(_02718__PTR1) );
  INV_X1 U11198 ( .A(_02717__PTR2), .ZN(_02718__PTR2) );
  INV_X1 U11199 ( .A(_02717__PTR3), .ZN(_02718__PTR3) );
  INV_X1 U11200 ( .A(_02717__PTR4), .ZN(_02718__PTR4) );
  INV_X1 U11201 ( .A(_01892__PTR159), .ZN(_02713__PTR31) );
  INV_X1 U11202 ( .A(P1_rEIP_PTR1), .ZN(_01882__PTR7) );
  INV_X1 U11203 ( .A(_02224__PTR56), .ZN(_02991__PTR0) );
  INV_X1 U11204 ( .A(_02224__PTR60), .ZN(_03188__PTR4) );
  INV_X1 U11205 ( .A(P2_P1_InstAddrPointer_PTR5), .ZN(_02990__PTR5) );
  INV_X1 U11206 ( .A(P2_P1_InstAddrPointer_PTR6), .ZN(_02990__PTR6) );
  INV_X1 U11207 ( .A(P2_P1_InstAddrPointer_PTR7), .ZN(_02990__PTR7) );
  INV_X1 U11208 ( .A(P2_P1_InstAddrPointer_PTR9), .ZN(_02990__PTR9) );
  INV_X1 U11209 ( .A(P2_P1_InstAddrPointer_PTR10), .ZN(_02990__PTR10) );
  INV_X1 U11210 ( .A(P2_P1_InstAddrPointer_PTR11), .ZN(_02990__PTR11) );
  INV_X1 U11211 ( .A(P2_P1_InstAddrPointer_PTR12), .ZN(_02990__PTR12) );
  INV_X1 U11212 ( .A(P2_P1_InstAddrPointer_PTR14), .ZN(_02990__PTR14) );
  INV_X1 U11213 ( .A(P2_P1_InstAddrPointer_PTR15), .ZN(_02990__PTR15) );
  INV_X1 U11214 ( .A(P2_P1_InstAddrPointer_PTR17), .ZN(_02990__PTR17) );
  INV_X1 U11215 ( .A(P2_P1_InstAddrPointer_PTR18), .ZN(_02990__PTR18) );
  INV_X1 U11216 ( .A(P2_P1_InstAddrPointer_PTR20), .ZN(_02990__PTR20) );
  INV_X1 U11217 ( .A(P2_P1_InstAddrPointer_PTR22), .ZN(_02990__PTR22) );
  INV_X1 U11218 ( .A(P2_P1_InstAddrPointer_PTR23), .ZN(_02990__PTR23) );
  INV_X1 U11219 ( .A(P2_P1_InstAddrPointer_PTR24), .ZN(_02990__PTR24) );
  INV_X1 U11220 ( .A(P2_P1_InstAddrPointer_PTR25), .ZN(_02990__PTR25) );
  INV_X1 U11221 ( .A(P2_P1_InstAddrPointer_PTR27), .ZN(_02990__PTR27) );
  INV_X1 U11222 ( .A(P2_P1_InstAddrPointer_PTR28), .ZN(_02990__PTR28) );
  INV_X1 U11223 ( .A(P2_P1_InstAddrPointer_PTR29), .ZN(_02990__PTR29) );
  INV_X1 U11224 ( .A(P2_P1_InstAddrPointer_PTR30), .ZN(_02990__PTR30) );
  INV_X1 U11225 ( .A(P2_P1_InstAddrPointer_PTR31), .ZN(_02988__PTR31) );
  INV_X1 U11226 ( .A(_02224__PTR42), .ZN(_02984__PTR2) );
  INV_X1 U11227 ( .A(_02224__PTR43), .ZN(_02984__PTR3) );
  INV_X1 U11228 ( .A(_02224__PTR44), .ZN(_03186__PTR4) );
  INV_X1 U11229 ( .A(P2_P1_InstQueueWr_Addr_PTR0), .ZN(_02129__PTR0) );
  INV_X1 U11230 ( .A(P2_P1_InstQueueWr_Addr_PTR1), .ZN(_02980__PTR1) );
  INV_X1 U11231 ( .A(P2_P1_InstQueueWr_Addr_PTR2), .ZN(_02980__PTR2) );
  INV_X1 U11232 ( .A(P2_P1_InstQueueWr_Addr_PTR3), .ZN(_02980__PTR3) );
  INV_X1 U11233 ( .A(P2_P1_InstQueueWr_Addr_PTR4), .ZN(_02980__PTR4) );
  INV_X1 U11234 ( .A(P2_EBX_PTR2), .ZN(_02979__PTR2) );
  INV_X1 U11235 ( .A(P2_EBX_PTR7), .ZN(_02979__PTR7) );
  INV_X1 U11236 ( .A(P2_EBX_PTR10), .ZN(_02979__PTR10) );
  INV_X1 U11237 ( .A(P2_EBX_PTR11), .ZN(_02979__PTR11) );
  INV_X1 U11238 ( .A(P2_EBX_PTR12), .ZN(_02979__PTR12) );
  INV_X1 U11239 ( .A(P2_EBX_PTR14), .ZN(_02979__PTR14) );
  INV_X1 U11240 ( .A(P2_EBX_PTR18), .ZN(_02979__PTR18) );
  INV_X1 U11241 ( .A(P2_EBX_PTR20), .ZN(_02979__PTR20) );
  INV_X1 U11242 ( .A(P2_EBX_PTR22), .ZN(_02979__PTR22) );
  INV_X1 U11243 ( .A(P2_EBX_PTR23), .ZN(_02979__PTR23) );
  INV_X1 U11244 ( .A(P2_EBX_PTR24), .ZN(_02979__PTR24) );
  INV_X1 U11245 ( .A(P2_EBX_PTR27), .ZN(_02979__PTR27) );
  INV_X1 U11246 ( .A(P2_EBX_PTR28), .ZN(_02979__PTR28) );
  INV_X1 U11247 ( .A(P2_EBX_PTR29), .ZN(_02979__PTR29) );
  INV_X1 U11248 ( .A(P2_EBX_PTR31), .ZN(_02977__PTR31) );
  INV_X1 U11249 ( .A(P2_P1_InstQueueRd_Addr_PTR1), .ZN(_02182__PTR4) );
  INV_X1 U11250 ( .A(P2_P1_InstQueueRd_Addr_PTR3), .ZN(_03175__PTR3) );
  INV_X1 U11251 ( .A(P2_P1_InstQueueRd_Addr_PTR4), .ZN(_02996__PTR4) );
  INV_X1 U11252 ( .A(_02962__PTR1), .ZN(_02963__PTR1) );
  INV_X1 U11253 ( .A(_02962__PTR2), .ZN(_02963__PTR2) );
  INV_X1 U11254 ( .A(_02177__PTR3), .ZN(_02968__PTR3) );
  INV_X1 U11255 ( .A(_02177__PTR7), .ZN(_02968__PTR7) );
  INV_X1 U11256 ( .A(_02962__PTR3), .ZN(_02963__PTR3) );
  INV_X1 U11257 ( .A(_02962__PTR4), .ZN(_02963__PTR4) );
  INV_X1 U11258 ( .A(_02177__PTR4), .ZN(_02968__PTR4) );
  INV_X1 U11259 ( .A(_02177__PTR5), .ZN(_02968__PTR5) );
  INV_X1 U11260 ( .A(_02970__PTR4), .ZN(_03181__PTR4) );
  INV_X1 U11261 ( .A(_02970__PTR5), .ZN(_03181__PTR5) );
  INV_X1 U11262 ( .A(_02970__PTR6), .ZN(_03181__PTR6) );
  INV_X1 U11263 ( .A(_03180__PTR7), .ZN(_03181__PTR7) );
  INV_X1 U11264 ( .A(_02177__PTR2), .ZN(_02968__PTR2) );
  INV_X1 U11265 ( .A(_02177__PTR6), .ZN(_02968__PTR6) );
  INV_X1 U11266 ( .A(P2_P1_PhyAddrPointer_PTR0), .ZN(_02960__PTR0) );
  INV_X1 U11267 ( .A(_02184__PTR132), .ZN(_02960__PTR4) );
  INV_X1 U11268 ( .A(_02184__PTR133), .ZN(_02960__PTR5) );
  INV_X1 U11269 ( .A(_02184__PTR136), .ZN(_02960__PTR8) );
  INV_X1 U11270 ( .A(_02184__PTR137), .ZN(_02960__PTR9) );
  INV_X1 U11271 ( .A(_02184__PTR139), .ZN(_02960__PTR11) );
  INV_X1 U11272 ( .A(_02184__PTR141), .ZN(_02960__PTR13) );
  INV_X1 U11273 ( .A(_02184__PTR143), .ZN(_02960__PTR15) );
  INV_X1 U11274 ( .A(_02184__PTR144), .ZN(_02960__PTR16) );
  INV_X1 U11275 ( .A(_02184__PTR149), .ZN(_02960__PTR21) );
  INV_X1 U11276 ( .A(_02184__PTR150), .ZN(_02960__PTR22) );
  INV_X1 U11277 ( .A(_02184__PTR151), .ZN(_02960__PTR23) );
  INV_X1 U11278 ( .A(_02184__PTR152), .ZN(_02960__PTR24) );
  INV_X1 U11279 ( .A(_02184__PTR153), .ZN(_02960__PTR25) );
  INV_X1 U11280 ( .A(_02184__PTR155), .ZN(_02960__PTR27) );
  INV_X1 U11281 ( .A(_02184__PTR156), .ZN(_02960__PTR28) );
  INV_X1 U11282 ( .A(_02184__PTR157), .ZN(_02960__PTR29) );
  INV_X1 U11283 ( .A(_02184__PTR159), .ZN(_02958__PTR31) );
  INV_X1 U11284 ( .A(_02513__PTR56), .ZN(_03236__PTR0) );
  INV_X1 U11285 ( .A(_02513__PTR57), .ZN(_03236__PTR1) );
  INV_X1 U11286 ( .A(_02513__PTR58), .ZN(_03236__PTR2) );
  INV_X1 U11287 ( .A(_02513__PTR60), .ZN(_03433__PTR4) );
  INV_X1 U11288 ( .A(P3_P1_InstAddrPointer_PTR2), .ZN(_03235__PTR2) );
  INV_X1 U11289 ( .A(P3_P1_InstAddrPointer_PTR3), .ZN(_03235__PTR3) );
  INV_X1 U11290 ( .A(P3_P1_InstAddrPointer_PTR5), .ZN(_03235__PTR5) );
  INV_X1 U11291 ( .A(P3_P1_InstAddrPointer_PTR6), .ZN(_03235__PTR6) );
  INV_X1 U11292 ( .A(P3_P1_InstAddrPointer_PTR8), .ZN(_03235__PTR8) );
  INV_X1 U11293 ( .A(P3_P1_InstAddrPointer_PTR9), .ZN(_03235__PTR9) );
  INV_X1 U11294 ( .A(P3_P1_InstAddrPointer_PTR12), .ZN(_03235__PTR12) );
  INV_X1 U11295 ( .A(P3_P1_InstAddrPointer_PTR13), .ZN(_03235__PTR13) );
  INV_X1 U11296 ( .A(P3_P1_InstAddrPointer_PTR14), .ZN(_03235__PTR14) );
  INV_X1 U11297 ( .A(P3_P1_InstAddrPointer_PTR15), .ZN(_03235__PTR15) );
  INV_X1 U11298 ( .A(P3_P1_InstAddrPointer_PTR16), .ZN(_03235__PTR16) );
  INV_X1 U11299 ( .A(P3_P1_InstAddrPointer_PTR18), .ZN(_03235__PTR18) );
  INV_X1 U11300 ( .A(P3_P1_InstAddrPointer_PTR19), .ZN(_03235__PTR19) );
  INV_X1 U11301 ( .A(P3_P1_InstAddrPointer_PTR23), .ZN(_03235__PTR23) );
  INV_X1 U11302 ( .A(P3_P1_InstAddrPointer_PTR24), .ZN(_03235__PTR24) );
  INV_X1 U11303 ( .A(P3_P1_InstAddrPointer_PTR25), .ZN(_03235__PTR25) );
  INV_X1 U11304 ( .A(P3_P1_InstAddrPointer_PTR26), .ZN(_03235__PTR26) );
  INV_X1 U11305 ( .A(P3_P1_InstAddrPointer_PTR27), .ZN(_03235__PTR27) );
  INV_X1 U11306 ( .A(P3_P1_InstAddrPointer_PTR29), .ZN(_03235__PTR29) );
  INV_X1 U11307 ( .A(P3_P1_InstAddrPointer_PTR30), .ZN(_03235__PTR30) );
  INV_X1 U11308 ( .A(P3_P1_InstAddrPointer_PTR31), .ZN(_03233__PTR31) );
  INV_X1 U11309 ( .A(_02513__PTR42), .ZN(_03229__PTR2) );
  INV_X1 U11310 ( .A(_02513__PTR43), .ZN(_03229__PTR3) );
  INV_X1 U11311 ( .A(_02513__PTR44), .ZN(_03431__PTR4) );
  INV_X1 U11312 ( .A(P3_P1_InstQueueWr_Addr_PTR0), .ZN(_02418__PTR0) );
  INV_X1 U11313 ( .A(P3_P1_InstQueueWr_Addr_PTR1), .ZN(_03225__PTR1) );
  INV_X1 U11314 ( .A(P3_P1_InstQueueWr_Addr_PTR2), .ZN(_03225__PTR2) );
  INV_X1 U11315 ( .A(P3_P1_InstQueueWr_Addr_PTR3), .ZN(_03225__PTR3) );
  INV_X1 U11316 ( .A(P3_P1_InstQueueWr_Addr_PTR4), .ZN(_03225__PTR4) );
  INV_X1 U11317 ( .A(P3_EBX_PTR1), .ZN(_03224__PTR1) );
  INV_X1 U11318 ( .A(P3_EBX_PTR4), .ZN(_03224__PTR4) );
  INV_X1 U11319 ( .A(P3_EBX_PTR5), .ZN(_03224__PTR5) );
  INV_X1 U11320 ( .A(P3_EBX_PTR6), .ZN(_03224__PTR6) );
  INV_X1 U11321 ( .A(P3_EBX_PTR7), .ZN(_03224__PTR7) );
  INV_X1 U11322 ( .A(P3_EBX_PTR8), .ZN(_03224__PTR8) );
  INV_X1 U11323 ( .A(P3_EBX_PTR9), .ZN(_03224__PTR9) );
  INV_X1 U11324 ( .A(P3_EBX_PTR10), .ZN(_03224__PTR10) );
  INV_X1 U11325 ( .A(P3_EBX_PTR11), .ZN(_03224__PTR11) );
  INV_X1 U11326 ( .A(P3_EBX_PTR12), .ZN(_03224__PTR12) );
  INV_X1 U11327 ( .A(P3_EBX_PTR13), .ZN(_03224__PTR13) );
  INV_X1 U11328 ( .A(P3_EBX_PTR14), .ZN(_03224__PTR14) );
  INV_X1 U11329 ( .A(P3_EBX_PTR15), .ZN(_03224__PTR15) );
  INV_X1 U11330 ( .A(P3_EBX_PTR16), .ZN(_03224__PTR16) );
  INV_X1 U11331 ( .A(P3_EBX_PTR17), .ZN(_03224__PTR17) );
  INV_X1 U11332 ( .A(P3_EBX_PTR18), .ZN(_03224__PTR18) );
  INV_X1 U11333 ( .A(P3_EBX_PTR19), .ZN(_03224__PTR19) );
  INV_X1 U11334 ( .A(P3_EBX_PTR21), .ZN(_03224__PTR21) );
  INV_X1 U11335 ( .A(P3_EBX_PTR22), .ZN(_03224__PTR22) );
  INV_X1 U11336 ( .A(P3_EBX_PTR23), .ZN(_03224__PTR23) );
  INV_X1 U11337 ( .A(P3_EBX_PTR24), .ZN(_03224__PTR24) );
  INV_X1 U11338 ( .A(P3_EBX_PTR25), .ZN(_03224__PTR25) );
  INV_X1 U11339 ( .A(P3_EBX_PTR26), .ZN(_03224__PTR26) );
  INV_X1 U11340 ( .A(P3_EBX_PTR27), .ZN(_03224__PTR27) );
  INV_X1 U11341 ( .A(P3_EBX_PTR28), .ZN(_03224__PTR28) );
  INV_X1 U11342 ( .A(P3_EBX_PTR29), .ZN(_03224__PTR29) );
  INV_X1 U11343 ( .A(P3_EBX_PTR30), .ZN(_03224__PTR30) );
  INV_X1 U11344 ( .A(P3_EBX_PTR31), .ZN(_03222__PTR31) );
  INV_X1 U11345 ( .A(P3_P1_InstQueueRd_Addr_PTR3), .ZN(_03420__PTR3) );
  INV_X1 U11346 ( .A(P3_P1_InstQueueRd_Addr_PTR4), .ZN(_03241__PTR4) );
  INV_X1 U11347 ( .A(_02466__PTR2), .ZN(_03213__PTR2) );
  INV_X1 U11348 ( .A(_02466__PTR3), .ZN(_03213__PTR3) );
  INV_X1 U11349 ( .A(_02466__PTR4), .ZN(_03213__PTR4) );
  INV_X1 U11350 ( .A(_02466__PTR5), .ZN(_03213__PTR5) );
  INV_X1 U11351 ( .A(_02466__PTR7), .ZN(_03213__PTR7) );
  INV_X1 U11352 ( .A(_03207__PTR1), .ZN(_03208__PTR1) );
  INV_X1 U11353 ( .A(_03207__PTR2), .ZN(_03208__PTR2) );
  INV_X1 U11354 ( .A(_03207__PTR3), .ZN(_03208__PTR3) );
  INV_X1 U11355 ( .A(_03207__PTR4), .ZN(_03208__PTR4) );
  INV_X1 U11356 ( .A(_02466__PTR6), .ZN(_03213__PTR6) );
  INV_X1 U11357 ( .A(_03215__PTR4), .ZN(_03426__PTR4) );
  INV_X1 U11358 ( .A(_03215__PTR5), .ZN(_03426__PTR5) );
  INV_X1 U11359 ( .A(_03215__PTR6), .ZN(_03426__PTR6) );
  INV_X1 U11360 ( .A(_03425__PTR7), .ZN(_03426__PTR7) );
  INV_X1 U11361 ( .A(_02473__PTR130), .ZN(_03205__PTR2) );
  INV_X1 U11362 ( .A(_02473__PTR134), .ZN(_03205__PTR6) );
  INV_X1 U11363 ( .A(_02473__PTR135), .ZN(_03205__PTR7) );
  INV_X1 U11364 ( .A(_02473__PTR136), .ZN(_03205__PTR8) );
  INV_X1 U11365 ( .A(_02473__PTR137), .ZN(_03205__PTR9) );
  INV_X1 U11366 ( .A(_02473__PTR138), .ZN(_03205__PTR10) );
  INV_X1 U11367 ( .A(_02473__PTR139), .ZN(_03205__PTR11) );
  INV_X1 U11368 ( .A(_02473__PTR140), .ZN(_03205__PTR12) );
  INV_X1 U11369 ( .A(_02473__PTR141), .ZN(_03205__PTR13) );
  INV_X1 U11370 ( .A(_02473__PTR142), .ZN(_03205__PTR14) );
  INV_X1 U11371 ( .A(_02473__PTR143), .ZN(_03205__PTR15) );
  INV_X1 U11372 ( .A(_02473__PTR144), .ZN(_03205__PTR16) );
  INV_X1 U11373 ( .A(_02473__PTR145), .ZN(_03205__PTR17) );
  INV_X1 U11374 ( .A(_02473__PTR146), .ZN(_03205__PTR18) );
  INV_X1 U11375 ( .A(_02473__PTR147), .ZN(_03205__PTR19) );
  INV_X1 U11376 ( .A(_02473__PTR148), .ZN(_03205__PTR20) );
  INV_X1 U11377 ( .A(_02473__PTR149), .ZN(_03205__PTR21) );
  INV_X1 U11378 ( .A(_02473__PTR150), .ZN(_03205__PTR22) );
  INV_X1 U11379 ( .A(_02473__PTR151), .ZN(_03205__PTR23) );
  INV_X1 U11380 ( .A(_02473__PTR152), .ZN(_03205__PTR24) );
  INV_X1 U11381 ( .A(_02473__PTR153), .ZN(_03205__PTR25) );
  INV_X1 U11382 ( .A(_02473__PTR154), .ZN(_03205__PTR26) );
  INV_X1 U11383 ( .A(_02473__PTR155), .ZN(_03205__PTR27) );
  INV_X1 U11384 ( .A(_02473__PTR156), .ZN(_03205__PTR28) );
  INV_X1 U11385 ( .A(_02473__PTR157), .ZN(_03205__PTR29) );
  INV_X1 U11386 ( .A(_02473__PTR158), .ZN(_03205__PTR30) );
  INV_X1 U11387 ( .A(_02473__PTR159), .ZN(_03203__PTR31) );
  INV_X1 U11388 ( .A(P1_ADS_n), .ZN(_05753_) );
  INV_X1 U11389 ( .A(P1_D_C_n), .ZN(_05754_) );
  INV_X1 U11390 ( .A(P2_ADS_n), .ZN(_05763_) );
  INV_X1 U11391 ( .A(P2_D_C_n), .ZN(_05764_) );
  INV_X1 U11392 ( .A(P3_ADS_n), .ZN(_05742_) );
  INV_X1 U11393 ( .A(P3_D_C_n), .ZN(_05743_) );
  INV_X1 U11394 ( .A(P3_W_R_n), .ZN(_05744_) );
  INV_X1 U11395 ( .A(_00135_), .ZN(_02124__PTR0) );
  INV_X1 U11396 ( .A(_01834_), .ZN(_02058_) );
  INV_X1 U11397 ( .A(P1_StateBS16), .ZN(_01894__PTR9) );
  INV_X1 U11398 ( .A(P1_READY_n), .ZN(_01894__PTR14) );
  INV_X1 U11399 ( .A(_01770__PTR2), .ZN(_01894__PTR32) );
  INV_X1 U11400 ( .A(_01853__PTR2), .ZN(_01857__PTR2) );
  INV_X1 U11401 ( .A(_01853__PTR3), .ZN(_01857__PTR3) );
  INV_X1 U11402 ( .A(_00136_), .ZN(_02413__PTR0) );
  INV_X1 U11403 ( .A(_02127_), .ZN(_02347_) );
  INV_X1 U11404 ( .A(P2_StateBS16), .ZN(_02186__PTR9) );
  INV_X1 U11405 ( .A(P2_READY_n), .ZN(_02186__PTR14) );
  INV_X1 U11406 ( .A(_01768__PTR2), .ZN(_02186__PTR32) );
  INV_X1 U11407 ( .A(_02146__PTR2), .ZN(_02150__PTR2) );
  INV_X1 U11408 ( .A(_02146__PTR3), .ZN(_02150__PTR3) );
  INV_X1 U11409 ( .A(na), .ZN(_02003_) );
  INV_X1 U11410 ( .A(hold), .ZN(_01999_) );
  INV_X1 U11411 ( .A(_00137_), .ZN(_02702__PTR0) );
  INV_X1 U11412 ( .A(_02416_), .ZN(_02636_) );
  INV_X1 U11413 ( .A(P3_StateBS16), .ZN(_02475__PTR9) );
  INV_X1 U11414 ( .A(P3_READY_n), .ZN(_02475__PTR14) );
  INV_X1 U11415 ( .A(_01766__PTR2), .ZN(_02475__PTR32) );
  INV_X1 U11416 ( .A(_02435__PTR2), .ZN(_02439__PTR2) );
  INV_X1 U11417 ( .A(_02435__PTR3), .ZN(_02439__PTR3) );
  INV_X1 U11418 ( .A(_05729__PTR31), .ZN(_05731_) );
  INV_X1 U11419 ( .A(_05725__PTR31), .ZN(_05727_) );
  INV_X1 U11420 ( .A(_05721__PTR31), .ZN(_05723_) );
  INV_X1 U11421 ( .A(_05715__PTR29), .ZN(_05716_) );
  INV_X1 U11422 ( .A(_05713__PTR29), .ZN(_05714_) );
  INV_X1 U11423 ( .A(_05718__PTR29), .ZN(_05719_) );
  DFFR_X1 ready11 ( .D(_05734_), .CK(clock), .RN(reset_n_DEFINE), .Q(ready11), .QN());
  DFFR_X1 ready12 ( .D(_05736_), .CK(clock), .RN(reset_n_DEFINE), .Q(ready12), .QN());
  DFFR_X1 ready21 ( .D(_05750_), .CK(clock), .RN(reset_n_DEFINE), .Q(ready21), .QN());
  DFFR_X1 ready22 ( .D(_05752_), .CK(clock), .RN(reset_n_DEFINE), .Q(ready22), .QN());
  DFFR_X1 P2_ByteEnable_PTR0 ( .D(_02414__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_ByteEnable_PTR0), .QN());
  DFFR_X1 P2_ByteEnable_PTR1 ( .D(_02414__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_ByteEnable_PTR1), .QN());
  DFFR_X1 P2_ByteEnable_PTR2 ( .D(_02414__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_ByteEnable_PTR2), .QN());
  DFFR_X1 P2_ByteEnable_PTR3 ( .D(_02414__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P2_ByteEnable_PTR3), .QN());
  DFFR_X1 buf2_PTR0 ( .D(P2_Datao_PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR0), .QN());
  DFFR_X1 buf2_PTR1 ( .D(P2_Datao_PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR1), .QN());
  DFFR_X1 buf2_PTR2 ( .D(P2_Datao_PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR2), .QN());
  DFFR_X1 buf2_PTR3 ( .D(P2_Datao_PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR3), .QN());
  DFFR_X1 buf2_PTR4 ( .D(P2_Datao_PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR4), .QN());
  DFFR_X1 buf2_PTR5 ( .D(P2_Datao_PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR5), .QN());
  DFFR_X1 buf2_PTR6 ( .D(P2_Datao_PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR6), .QN());
  DFFR_X1 buf2_PTR7 ( .D(P2_Datao_PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR7), .QN());
  DFFR_X1 buf2_PTR8 ( .D(P2_Datao_PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR8), .QN());
  DFFR_X1 buf2_PTR9 ( .D(P2_Datao_PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR9), .QN());
  DFFR_X1 buf2_PTR10 ( .D(P2_Datao_PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR10), .QN());
  DFFR_X1 buf2_PTR11 ( .D(P2_Datao_PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR11), .QN());
  DFFR_X1 buf2_PTR12 ( .D(P2_Datao_PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR12), .QN());
  DFFR_X1 buf2_PTR13 ( .D(P2_Datao_PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR13), .QN());
  DFFR_X1 buf2_PTR14 ( .D(P2_Datao_PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR14), .QN());
  DFFR_X1 buf2_PTR15 ( .D(P2_Datao_PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR15), .QN());
  DFFR_X1 buf2_PTR16 ( .D(P2_Datao_PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR16), .QN());
  DFFR_X1 buf2_PTR17 ( .D(P2_Datao_PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR17), .QN());
  DFFR_X1 buf2_PTR18 ( .D(P2_Datao_PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR18), .QN());
  DFFR_X1 buf2_PTR19 ( .D(P2_Datao_PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR19), .QN());
  DFFR_X1 buf2_PTR20 ( .D(P2_Datao_PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR20), .QN());
  DFFR_X1 buf2_PTR21 ( .D(P2_Datao_PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR21), .QN());
  DFFR_X1 buf2_PTR22 ( .D(P2_Datao_PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR22), .QN());
  DFFR_X1 buf2_PTR23 ( .D(P2_Datao_PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR23), .QN());
  DFFR_X1 buf2_PTR24 ( .D(P2_Datao_PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR24), .QN());
  DFFR_X1 buf2_PTR25 ( .D(P2_Datao_PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR25), .QN());
  DFFR_X1 buf2_PTR26 ( .D(P2_Datao_PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR26), .QN());
  DFFR_X1 buf2_PTR27 ( .D(P2_Datao_PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR27), .QN());
  DFFR_X1 buf2_PTR28 ( .D(P2_Datao_PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR28), .QN());
  DFFR_X1 buf2_PTR29 ( .D(P2_Datao_PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR29), .QN());
  DFFR_X1 buf2_PTR30 ( .D(P2_Datao_PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR30), .QN());
  DFFR_X1 buf2_PTR31 ( .D(P2_Datao_PTR31), .CK(clock), .RN(reset_n_DEFINE), .Q(buf2_PTR31), .QN());
  DFFR_X1 buf1_PTR0 ( .D(_05733__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR0), .QN());
  DFFR_X1 buf1_PTR1 ( .D(_05733__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR1), .QN());
  DFFR_X1 buf1_PTR2 ( .D(_05733__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR2), .QN());
  DFFR_X1 buf1_PTR3 ( .D(_05733__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR3), .QN());
  DFFR_X1 buf1_PTR4 ( .D(_05733__PTR4), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR4), .QN());
  DFFR_X1 buf1_PTR5 ( .D(_05733__PTR5), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR5), .QN());
  DFFR_X1 buf1_PTR6 ( .D(_05733__PTR6), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR6), .QN());
  DFFR_X1 buf1_PTR7 ( .D(_05733__PTR7), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR7), .QN());
  DFFR_X1 buf1_PTR8 ( .D(_05733__PTR8), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR8), .QN());
  DFFR_X1 buf1_PTR9 ( .D(_05733__PTR9), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR9), .QN());
  DFFR_X1 buf1_PTR10 ( .D(_05733__PTR10), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR10), .QN());
  DFFR_X1 buf1_PTR11 ( .D(_05733__PTR11), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR11), .QN());
  DFFR_X1 buf1_PTR12 ( .D(_05733__PTR12), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR12), .QN());
  DFFR_X1 buf1_PTR13 ( .D(_05733__PTR13), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR13), .QN());
  DFFR_X1 buf1_PTR14 ( .D(_05733__PTR14), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR14), .QN());
  DFFR_X1 buf1_PTR15 ( .D(_05733__PTR15), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR15), .QN());
  DFFR_X1 buf1_PTR16 ( .D(_05733__PTR16), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR16), .QN());
  DFFR_X1 buf1_PTR17 ( .D(_05733__PTR17), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR17), .QN());
  DFFR_X1 buf1_PTR18 ( .D(_05733__PTR18), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR18), .QN());
  DFFR_X1 buf1_PTR19 ( .D(_05733__PTR19), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR19), .QN());
  DFFR_X1 buf1_PTR20 ( .D(_05733__PTR20), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR20), .QN());
  DFFR_X1 buf1_PTR21 ( .D(_05733__PTR21), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR21), .QN());
  DFFR_X1 buf1_PTR22 ( .D(_05733__PTR22), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR22), .QN());
  DFFR_X1 buf1_PTR23 ( .D(_05733__PTR23), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR23), .QN());
  DFFR_X1 buf1_PTR24 ( .D(_05733__PTR24), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR24), .QN());
  DFFR_X1 buf1_PTR25 ( .D(_05733__PTR25), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR25), .QN());
  DFFR_X1 buf1_PTR26 ( .D(_05733__PTR26), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR26), .QN());
  DFFR_X1 buf1_PTR27 ( .D(_05733__PTR27), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR27), .QN());
  DFFR_X1 buf1_PTR28 ( .D(_05733__PTR28), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR28), .QN());
  DFFR_X1 buf1_PTR29 ( .D(_05733__PTR29), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR29), .QN());
  DFFR_X1 buf1_PTR30 ( .D(_05733__PTR30), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR30), .QN());
  DFFR_X1 buf1_PTR31 ( .D(_05733__PTR31), .CK(clock), .RN(reset_n_DEFINE), .Q(buf1_PTR31), .QN());
  DFFR_X1 P1_ByteEnable_PTR0 ( .D(_02125__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_ByteEnable_PTR0), .QN());
  DFFR_X1 P1_ByteEnable_PTR1 ( .D(_02125__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_ByteEnable_PTR1), .QN());
  DFFR_X1 P1_ByteEnable_PTR2 ( .D(_02125__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_ByteEnable_PTR2), .QN());
  DFFR_X1 P1_ByteEnable_PTR3 ( .D(_02125__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P1_ByteEnable_PTR3), .QN());
  DFFR_X1 P3_ByteEnable_PTR0 ( .D(_02703__PTR0), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_ByteEnable_PTR0), .QN());
  DFFR_X1 P3_ByteEnable_PTR1 ( .D(_02703__PTR1), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_ByteEnable_PTR1), .QN());
  DFFR_X1 P3_ByteEnable_PTR2 ( .D(_02703__PTR2), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_ByteEnable_PTR2), .QN());
  DFFR_X1 P3_ByteEnable_PTR3 ( .D(_02703__PTR3), .CK(clock), .RN(reset_n_DEFINE), .Q(P3_ByteEnable_PTR3), .QN());
  AND2_X1 U11424 ( .A1(_02114__PTR64), .A2(_01863__PTR2), .ZN(_02115__PTR64) );
  AND2_X1 U11425 ( .A1(_02114__PTR65), .A2(_01863__PTR2), .ZN(_02115__PTR65) );
  AND2_X1 U11426 ( .A1(_02114__PTR66), .A2(_01863__PTR2), .ZN(_02115__PTR66) );
  AND2_X1 U11427 ( .A1(_02114__PTR67), .A2(_01863__PTR2), .ZN(_02115__PTR67) );
  AND2_X1 U11428 ( .A1(_02114__PTR68), .A2(_01863__PTR2), .ZN(_02115__PTR68) );
  AND2_X1 U11429 ( .A1(_02114__PTR69), .A2(_01863__PTR2), .ZN(_02115__PTR69) );
  AND2_X1 U11430 ( .A1(_02114__PTR70), .A2(_01863__PTR2), .ZN(_02115__PTR70) );
  AND2_X1 U11431 ( .A1(_02114__PTR71), .A2(_01863__PTR2), .ZN(_02115__PTR71) );
  AND2_X1 U11432 ( .A1(_02114__PTR72), .A2(_01863__PTR2), .ZN(_02115__PTR72) );
  AND2_X1 U11433 ( .A1(_02114__PTR73), .A2(_01863__PTR2), .ZN(_02115__PTR73) );
  AND2_X1 U11434 ( .A1(_02114__PTR74), .A2(_01863__PTR2), .ZN(_02115__PTR74) );
  AND2_X1 U11435 ( .A1(_02114__PTR75), .A2(_01863__PTR2), .ZN(_02115__PTR75) );
  AND2_X1 U11436 ( .A1(_02114__PTR76), .A2(_01863__PTR2), .ZN(_02115__PTR76) );
  AND2_X1 U11437 ( .A1(_02114__PTR77), .A2(_01863__PTR2), .ZN(_02115__PTR77) );
  AND2_X1 U11438 ( .A1(_02114__PTR78), .A2(_01863__PTR2), .ZN(_02115__PTR78) );
  AND2_X1 U11439 ( .A1(_02114__PTR79), .A2(_01863__PTR2), .ZN(_02115__PTR79) );
  AND2_X1 U11440 ( .A1(_02114__PTR80), .A2(_01863__PTR2), .ZN(_02115__PTR80) );
  AND2_X1 U11441 ( .A1(_02114__PTR81), .A2(_01863__PTR2), .ZN(_02115__PTR81) );
  AND2_X1 U11442 ( .A1(_02114__PTR82), .A2(_01863__PTR2), .ZN(_02115__PTR82) );
  AND2_X1 U11443 ( .A1(_02114__PTR83), .A2(_01863__PTR2), .ZN(_02115__PTR83) );
  AND2_X1 U11444 ( .A1(_02114__PTR84), .A2(_01863__PTR2), .ZN(_02115__PTR84) );
  AND2_X1 U11445 ( .A1(_02114__PTR85), .A2(_01863__PTR2), .ZN(_02115__PTR85) );
  AND2_X1 U11446 ( .A1(_02114__PTR86), .A2(_01863__PTR2), .ZN(_02115__PTR86) );
  AND2_X1 U11447 ( .A1(_02114__PTR87), .A2(_01863__PTR2), .ZN(_02115__PTR87) );
  AND2_X1 U11448 ( .A1(_02114__PTR88), .A2(_01863__PTR2), .ZN(_02115__PTR88) );
  AND2_X1 U11449 ( .A1(_02114__PTR89), .A2(_01863__PTR2), .ZN(_02115__PTR89) );
  AND2_X1 U11450 ( .A1(_02114__PTR90), .A2(_01863__PTR2), .ZN(_02115__PTR90) );
  AND2_X1 U11451 ( .A1(_02114__PTR91), .A2(_01863__PTR2), .ZN(_02115__PTR91) );
  AND2_X1 U11452 ( .A1(_02114__PTR92), .A2(_01863__PTR2), .ZN(_02115__PTR92) );
  AND2_X1 U11453 ( .A1(_02114__PTR93), .A2(_01863__PTR2), .ZN(_02115__PTR93) );
  AND2_X1 U11454 ( .A1(_02114__PTR94), .A2(_01863__PTR2), .ZN(_02115__PTR94) );
  AND2_X1 U11455 ( .A1(_02114__PTR95), .A2(_01863__PTR2), .ZN(_02115__PTR95) );
  AND2_X1 U11456 ( .A1(_02114__PTR64), .A2(_01863__PTR0), .ZN(_02115__PTR32) );
  AND2_X1 U11457 ( .A1(_02114__PTR65), .A2(_01863__PTR0), .ZN(_02115__PTR33) );
  AND2_X1 U11458 ( .A1(_02114__PTR66), .A2(_01863__PTR0), .ZN(_02115__PTR34) );
  AND2_X1 U11459 ( .A1(_02114__PTR67), .A2(_01863__PTR0), .ZN(_02115__PTR35) );
  AND2_X1 U11460 ( .A1(_02114__PTR68), .A2(_01863__PTR0), .ZN(_02115__PTR36) );
  AND2_X1 U11461 ( .A1(_02114__PTR69), .A2(_01863__PTR0), .ZN(_02115__PTR37) );
  AND2_X1 U11462 ( .A1(_02114__PTR70), .A2(_01863__PTR0), .ZN(_02115__PTR38) );
  AND2_X1 U11463 ( .A1(_02114__PTR71), .A2(_01863__PTR0), .ZN(_02115__PTR39) );
  AND2_X1 U11464 ( .A1(_02114__PTR72), .A2(_01863__PTR0), .ZN(_02115__PTR40) );
  AND2_X1 U11465 ( .A1(_02114__PTR73), .A2(_01863__PTR0), .ZN(_02115__PTR41) );
  AND2_X1 U11466 ( .A1(_02114__PTR74), .A2(_01863__PTR0), .ZN(_02115__PTR42) );
  AND2_X1 U11467 ( .A1(_02114__PTR75), .A2(_01863__PTR0), .ZN(_02115__PTR43) );
  AND2_X1 U11468 ( .A1(_02114__PTR76), .A2(_01863__PTR0), .ZN(_02115__PTR44) );
  AND2_X1 U11469 ( .A1(_02114__PTR77), .A2(_01863__PTR0), .ZN(_02115__PTR45) );
  AND2_X1 U11470 ( .A1(_02114__PTR78), .A2(_01863__PTR0), .ZN(_02115__PTR46) );
  AND2_X1 U11471 ( .A1(_02114__PTR79), .A2(_01863__PTR0), .ZN(_02115__PTR47) );
  AND2_X1 U11472 ( .A1(_02114__PTR48), .A2(_01863__PTR0), .ZN(_02115__PTR48) );
  AND2_X1 U11473 ( .A1(_02114__PTR49), .A2(_01863__PTR0), .ZN(_02115__PTR49) );
  AND2_X1 U11474 ( .A1(_02114__PTR50), .A2(_01863__PTR0), .ZN(_02115__PTR50) );
  AND2_X1 U11475 ( .A1(_02114__PTR51), .A2(_01863__PTR0), .ZN(_02115__PTR51) );
  AND2_X1 U11476 ( .A1(_02114__PTR52), .A2(_01863__PTR0), .ZN(_02115__PTR52) );
  AND2_X1 U11477 ( .A1(_02114__PTR53), .A2(_01863__PTR0), .ZN(_02115__PTR53) );
  AND2_X1 U11478 ( .A1(_02114__PTR54), .A2(_01863__PTR0), .ZN(_02115__PTR54) );
  AND2_X1 U11479 ( .A1(_02114__PTR55), .A2(_01863__PTR0), .ZN(_02115__PTR55) );
  AND2_X1 U11480 ( .A1(_02114__PTR56), .A2(_01863__PTR0), .ZN(_02115__PTR56) );
  AND2_X1 U11481 ( .A1(_02114__PTR57), .A2(_01863__PTR0), .ZN(_02115__PTR57) );
  AND2_X1 U11482 ( .A1(_02114__PTR58), .A2(_01863__PTR0), .ZN(_02115__PTR58) );
  AND2_X1 U11483 ( .A1(_02114__PTR59), .A2(_01863__PTR0), .ZN(_02115__PTR59) );
  AND2_X1 U11484 ( .A1(_02114__PTR60), .A2(_01863__PTR0), .ZN(_02115__PTR60) );
  AND2_X1 U11485 ( .A1(_02114__PTR61), .A2(_01863__PTR0), .ZN(_02115__PTR61) );
  AND2_X1 U11486 ( .A1(_02114__PTR62), .A2(_01863__PTR0), .ZN(_02115__PTR62) );
  AND2_X1 U11487 ( .A1(_02114__PTR95), .A2(_01863__PTR0), .ZN(_02115__PTR63) );
  AND2_X1 U11488 ( .A1(P1_Datao_PTR0), .A2(_02116__PTR0), .ZN(_02115__PTR0) );
  AND2_X1 U11489 ( .A1(P1_Datao_PTR1), .A2(_02116__PTR0), .ZN(_02115__PTR1) );
  AND2_X1 U11490 ( .A1(P1_Datao_PTR2), .A2(_02116__PTR0), .ZN(_02115__PTR2) );
  AND2_X1 U11491 ( .A1(P1_Datao_PTR3), .A2(_02116__PTR0), .ZN(_02115__PTR3) );
  AND2_X1 U11492 ( .A1(P1_Datao_PTR4), .A2(_02116__PTR0), .ZN(_02115__PTR4) );
  AND2_X1 U11493 ( .A1(P1_Datao_PTR5), .A2(_02116__PTR0), .ZN(_02115__PTR5) );
  AND2_X1 U11494 ( .A1(P1_Datao_PTR6), .A2(_02116__PTR0), .ZN(_02115__PTR6) );
  AND2_X1 U11495 ( .A1(P1_Datao_PTR7), .A2(_02116__PTR0), .ZN(_02115__PTR7) );
  AND2_X1 U11496 ( .A1(P1_Datao_PTR8), .A2(_02116__PTR0), .ZN(_02115__PTR8) );
  AND2_X1 U11497 ( .A1(P1_Datao_PTR9), .A2(_02116__PTR0), .ZN(_02115__PTR9) );
  AND2_X1 U11498 ( .A1(P1_Datao_PTR10), .A2(_02116__PTR0), .ZN(_02115__PTR10) );
  AND2_X1 U11499 ( .A1(P1_Datao_PTR11), .A2(_02116__PTR0), .ZN(_02115__PTR11) );
  AND2_X1 U11500 ( .A1(P1_Datao_PTR12), .A2(_02116__PTR0), .ZN(_02115__PTR12) );
  AND2_X1 U11501 ( .A1(P1_Datao_PTR13), .A2(_02116__PTR0), .ZN(_02115__PTR13) );
  AND2_X1 U11502 ( .A1(P1_Datao_PTR14), .A2(_02116__PTR0), .ZN(_02115__PTR14) );
  AND2_X1 U11503 ( .A1(P1_Datao_PTR15), .A2(_02116__PTR0), .ZN(_02115__PTR15) );
  AND2_X1 U11504 ( .A1(P1_Datao_PTR16), .A2(_02116__PTR0), .ZN(_02115__PTR16) );
  AND2_X1 U11505 ( .A1(P1_Datao_PTR17), .A2(_02116__PTR0), .ZN(_02115__PTR17) );
  AND2_X1 U11506 ( .A1(P1_Datao_PTR18), .A2(_02116__PTR0), .ZN(_02115__PTR18) );
  AND2_X1 U11507 ( .A1(P1_Datao_PTR19), .A2(_02116__PTR0), .ZN(_02115__PTR19) );
  AND2_X1 U11508 ( .A1(P1_Datao_PTR20), .A2(_02116__PTR0), .ZN(_02115__PTR20) );
  AND2_X1 U11509 ( .A1(P1_Datao_PTR21), .A2(_02116__PTR0), .ZN(_02115__PTR21) );
  AND2_X1 U11510 ( .A1(P1_Datao_PTR22), .A2(_02116__PTR0), .ZN(_02115__PTR22) );
  AND2_X1 U11511 ( .A1(P1_Datao_PTR23), .A2(_02116__PTR0), .ZN(_02115__PTR23) );
  AND2_X1 U11512 ( .A1(P1_Datao_PTR24), .A2(_02116__PTR0), .ZN(_02115__PTR24) );
  AND2_X1 U11513 ( .A1(P1_Datao_PTR25), .A2(_02116__PTR0), .ZN(_02115__PTR25) );
  AND2_X1 U11514 ( .A1(P1_Datao_PTR26), .A2(_02116__PTR0), .ZN(_02115__PTR26) );
  AND2_X1 U11515 ( .A1(P1_Datao_PTR27), .A2(_02116__PTR0), .ZN(_02115__PTR27) );
  AND2_X1 U11516 ( .A1(P1_Datao_PTR28), .A2(_02116__PTR0), .ZN(_02115__PTR28) );
  AND2_X1 U11517 ( .A1(P1_Datao_PTR29), .A2(_02116__PTR0), .ZN(_02115__PTR29) );
  AND2_X1 U11518 ( .A1(P1_Datao_PTR30), .A2(_02116__PTR0), .ZN(_02115__PTR30) );
  AND2_X1 U11519 ( .A1(P1_Datao_PTR31), .A2(_02116__PTR0), .ZN(_02115__PTR31) );
  AND2_X1 U11520 ( .A1(_02111__PTR32), .A2(_02090__PTR4), .ZN(_02112__PTR32) );
  AND2_X1 U11521 ( .A1(_02111__PTR33), .A2(_02090__PTR4), .ZN(_02112__PTR33) );
  AND2_X1 U11522 ( .A1(_02111__PTR34), .A2(_02090__PTR4), .ZN(_02112__PTR34) );
  AND2_X1 U11523 ( .A1(_02111__PTR35), .A2(_02090__PTR4), .ZN(_02112__PTR35) );
  AND2_X1 U11524 ( .A1(_02111__PTR36), .A2(_02090__PTR4), .ZN(_02112__PTR36) );
  AND2_X1 U11525 ( .A1(_02111__PTR37), .A2(_02090__PTR4), .ZN(_02112__PTR37) );
  AND2_X1 U11526 ( .A1(_02111__PTR38), .A2(_02090__PTR4), .ZN(_02112__PTR38) );
  AND2_X1 U11527 ( .A1(_02111__PTR39), .A2(_02090__PTR4), .ZN(_02112__PTR39) );
  AND2_X1 U11528 ( .A1(_02111__PTR40), .A2(_02090__PTR4), .ZN(_02112__PTR40) );
  AND2_X1 U11529 ( .A1(_02111__PTR41), .A2(_02090__PTR4), .ZN(_02112__PTR41) );
  AND2_X1 U11530 ( .A1(_02111__PTR42), .A2(_02090__PTR4), .ZN(_02112__PTR42) );
  AND2_X1 U11531 ( .A1(_02111__PTR43), .A2(_02090__PTR4), .ZN(_02112__PTR43) );
  AND2_X1 U11532 ( .A1(_02111__PTR44), .A2(_02090__PTR4), .ZN(_02112__PTR44) );
  AND2_X1 U11533 ( .A1(_02111__PTR45), .A2(_02090__PTR4), .ZN(_02112__PTR45) );
  AND2_X1 U11534 ( .A1(_02111__PTR46), .A2(_02090__PTR4), .ZN(_02112__PTR46) );
  AND2_X1 U11535 ( .A1(_02111__PTR47), .A2(_02090__PTR4), .ZN(_02112__PTR47) );
  AND2_X1 U11536 ( .A1(_02111__PTR16), .A2(_01863__PTR2), .ZN(_02112__PTR16) );
  AND2_X1 U11537 ( .A1(_02111__PTR17), .A2(_01863__PTR2), .ZN(_02112__PTR17) );
  AND2_X1 U11538 ( .A1(_02111__PTR18), .A2(_01863__PTR2), .ZN(_02112__PTR18) );
  AND2_X1 U11539 ( .A1(_02111__PTR19), .A2(_01863__PTR2), .ZN(_02112__PTR19) );
  AND2_X1 U11540 ( .A1(_02111__PTR20), .A2(_01863__PTR2), .ZN(_02112__PTR20) );
  AND2_X1 U11541 ( .A1(_02111__PTR21), .A2(_01863__PTR2), .ZN(_02112__PTR21) );
  AND2_X1 U11542 ( .A1(_02111__PTR22), .A2(_01863__PTR2), .ZN(_02112__PTR22) );
  AND2_X1 U11543 ( .A1(_02111__PTR23), .A2(_01863__PTR2), .ZN(_02112__PTR23) );
  AND2_X1 U11544 ( .A1(_02111__PTR24), .A2(_01863__PTR2), .ZN(_02112__PTR24) );
  AND2_X1 U11545 ( .A1(_02111__PTR25), .A2(_01863__PTR2), .ZN(_02112__PTR25) );
  AND2_X1 U11546 ( .A1(_02111__PTR26), .A2(_01863__PTR2), .ZN(_02112__PTR26) );
  AND2_X1 U11547 ( .A1(_02111__PTR27), .A2(_01863__PTR2), .ZN(_02112__PTR27) );
  AND2_X1 U11548 ( .A1(_02111__PTR28), .A2(_01863__PTR2), .ZN(_02112__PTR28) );
  AND2_X1 U11549 ( .A1(_02111__PTR29), .A2(_01863__PTR2), .ZN(_02112__PTR29) );
  AND2_X1 U11550 ( .A1(_02111__PTR30), .A2(_01863__PTR2), .ZN(_02112__PTR30) );
  AND2_X1 U11551 ( .A1(_02111__PTR31), .A2(_01863__PTR2), .ZN(_02112__PTR31) );
  AND2_X1 U11552 ( .A1(P1_P1_lWord_PTR0), .A2(_02109__PTR0), .ZN(_02112__PTR0) );
  AND2_X1 U11553 ( .A1(P1_P1_lWord_PTR1), .A2(_02109__PTR0), .ZN(_02112__PTR1) );
  AND2_X1 U11554 ( .A1(P1_P1_lWord_PTR2), .A2(_02109__PTR0), .ZN(_02112__PTR2) );
  AND2_X1 U11555 ( .A1(P1_P1_lWord_PTR3), .A2(_02109__PTR0), .ZN(_02112__PTR3) );
  AND2_X1 U11556 ( .A1(P1_P1_lWord_PTR4), .A2(_02109__PTR0), .ZN(_02112__PTR4) );
  AND2_X1 U11557 ( .A1(P1_P1_lWord_PTR5), .A2(_02109__PTR0), .ZN(_02112__PTR5) );
  AND2_X1 U11558 ( .A1(P1_P1_lWord_PTR6), .A2(_02109__PTR0), .ZN(_02112__PTR6) );
  AND2_X1 U11559 ( .A1(P1_P1_lWord_PTR7), .A2(_02109__PTR0), .ZN(_02112__PTR7) );
  AND2_X1 U11560 ( .A1(P1_P1_lWord_PTR8), .A2(_02109__PTR0), .ZN(_02112__PTR8) );
  AND2_X1 U11561 ( .A1(P1_P1_lWord_PTR9), .A2(_02109__PTR0), .ZN(_02112__PTR9) );
  AND2_X1 U11562 ( .A1(P1_P1_lWord_PTR10), .A2(_02109__PTR0), .ZN(_02112__PTR10) );
  AND2_X1 U11563 ( .A1(P1_P1_lWord_PTR11), .A2(_02109__PTR0), .ZN(_02112__PTR11) );
  AND2_X1 U11564 ( .A1(P1_P1_lWord_PTR12), .A2(_02109__PTR0), .ZN(_02112__PTR12) );
  AND2_X1 U11565 ( .A1(P1_P1_lWord_PTR13), .A2(_02109__PTR0), .ZN(_02112__PTR13) );
  AND2_X1 U11566 ( .A1(P1_P1_lWord_PTR14), .A2(_02109__PTR0), .ZN(_02112__PTR14) );
  AND2_X1 U11567 ( .A1(P1_P1_lWord_PTR15), .A2(_02109__PTR0), .ZN(_02112__PTR15) );
  AND2_X1 U11568 ( .A1(_02107__PTR30), .A2(_02090__PTR4), .ZN(_02108__PTR30) );
  AND2_X1 U11569 ( .A1(_02107__PTR31), .A2(_02090__PTR4), .ZN(_02108__PTR31) );
  AND2_X1 U11570 ( .A1(_02107__PTR32), .A2(_02090__PTR4), .ZN(_02108__PTR32) );
  AND2_X1 U11571 ( .A1(_02107__PTR33), .A2(_02090__PTR4), .ZN(_02108__PTR33) );
  AND2_X1 U11572 ( .A1(_02107__PTR34), .A2(_02090__PTR4), .ZN(_02108__PTR34) );
  AND2_X1 U11573 ( .A1(_02107__PTR35), .A2(_02090__PTR4), .ZN(_02108__PTR35) );
  AND2_X1 U11574 ( .A1(_02107__PTR36), .A2(_02090__PTR4), .ZN(_02108__PTR36) );
  AND2_X1 U11575 ( .A1(_02107__PTR37), .A2(_02090__PTR4), .ZN(_02108__PTR37) );
  AND2_X1 U11576 ( .A1(_02107__PTR38), .A2(_02090__PTR4), .ZN(_02108__PTR38) );
  AND2_X1 U11577 ( .A1(_02107__PTR39), .A2(_02090__PTR4), .ZN(_02108__PTR39) );
  AND2_X1 U11578 ( .A1(_02107__PTR40), .A2(_02090__PTR4), .ZN(_02108__PTR40) );
  AND2_X1 U11579 ( .A1(_02107__PTR41), .A2(_02090__PTR4), .ZN(_02108__PTR41) );
  AND2_X1 U11580 ( .A1(_02107__PTR42), .A2(_02090__PTR4), .ZN(_02108__PTR42) );
  AND2_X1 U11581 ( .A1(_02107__PTR43), .A2(_02090__PTR4), .ZN(_02108__PTR43) );
  AND2_X1 U11582 ( .A1(_02107__PTR44), .A2(_02090__PTR4), .ZN(_02108__PTR44) );
  AND2_X1 U11583 ( .A1(_02107__PTR15), .A2(_01863__PTR2), .ZN(_02108__PTR15) );
  AND2_X1 U11584 ( .A1(_02107__PTR16), .A2(_01863__PTR2), .ZN(_02108__PTR16) );
  AND2_X1 U11585 ( .A1(_02107__PTR17), .A2(_01863__PTR2), .ZN(_02108__PTR17) );
  AND2_X1 U11586 ( .A1(_02107__PTR18), .A2(_01863__PTR2), .ZN(_02108__PTR18) );
  AND2_X1 U11587 ( .A1(_02107__PTR19), .A2(_01863__PTR2), .ZN(_02108__PTR19) );
  AND2_X1 U11588 ( .A1(_02107__PTR20), .A2(_01863__PTR2), .ZN(_02108__PTR20) );
  AND2_X1 U11589 ( .A1(_02107__PTR21), .A2(_01863__PTR2), .ZN(_02108__PTR21) );
  AND2_X1 U11590 ( .A1(_02107__PTR22), .A2(_01863__PTR2), .ZN(_02108__PTR22) );
  AND2_X1 U11591 ( .A1(_02107__PTR23), .A2(_01863__PTR2), .ZN(_02108__PTR23) );
  AND2_X1 U11592 ( .A1(_02107__PTR24), .A2(_01863__PTR2), .ZN(_02108__PTR24) );
  AND2_X1 U11593 ( .A1(_02107__PTR25), .A2(_01863__PTR2), .ZN(_02108__PTR25) );
  AND2_X1 U11594 ( .A1(_02107__PTR26), .A2(_01863__PTR2), .ZN(_02108__PTR26) );
  AND2_X1 U11595 ( .A1(_02107__PTR27), .A2(_01863__PTR2), .ZN(_02108__PTR27) );
  AND2_X1 U11596 ( .A1(_02107__PTR28), .A2(_01863__PTR2), .ZN(_02108__PTR28) );
  AND2_X1 U11597 ( .A1(_02107__PTR29), .A2(_01863__PTR2), .ZN(_02108__PTR29) );
  AND2_X1 U11598 ( .A1(P1_P1_uWord_PTR0), .A2(_02109__PTR0), .ZN(_02108__PTR0) );
  AND2_X1 U11599 ( .A1(P1_P1_uWord_PTR1), .A2(_02109__PTR0), .ZN(_02108__PTR1) );
  AND2_X1 U11600 ( .A1(P1_P1_uWord_PTR2), .A2(_02109__PTR0), .ZN(_02108__PTR2) );
  AND2_X1 U11601 ( .A1(P1_P1_uWord_PTR3), .A2(_02109__PTR0), .ZN(_02108__PTR3) );
  AND2_X1 U11602 ( .A1(P1_P1_uWord_PTR4), .A2(_02109__PTR0), .ZN(_02108__PTR4) );
  AND2_X1 U11603 ( .A1(P1_P1_uWord_PTR5), .A2(_02109__PTR0), .ZN(_02108__PTR5) );
  AND2_X1 U11604 ( .A1(P1_P1_uWord_PTR6), .A2(_02109__PTR0), .ZN(_02108__PTR6) );
  AND2_X1 U11605 ( .A1(P1_P1_uWord_PTR7), .A2(_02109__PTR0), .ZN(_02108__PTR7) );
  AND2_X1 U11606 ( .A1(P1_P1_uWord_PTR8), .A2(_02109__PTR0), .ZN(_02108__PTR8) );
  AND2_X1 U11607 ( .A1(P1_P1_uWord_PTR9), .A2(_02109__PTR0), .ZN(_02108__PTR9) );
  AND2_X1 U11608 ( .A1(P1_P1_uWord_PTR10), .A2(_02109__PTR0), .ZN(_02108__PTR10) );
  AND2_X1 U11609 ( .A1(P1_P1_uWord_PTR11), .A2(_02109__PTR0), .ZN(_02108__PTR11) );
  AND2_X1 U11610 ( .A1(P1_P1_uWord_PTR12), .A2(_02109__PTR0), .ZN(_02108__PTR12) );
  AND2_X1 U11611 ( .A1(P1_P1_uWord_PTR13), .A2(_02109__PTR0), .ZN(_02108__PTR13) );
  AND2_X1 U11612 ( .A1(P1_P1_uWord_PTR14), .A2(_02109__PTR0), .ZN(_02108__PTR14) );
  AND2_X1 U11613 ( .A1(P1_EBX_PTR0), .A2(_02102__PTR0), .ZN(_02101__PTR0) );
  AND2_X1 U11614 ( .A1(P1_EBX_PTR1), .A2(_02102__PTR0), .ZN(_02101__PTR1) );
  AND2_X1 U11615 ( .A1(P1_EBX_PTR2), .A2(_02102__PTR0), .ZN(_02101__PTR2) );
  AND2_X1 U11616 ( .A1(P1_EBX_PTR3), .A2(_02102__PTR0), .ZN(_02101__PTR3) );
  AND2_X1 U11617 ( .A1(P1_EBX_PTR4), .A2(_02102__PTR0), .ZN(_02101__PTR4) );
  AND2_X1 U11618 ( .A1(P1_EBX_PTR5), .A2(_02102__PTR0), .ZN(_02101__PTR5) );
  AND2_X1 U11619 ( .A1(P1_EBX_PTR6), .A2(_02102__PTR0), .ZN(_02101__PTR6) );
  AND2_X1 U11620 ( .A1(P1_EBX_PTR7), .A2(_02102__PTR0), .ZN(_02101__PTR7) );
  AND2_X1 U11621 ( .A1(P1_EBX_PTR8), .A2(_02102__PTR0), .ZN(_02101__PTR8) );
  AND2_X1 U11622 ( .A1(P1_EBX_PTR9), .A2(_02102__PTR0), .ZN(_02101__PTR9) );
  AND2_X1 U11623 ( .A1(P1_EBX_PTR10), .A2(_02102__PTR0), .ZN(_02101__PTR10) );
  AND2_X1 U11624 ( .A1(P1_EBX_PTR11), .A2(_02102__PTR0), .ZN(_02101__PTR11) );
  AND2_X1 U11625 ( .A1(P1_EBX_PTR12), .A2(_02102__PTR0), .ZN(_02101__PTR12) );
  AND2_X1 U11626 ( .A1(P1_EBX_PTR13), .A2(_02102__PTR0), .ZN(_02101__PTR13) );
  AND2_X1 U11627 ( .A1(P1_EBX_PTR14), .A2(_02102__PTR0), .ZN(_02101__PTR14) );
  AND2_X1 U11628 ( .A1(P1_EBX_PTR15), .A2(_02102__PTR0), .ZN(_02101__PTR15) );
  AND2_X1 U11629 ( .A1(P1_EBX_PTR16), .A2(_02102__PTR0), .ZN(_02101__PTR16) );
  AND2_X1 U11630 ( .A1(P1_EBX_PTR17), .A2(_02102__PTR0), .ZN(_02101__PTR17) );
  AND2_X1 U11631 ( .A1(P1_EBX_PTR18), .A2(_02102__PTR0), .ZN(_02101__PTR18) );
  AND2_X1 U11632 ( .A1(P1_EBX_PTR19), .A2(_02102__PTR0), .ZN(_02101__PTR19) );
  AND2_X1 U11633 ( .A1(P1_EBX_PTR20), .A2(_02102__PTR0), .ZN(_02101__PTR20) );
  AND2_X1 U11634 ( .A1(P1_EBX_PTR21), .A2(_02102__PTR0), .ZN(_02101__PTR21) );
  AND2_X1 U11635 ( .A1(P1_EBX_PTR22), .A2(_02102__PTR0), .ZN(_02101__PTR22) );
  AND2_X1 U11636 ( .A1(P1_EBX_PTR23), .A2(_02102__PTR0), .ZN(_02101__PTR23) );
  AND2_X1 U11637 ( .A1(P1_EBX_PTR24), .A2(_02102__PTR0), .ZN(_02101__PTR24) );
  AND2_X1 U11638 ( .A1(P1_EBX_PTR25), .A2(_02102__PTR0), .ZN(_02101__PTR25) );
  AND2_X1 U11639 ( .A1(P1_EBX_PTR26), .A2(_02102__PTR0), .ZN(_02101__PTR26) );
  AND2_X1 U11640 ( .A1(P1_EBX_PTR27), .A2(_02102__PTR0), .ZN(_02101__PTR27) );
  AND2_X1 U11641 ( .A1(P1_EBX_PTR28), .A2(_02102__PTR0), .ZN(_02101__PTR28) );
  AND2_X1 U11642 ( .A1(P1_EBX_PTR29), .A2(_02102__PTR0), .ZN(_02101__PTR29) );
  AND2_X1 U11643 ( .A1(P1_EBX_PTR30), .A2(_02102__PTR0), .ZN(_02101__PTR30) );
  AND2_X1 U11644 ( .A1(P1_EBX_PTR31), .A2(_02102__PTR0), .ZN(_02101__PTR31) );
  AND2_X1 U11645 ( .A1(_02100__PTR32), .A2(_02102__PTR1), .ZN(_02101__PTR32) );
  AND2_X1 U11646 ( .A1(_02100__PTR33), .A2(_02102__PTR1), .ZN(_02101__PTR33) );
  AND2_X1 U11647 ( .A1(_02100__PTR34), .A2(_02102__PTR1), .ZN(_02101__PTR34) );
  AND2_X1 U11648 ( .A1(_02100__PTR35), .A2(_02102__PTR1), .ZN(_02101__PTR35) );
  AND2_X1 U11649 ( .A1(_02100__PTR36), .A2(_02102__PTR1), .ZN(_02101__PTR36) );
  AND2_X1 U11650 ( .A1(_02100__PTR37), .A2(_02102__PTR1), .ZN(_02101__PTR37) );
  AND2_X1 U11651 ( .A1(_02100__PTR38), .A2(_02102__PTR1), .ZN(_02101__PTR38) );
  AND2_X1 U11652 ( .A1(_02100__PTR39), .A2(_02102__PTR1), .ZN(_02101__PTR39) );
  AND2_X1 U11653 ( .A1(_02100__PTR40), .A2(_02102__PTR1), .ZN(_02101__PTR40) );
  AND2_X1 U11654 ( .A1(_02100__PTR41), .A2(_02102__PTR1), .ZN(_02101__PTR41) );
  AND2_X1 U11655 ( .A1(_02100__PTR42), .A2(_02102__PTR1), .ZN(_02101__PTR42) );
  AND2_X1 U11656 ( .A1(_02100__PTR43), .A2(_02102__PTR1), .ZN(_02101__PTR43) );
  AND2_X1 U11657 ( .A1(_02100__PTR44), .A2(_02102__PTR1), .ZN(_02101__PTR44) );
  AND2_X1 U11658 ( .A1(_02100__PTR45), .A2(_02102__PTR1), .ZN(_02101__PTR45) );
  AND2_X1 U11659 ( .A1(_02100__PTR46), .A2(_02102__PTR1), .ZN(_02101__PTR46) );
  AND2_X1 U11660 ( .A1(_02100__PTR47), .A2(_02102__PTR1), .ZN(_02101__PTR47) );
  AND2_X1 U11661 ( .A1(_02100__PTR48), .A2(_02102__PTR1), .ZN(_02101__PTR48) );
  AND2_X1 U11662 ( .A1(_02100__PTR49), .A2(_02102__PTR1), .ZN(_02101__PTR49) );
  AND2_X1 U11663 ( .A1(_02100__PTR50), .A2(_02102__PTR1), .ZN(_02101__PTR50) );
  AND2_X1 U11664 ( .A1(_02100__PTR51), .A2(_02102__PTR1), .ZN(_02101__PTR51) );
  AND2_X1 U11665 ( .A1(_02100__PTR52), .A2(_02102__PTR1), .ZN(_02101__PTR52) );
  AND2_X1 U11666 ( .A1(_02100__PTR53), .A2(_02102__PTR1), .ZN(_02101__PTR53) );
  AND2_X1 U11667 ( .A1(_02100__PTR54), .A2(_02102__PTR1), .ZN(_02101__PTR54) );
  AND2_X1 U11668 ( .A1(_02100__PTR55), .A2(_02102__PTR1), .ZN(_02101__PTR55) );
  AND2_X1 U11669 ( .A1(_02100__PTR56), .A2(_02102__PTR1), .ZN(_02101__PTR56) );
  AND2_X1 U11670 ( .A1(_02100__PTR57), .A2(_02102__PTR1), .ZN(_02101__PTR57) );
  AND2_X1 U11671 ( .A1(_02100__PTR58), .A2(_02102__PTR1), .ZN(_02101__PTR58) );
  AND2_X1 U11672 ( .A1(_02100__PTR59), .A2(_02102__PTR1), .ZN(_02101__PTR59) );
  AND2_X1 U11673 ( .A1(_02100__PTR60), .A2(_02102__PTR1), .ZN(_02101__PTR60) );
  AND2_X1 U11674 ( .A1(_02100__PTR61), .A2(_02102__PTR1), .ZN(_02101__PTR61) );
  AND2_X1 U11675 ( .A1(_02100__PTR62), .A2(_02102__PTR1), .ZN(_02101__PTR62) );
  AND2_X1 U11676 ( .A1(_02100__PTR63), .A2(_02102__PTR1), .ZN(_02101__PTR63) );
  AND2_X1 U11677 ( .A1(_02100__PTR64), .A2(_02102__PTR2), .ZN(_02101__PTR64) );
  AND2_X1 U11678 ( .A1(_02100__PTR65), .A2(_02102__PTR2), .ZN(_02101__PTR65) );
  AND2_X1 U11679 ( .A1(_02100__PTR66), .A2(_02102__PTR2), .ZN(_02101__PTR66) );
  AND2_X1 U11680 ( .A1(_02100__PTR67), .A2(_02102__PTR2), .ZN(_02101__PTR67) );
  AND2_X1 U11681 ( .A1(_02100__PTR68), .A2(_02102__PTR2), .ZN(_02101__PTR68) );
  AND2_X1 U11682 ( .A1(_02100__PTR69), .A2(_02102__PTR2), .ZN(_02101__PTR69) );
  AND2_X1 U11683 ( .A1(_02100__PTR70), .A2(_02102__PTR2), .ZN(_02101__PTR70) );
  AND2_X1 U11684 ( .A1(_02100__PTR71), .A2(_02102__PTR2), .ZN(_02101__PTR71) );
  AND2_X1 U11685 ( .A1(_02100__PTR72), .A2(_02102__PTR2), .ZN(_02101__PTR72) );
  AND2_X1 U11686 ( .A1(_02100__PTR73), .A2(_02102__PTR2), .ZN(_02101__PTR73) );
  AND2_X1 U11687 ( .A1(_02100__PTR74), .A2(_02102__PTR2), .ZN(_02101__PTR74) );
  AND2_X1 U11688 ( .A1(_02100__PTR75), .A2(_02102__PTR2), .ZN(_02101__PTR75) );
  AND2_X1 U11689 ( .A1(_02100__PTR76), .A2(_02102__PTR2), .ZN(_02101__PTR76) );
  AND2_X1 U11690 ( .A1(_02100__PTR77), .A2(_02102__PTR2), .ZN(_02101__PTR77) );
  AND2_X1 U11691 ( .A1(_02100__PTR78), .A2(_02102__PTR2), .ZN(_02101__PTR78) );
  AND2_X1 U11692 ( .A1(_02100__PTR79), .A2(_02102__PTR2), .ZN(_02101__PTR79) );
  AND2_X1 U11693 ( .A1(_02100__PTR80), .A2(_02102__PTR2), .ZN(_02101__PTR80) );
  AND2_X1 U11694 ( .A1(_02100__PTR81), .A2(_02102__PTR2), .ZN(_02101__PTR81) );
  AND2_X1 U11695 ( .A1(_02100__PTR82), .A2(_02102__PTR2), .ZN(_02101__PTR82) );
  AND2_X1 U11696 ( .A1(_02100__PTR83), .A2(_02102__PTR2), .ZN(_02101__PTR83) );
  AND2_X1 U11697 ( .A1(_02100__PTR84), .A2(_02102__PTR2), .ZN(_02101__PTR84) );
  AND2_X1 U11698 ( .A1(_02100__PTR85), .A2(_02102__PTR2), .ZN(_02101__PTR85) );
  AND2_X1 U11699 ( .A1(_02100__PTR86), .A2(_02102__PTR2), .ZN(_02101__PTR86) );
  AND2_X1 U11700 ( .A1(_02100__PTR87), .A2(_02102__PTR2), .ZN(_02101__PTR87) );
  AND2_X1 U11701 ( .A1(_02100__PTR88), .A2(_02102__PTR2), .ZN(_02101__PTR88) );
  AND2_X1 U11702 ( .A1(_02100__PTR89), .A2(_02102__PTR2), .ZN(_02101__PTR89) );
  AND2_X1 U11703 ( .A1(_02100__PTR90), .A2(_02102__PTR2), .ZN(_02101__PTR90) );
  AND2_X1 U11704 ( .A1(_02100__PTR91), .A2(_02102__PTR2), .ZN(_02101__PTR91) );
  AND2_X1 U11705 ( .A1(_02100__PTR92), .A2(_02102__PTR2), .ZN(_02101__PTR92) );
  AND2_X1 U11706 ( .A1(_02100__PTR93), .A2(_02102__PTR2), .ZN(_02101__PTR93) );
  AND2_X1 U11707 ( .A1(_02100__PTR94), .A2(_02102__PTR2), .ZN(_02101__PTR94) );
  AND2_X1 U11708 ( .A1(_02100__PTR95), .A2(_02102__PTR2), .ZN(_02101__PTR95) );
  AND2_X1 U11709 ( .A1(_02096__PTR128), .A2(_02098__PTR4), .ZN(_02097__PTR128) );
  AND2_X1 U11710 ( .A1(_02096__PTR129), .A2(_02098__PTR4), .ZN(_02097__PTR129) );
  AND2_X1 U11711 ( .A1(_02096__PTR130), .A2(_02098__PTR4), .ZN(_02097__PTR130) );
  AND2_X1 U11712 ( .A1(_02096__PTR131), .A2(_02098__PTR4), .ZN(_02097__PTR131) );
  AND2_X1 U11713 ( .A1(_02096__PTR132), .A2(_02098__PTR4), .ZN(_02097__PTR132) );
  AND2_X1 U11714 ( .A1(_02096__PTR133), .A2(_02098__PTR4), .ZN(_02097__PTR133) );
  AND2_X1 U11715 ( .A1(_02096__PTR134), .A2(_02098__PTR4), .ZN(_02097__PTR134) );
  AND2_X1 U11716 ( .A1(_02096__PTR135), .A2(_02098__PTR4), .ZN(_02097__PTR135) );
  AND2_X1 U11717 ( .A1(_02096__PTR136), .A2(_02098__PTR4), .ZN(_02097__PTR136) );
  AND2_X1 U11718 ( .A1(_02096__PTR137), .A2(_02098__PTR4), .ZN(_02097__PTR137) );
  AND2_X1 U11719 ( .A1(_02096__PTR138), .A2(_02098__PTR4), .ZN(_02097__PTR138) );
  AND2_X1 U11720 ( .A1(_02096__PTR139), .A2(_02098__PTR4), .ZN(_02097__PTR139) );
  AND2_X1 U11721 ( .A1(_02096__PTR140), .A2(_02098__PTR4), .ZN(_02097__PTR140) );
  AND2_X1 U11722 ( .A1(_02096__PTR141), .A2(_02098__PTR4), .ZN(_02097__PTR141) );
  AND2_X1 U11723 ( .A1(_02096__PTR142), .A2(_02098__PTR4), .ZN(_02097__PTR142) );
  AND2_X1 U11724 ( .A1(_02096__PTR143), .A2(_02098__PTR4), .ZN(_02097__PTR143) );
  AND2_X1 U11725 ( .A1(_02096__PTR144), .A2(_02098__PTR4), .ZN(_02097__PTR144) );
  AND2_X1 U11726 ( .A1(_02096__PTR145), .A2(_02098__PTR4), .ZN(_02097__PTR145) );
  AND2_X1 U11727 ( .A1(_02096__PTR146), .A2(_02098__PTR4), .ZN(_02097__PTR146) );
  AND2_X1 U11728 ( .A1(_02096__PTR147), .A2(_02098__PTR4), .ZN(_02097__PTR147) );
  AND2_X1 U11729 ( .A1(_02096__PTR148), .A2(_02098__PTR4), .ZN(_02097__PTR148) );
  AND2_X1 U11730 ( .A1(_02096__PTR149), .A2(_02098__PTR4), .ZN(_02097__PTR149) );
  AND2_X1 U11731 ( .A1(_02096__PTR150), .A2(_02098__PTR4), .ZN(_02097__PTR150) );
  AND2_X1 U11732 ( .A1(_02096__PTR151), .A2(_02098__PTR4), .ZN(_02097__PTR151) );
  AND2_X1 U11733 ( .A1(_02096__PTR152), .A2(_02098__PTR4), .ZN(_02097__PTR152) );
  AND2_X1 U11734 ( .A1(_02096__PTR153), .A2(_02098__PTR4), .ZN(_02097__PTR153) );
  AND2_X1 U11735 ( .A1(_02096__PTR154), .A2(_02098__PTR4), .ZN(_02097__PTR154) );
  AND2_X1 U11736 ( .A1(_02096__PTR155), .A2(_02098__PTR4), .ZN(_02097__PTR155) );
  AND2_X1 U11737 ( .A1(_02096__PTR156), .A2(_02098__PTR4), .ZN(_02097__PTR156) );
  AND2_X1 U11738 ( .A1(_02096__PTR157), .A2(_02098__PTR4), .ZN(_02097__PTR157) );
  AND2_X1 U11739 ( .A1(_02096__PTR158), .A2(_02098__PTR4), .ZN(_02097__PTR158) );
  AND2_X1 U11740 ( .A1(_02096__PTR159), .A2(_02098__PTR4), .ZN(_02097__PTR159) );
  AND2_X1 U11741 ( .A1(_02096__PTR96), .A2(_02090__PTR4), .ZN(_02097__PTR96) );
  AND2_X1 U11742 ( .A1(_02096__PTR97), .A2(_02090__PTR4), .ZN(_02097__PTR97) );
  AND2_X1 U11743 ( .A1(_02096__PTR98), .A2(_02090__PTR4), .ZN(_02097__PTR98) );
  AND2_X1 U11744 ( .A1(_02096__PTR99), .A2(_02090__PTR4), .ZN(_02097__PTR99) );
  AND2_X1 U11745 ( .A1(_02096__PTR100), .A2(_02090__PTR4), .ZN(_02097__PTR100) );
  AND2_X1 U11746 ( .A1(_02096__PTR101), .A2(_02090__PTR4), .ZN(_02097__PTR101) );
  AND2_X1 U11747 ( .A1(_02096__PTR102), .A2(_02090__PTR4), .ZN(_02097__PTR102) );
  AND2_X1 U11748 ( .A1(_02096__PTR103), .A2(_02090__PTR4), .ZN(_02097__PTR103) );
  AND2_X1 U11749 ( .A1(_02096__PTR104), .A2(_02090__PTR4), .ZN(_02097__PTR104) );
  AND2_X1 U11750 ( .A1(_02096__PTR105), .A2(_02090__PTR4), .ZN(_02097__PTR105) );
  AND2_X1 U11751 ( .A1(_02096__PTR106), .A2(_02090__PTR4), .ZN(_02097__PTR106) );
  AND2_X1 U11752 ( .A1(_02096__PTR107), .A2(_02090__PTR4), .ZN(_02097__PTR107) );
  AND2_X1 U11753 ( .A1(_02096__PTR108), .A2(_02090__PTR4), .ZN(_02097__PTR108) );
  AND2_X1 U11754 ( .A1(_02096__PTR109), .A2(_02090__PTR4), .ZN(_02097__PTR109) );
  AND2_X1 U11755 ( .A1(_02096__PTR110), .A2(_02090__PTR4), .ZN(_02097__PTR110) );
  AND2_X1 U11756 ( .A1(_02096__PTR111), .A2(_02090__PTR4), .ZN(_02097__PTR111) );
  AND2_X1 U11757 ( .A1(_02096__PTR112), .A2(_02090__PTR4), .ZN(_02097__PTR112) );
  AND2_X1 U11758 ( .A1(_02096__PTR113), .A2(_02090__PTR4), .ZN(_02097__PTR113) );
  AND2_X1 U11759 ( .A1(_02096__PTR114), .A2(_02090__PTR4), .ZN(_02097__PTR114) );
  AND2_X1 U11760 ( .A1(_02096__PTR115), .A2(_02090__PTR4), .ZN(_02097__PTR115) );
  AND2_X1 U11761 ( .A1(_02096__PTR116), .A2(_02090__PTR4), .ZN(_02097__PTR116) );
  AND2_X1 U11762 ( .A1(_02096__PTR117), .A2(_02090__PTR4), .ZN(_02097__PTR117) );
  AND2_X1 U11763 ( .A1(_02096__PTR118), .A2(_02090__PTR4), .ZN(_02097__PTR118) );
  AND2_X1 U11764 ( .A1(_02096__PTR119), .A2(_02090__PTR4), .ZN(_02097__PTR119) );
  AND2_X1 U11765 ( .A1(_02096__PTR120), .A2(_02090__PTR4), .ZN(_02097__PTR120) );
  AND2_X1 U11766 ( .A1(_02096__PTR121), .A2(_02090__PTR4), .ZN(_02097__PTR121) );
  AND2_X1 U11767 ( .A1(_02096__PTR122), .A2(_02090__PTR4), .ZN(_02097__PTR122) );
  AND2_X1 U11768 ( .A1(_02096__PTR123), .A2(_02090__PTR4), .ZN(_02097__PTR123) );
  AND2_X1 U11769 ( .A1(_02096__PTR124), .A2(_02090__PTR4), .ZN(_02097__PTR124) );
  AND2_X1 U11770 ( .A1(_02096__PTR125), .A2(_02090__PTR4), .ZN(_02097__PTR125) );
  AND2_X1 U11771 ( .A1(_02096__PTR126), .A2(_02090__PTR4), .ZN(_02097__PTR126) );
  AND2_X1 U11772 ( .A1(_02096__PTR127), .A2(_02090__PTR4), .ZN(_02097__PTR127) );
  AND2_X1 U11773 ( .A1(_02096__PTR96), .A2(_02090__PTR3), .ZN(_02097__PTR64) );
  AND2_X1 U11774 ( .A1(_02096__PTR97), .A2(_02090__PTR3), .ZN(_02097__PTR65) );
  AND2_X1 U11775 ( .A1(_02096__PTR98), .A2(_02090__PTR3), .ZN(_02097__PTR66) );
  AND2_X1 U11776 ( .A1(_02096__PTR99), .A2(_02090__PTR3), .ZN(_02097__PTR67) );
  AND2_X1 U11777 ( .A1(_02096__PTR100), .A2(_02090__PTR3), .ZN(_02097__PTR68) );
  AND2_X1 U11778 ( .A1(_02096__PTR101), .A2(_02090__PTR3), .ZN(_02097__PTR69) );
  AND2_X1 U11779 ( .A1(_02096__PTR102), .A2(_02090__PTR3), .ZN(_02097__PTR70) );
  AND2_X1 U11780 ( .A1(_02096__PTR103), .A2(_02090__PTR3), .ZN(_02097__PTR71) );
  AND2_X1 U11781 ( .A1(_02096__PTR104), .A2(_02090__PTR3), .ZN(_02097__PTR72) );
  AND2_X1 U11782 ( .A1(_02096__PTR105), .A2(_02090__PTR3), .ZN(_02097__PTR73) );
  AND2_X1 U11783 ( .A1(_02096__PTR106), .A2(_02090__PTR3), .ZN(_02097__PTR74) );
  AND2_X1 U11784 ( .A1(_02096__PTR107), .A2(_02090__PTR3), .ZN(_02097__PTR75) );
  AND2_X1 U11785 ( .A1(_02096__PTR108), .A2(_02090__PTR3), .ZN(_02097__PTR76) );
  AND2_X1 U11786 ( .A1(_02096__PTR109), .A2(_02090__PTR3), .ZN(_02097__PTR77) );
  AND2_X1 U11787 ( .A1(_02096__PTR110), .A2(_02090__PTR3), .ZN(_02097__PTR78) );
  AND2_X1 U11788 ( .A1(_02096__PTR111), .A2(_02090__PTR3), .ZN(_02097__PTR79) );
  AND2_X1 U11789 ( .A1(_02096__PTR80), .A2(_02090__PTR3), .ZN(_02097__PTR80) );
  AND2_X1 U11790 ( .A1(_02096__PTR81), .A2(_02090__PTR3), .ZN(_02097__PTR81) );
  AND2_X1 U11791 ( .A1(_02096__PTR82), .A2(_02090__PTR3), .ZN(_02097__PTR82) );
  AND2_X1 U11792 ( .A1(_02096__PTR83), .A2(_02090__PTR3), .ZN(_02097__PTR83) );
  AND2_X1 U11793 ( .A1(_02096__PTR84), .A2(_02090__PTR3), .ZN(_02097__PTR84) );
  AND2_X1 U11794 ( .A1(_02096__PTR85), .A2(_02090__PTR3), .ZN(_02097__PTR85) );
  AND2_X1 U11795 ( .A1(_02096__PTR86), .A2(_02090__PTR3), .ZN(_02097__PTR86) );
  AND2_X1 U11796 ( .A1(_02096__PTR87), .A2(_02090__PTR3), .ZN(_02097__PTR87) );
  AND2_X1 U11797 ( .A1(_02096__PTR88), .A2(_02090__PTR3), .ZN(_02097__PTR88) );
  AND2_X1 U11798 ( .A1(_02096__PTR89), .A2(_02090__PTR3), .ZN(_02097__PTR89) );
  AND2_X1 U11799 ( .A1(_02096__PTR90), .A2(_02090__PTR3), .ZN(_02097__PTR90) );
  AND2_X1 U11800 ( .A1(_02096__PTR91), .A2(_02090__PTR3), .ZN(_02097__PTR91) );
  AND2_X1 U11801 ( .A1(_02096__PTR92), .A2(_02090__PTR3), .ZN(_02097__PTR92) );
  AND2_X1 U11802 ( .A1(_02096__PTR93), .A2(_02090__PTR3), .ZN(_02097__PTR93) );
  AND2_X1 U11803 ( .A1(_02096__PTR94), .A2(_02090__PTR3), .ZN(_02097__PTR94) );
  AND2_X1 U11804 ( .A1(_02096__PTR95), .A2(_02090__PTR3), .ZN(_02097__PTR95) );
  AND2_X1 U11805 ( .A1(_02096__PTR32), .A2(_02098__PTR1), .ZN(_02097__PTR32) );
  AND2_X1 U11806 ( .A1(_02096__PTR33), .A2(_02098__PTR1), .ZN(_02097__PTR33) );
  AND2_X1 U11807 ( .A1(_02096__PTR34), .A2(_02098__PTR1), .ZN(_02097__PTR34) );
  AND2_X1 U11808 ( .A1(_02096__PTR35), .A2(_02098__PTR1), .ZN(_02097__PTR35) );
  AND2_X1 U11809 ( .A1(_02096__PTR36), .A2(_02098__PTR1), .ZN(_02097__PTR36) );
  AND2_X1 U11810 ( .A1(_02096__PTR37), .A2(_02098__PTR1), .ZN(_02097__PTR37) );
  AND2_X1 U11811 ( .A1(_02096__PTR38), .A2(_02098__PTR1), .ZN(_02097__PTR38) );
  AND2_X1 U11812 ( .A1(_02096__PTR39), .A2(_02098__PTR1), .ZN(_02097__PTR39) );
  AND2_X1 U11813 ( .A1(_02096__PTR40), .A2(_02098__PTR1), .ZN(_02097__PTR40) );
  AND2_X1 U11814 ( .A1(_02096__PTR41), .A2(_02098__PTR1), .ZN(_02097__PTR41) );
  AND2_X1 U11815 ( .A1(_02096__PTR42), .A2(_02098__PTR1), .ZN(_02097__PTR42) );
  AND2_X1 U11816 ( .A1(_02096__PTR43), .A2(_02098__PTR1), .ZN(_02097__PTR43) );
  AND2_X1 U11817 ( .A1(_02096__PTR44), .A2(_02098__PTR1), .ZN(_02097__PTR44) );
  AND2_X1 U11818 ( .A1(_02096__PTR45), .A2(_02098__PTR1), .ZN(_02097__PTR45) );
  AND2_X1 U11819 ( .A1(_02096__PTR46), .A2(_02098__PTR1), .ZN(_02097__PTR46) );
  AND2_X1 U11820 ( .A1(_02096__PTR47), .A2(_02098__PTR1), .ZN(_02097__PTR47) );
  AND2_X1 U11821 ( .A1(_02096__PTR48), .A2(_02098__PTR1), .ZN(_02097__PTR48) );
  AND2_X1 U11822 ( .A1(_02096__PTR49), .A2(_02098__PTR1), .ZN(_02097__PTR49) );
  AND2_X1 U11823 ( .A1(_02096__PTR50), .A2(_02098__PTR1), .ZN(_02097__PTR50) );
  AND2_X1 U11824 ( .A1(_02096__PTR51), .A2(_02098__PTR1), .ZN(_02097__PTR51) );
  AND2_X1 U11825 ( .A1(_02096__PTR52), .A2(_02098__PTR1), .ZN(_02097__PTR52) );
  AND2_X1 U11826 ( .A1(_02096__PTR53), .A2(_02098__PTR1), .ZN(_02097__PTR53) );
  AND2_X1 U11827 ( .A1(_02096__PTR54), .A2(_02098__PTR1), .ZN(_02097__PTR54) );
  AND2_X1 U11828 ( .A1(_02096__PTR55), .A2(_02098__PTR1), .ZN(_02097__PTR55) );
  AND2_X1 U11829 ( .A1(_02096__PTR56), .A2(_02098__PTR1), .ZN(_02097__PTR56) );
  AND2_X1 U11830 ( .A1(_02096__PTR57), .A2(_02098__PTR1), .ZN(_02097__PTR57) );
  AND2_X1 U11831 ( .A1(_02096__PTR58), .A2(_02098__PTR1), .ZN(_02097__PTR58) );
  AND2_X1 U11832 ( .A1(_02096__PTR59), .A2(_02098__PTR1), .ZN(_02097__PTR59) );
  AND2_X1 U11833 ( .A1(_02096__PTR60), .A2(_02098__PTR1), .ZN(_02097__PTR60) );
  AND2_X1 U11834 ( .A1(_02096__PTR61), .A2(_02098__PTR1), .ZN(_02097__PTR61) );
  AND2_X1 U11835 ( .A1(_02096__PTR62), .A2(_02098__PTR1), .ZN(_02097__PTR62) );
  AND2_X1 U11836 ( .A1(_02096__PTR63), .A2(_02098__PTR1), .ZN(_02097__PTR63) );
  AND2_X1 U11837 ( .A1(P1_EAX_PTR0), .A2(_02098__PTR0), .ZN(_02097__PTR0) );
  AND2_X1 U11838 ( .A1(P1_EAX_PTR1), .A2(_02098__PTR0), .ZN(_02097__PTR1) );
  AND2_X1 U11839 ( .A1(P1_EAX_PTR2), .A2(_02098__PTR0), .ZN(_02097__PTR2) );
  AND2_X1 U11840 ( .A1(P1_EAX_PTR3), .A2(_02098__PTR0), .ZN(_02097__PTR3) );
  AND2_X1 U11841 ( .A1(P1_EAX_PTR4), .A2(_02098__PTR0), .ZN(_02097__PTR4) );
  AND2_X1 U11842 ( .A1(P1_EAX_PTR5), .A2(_02098__PTR0), .ZN(_02097__PTR5) );
  AND2_X1 U11843 ( .A1(P1_EAX_PTR6), .A2(_02098__PTR0), .ZN(_02097__PTR6) );
  AND2_X1 U11844 ( .A1(P1_EAX_PTR7), .A2(_02098__PTR0), .ZN(_02097__PTR7) );
  AND2_X1 U11845 ( .A1(P1_EAX_PTR8), .A2(_02098__PTR0), .ZN(_02097__PTR8) );
  AND2_X1 U11846 ( .A1(P1_EAX_PTR9), .A2(_02098__PTR0), .ZN(_02097__PTR9) );
  AND2_X1 U11847 ( .A1(P1_EAX_PTR10), .A2(_02098__PTR0), .ZN(_02097__PTR10) );
  AND2_X1 U11848 ( .A1(P1_EAX_PTR11), .A2(_02098__PTR0), .ZN(_02097__PTR11) );
  AND2_X1 U11849 ( .A1(P1_EAX_PTR12), .A2(_02098__PTR0), .ZN(_02097__PTR12) );
  AND2_X1 U11850 ( .A1(P1_EAX_PTR13), .A2(_02098__PTR0), .ZN(_02097__PTR13) );
  AND2_X1 U11851 ( .A1(P1_EAX_PTR14), .A2(_02098__PTR0), .ZN(_02097__PTR14) );
  AND2_X1 U11852 ( .A1(P1_EAX_PTR15), .A2(_02098__PTR0), .ZN(_02097__PTR15) );
  AND2_X1 U11853 ( .A1(P1_EAX_PTR16), .A2(_02098__PTR0), .ZN(_02097__PTR16) );
  AND2_X1 U11854 ( .A1(P1_EAX_PTR17), .A2(_02098__PTR0), .ZN(_02097__PTR17) );
  AND2_X1 U11855 ( .A1(P1_EAX_PTR18), .A2(_02098__PTR0), .ZN(_02097__PTR18) );
  AND2_X1 U11856 ( .A1(P1_EAX_PTR19), .A2(_02098__PTR0), .ZN(_02097__PTR19) );
  AND2_X1 U11857 ( .A1(P1_EAX_PTR20), .A2(_02098__PTR0), .ZN(_02097__PTR20) );
  AND2_X1 U11858 ( .A1(P1_EAX_PTR21), .A2(_02098__PTR0), .ZN(_02097__PTR21) );
  AND2_X1 U11859 ( .A1(P1_EAX_PTR22), .A2(_02098__PTR0), .ZN(_02097__PTR22) );
  AND2_X1 U11860 ( .A1(P1_EAX_PTR23), .A2(_02098__PTR0), .ZN(_02097__PTR23) );
  AND2_X1 U11861 ( .A1(P1_EAX_PTR24), .A2(_02098__PTR0), .ZN(_02097__PTR24) );
  AND2_X1 U11862 ( .A1(P1_EAX_PTR25), .A2(_02098__PTR0), .ZN(_02097__PTR25) );
  AND2_X1 U11863 ( .A1(P1_EAX_PTR26), .A2(_02098__PTR0), .ZN(_02097__PTR26) );
  AND2_X1 U11864 ( .A1(P1_EAX_PTR27), .A2(_02098__PTR0), .ZN(_02097__PTR27) );
  AND2_X1 U11865 ( .A1(P1_EAX_PTR28), .A2(_02098__PTR0), .ZN(_02097__PTR28) );
  AND2_X1 U11866 ( .A1(P1_EAX_PTR29), .A2(_02098__PTR0), .ZN(_02097__PTR29) );
  AND2_X1 U11867 ( .A1(P1_EAX_PTR30), .A2(_02098__PTR0), .ZN(_02097__PTR30) );
  AND2_X1 U11868 ( .A1(P1_EAX_PTR31), .A2(_02098__PTR0), .ZN(_02097__PTR31) );
  AND2_X1 U11869 ( .A1(_01857__PTR3), .A2(_01855__PTR3), .ZN(_01858__PTR3) );
  AND2_X1 U11870 ( .A1(_01857__PTR2), .A2(_01859__PTR2), .ZN(_01858__PTR2) );
  AND2_X1 U11871 ( .A1(_01857__PTR1), .A2(_01855__PTR1), .ZN(_01858__PTR1) );
  AND2_X1 U11872 ( .A1(_01857__PTR0), .A2(_01855__PTR0), .ZN(_01858__PTR0) );
  AND2_X1 U11873 ( .A1(_01853__PTR0), .A2(_01855__PTR0), .ZN(_01854__PTR0) );
  AND2_X1 U11874 ( .A1(_01853__PTR1), .A2(_01855__PTR1), .ZN(_01854__PTR1) );
  AND2_X1 U11875 ( .A1(_01853__PTR2), .A2(_01855__PTR2), .ZN(_01854__PTR2) );
  AND2_X1 U11876 ( .A1(_01853__PTR3), .A2(_01855__PTR3), .ZN(_01854__PTR3) );
  AND2_X1 U11877 ( .A1(P1_P1_InstQueueRd_Addr_PTR0), .A2(_02090__PTR6), .ZN(_02089__PTR30) );
  AND2_X1 U11878 ( .A1(P1_P1_InstQueueRd_Addr_PTR1), .A2(_02090__PTR6), .ZN(_02089__PTR31) );
  AND2_X1 U11879 ( .A1(P1_P1_InstQueueRd_Addr_PTR2), .A2(_02090__PTR6), .ZN(_02089__PTR32) );
  AND2_X1 U11880 ( .A1(P1_P1_InstQueueRd_Addr_PTR3), .A2(_02090__PTR6), .ZN(_02089__PTR33) );
  AND2_X1 U11881 ( .A1(P1_P1_InstQueueRd_Addr_PTR4), .A2(_02090__PTR6), .ZN(_02089__PTR34) );
  AND2_X1 U11882 ( .A1(_02088__PTR25), .A2(_02086__PTR4), .ZN(_02089__PTR25) );
  AND2_X1 U11883 ( .A1(_02088__PTR26), .A2(_02086__PTR4), .ZN(_02089__PTR26) );
  AND2_X1 U11884 ( .A1(_02088__PTR27), .A2(_02086__PTR4), .ZN(_02089__PTR27) );
  AND2_X1 U11885 ( .A1(_02088__PTR28), .A2(_02086__PTR4), .ZN(_02089__PTR28) );
  AND2_X1 U11886 ( .A1(_02088__PTR29), .A2(_02086__PTR4), .ZN(_02089__PTR29) );
  AND2_X1 U11887 ( .A1(P1_P1_InstQueueRd_Addr_PTR0), .A2(_02090__PTR4), .ZN(_02089__PTR20) );
  AND2_X1 U11888 ( .A1(_02088__PTR21), .A2(_02090__PTR4), .ZN(_02089__PTR21) );
  AND2_X1 U11889 ( .A1(_02088__PTR22), .A2(_02090__PTR4), .ZN(_02089__PTR22) );
  AND2_X1 U11890 ( .A1(_02088__PTR23), .A2(_02090__PTR4), .ZN(_02089__PTR23) );
  AND2_X1 U11891 ( .A1(_02088__PTR24), .A2(_02090__PTR4), .ZN(_02089__PTR24) );
  AND2_X1 U11892 ( .A1(P1_P1_InstQueueRd_Addr_PTR0), .A2(_02090__PTR3), .ZN(_02089__PTR15) );
  AND2_X1 U11893 ( .A1(_02088__PTR21), .A2(_02090__PTR3), .ZN(_02089__PTR16) );
  AND2_X1 U11894 ( .A1(_02088__PTR22), .A2(_02090__PTR3), .ZN(_02089__PTR17) );
  AND2_X1 U11895 ( .A1(_02088__PTR23), .A2(_02090__PTR3), .ZN(_02089__PTR18) );
  AND2_X1 U11896 ( .A1(_02088__PTR19), .A2(_02090__PTR3), .ZN(_02089__PTR19) );
  AND2_X1 U11897 ( .A1(P1_P1_InstQueueRd_Addr_PTR0), .A2(_01855__PTR0), .ZN(_02089__PTR10) );
  AND2_X1 U11898 ( .A1(_02088__PTR11), .A2(_01855__PTR0), .ZN(_02089__PTR11) );
  AND2_X1 U11899 ( .A1(_02088__PTR12), .A2(_01855__PTR0), .ZN(_02089__PTR12) );
  AND2_X1 U11900 ( .A1(_02088__PTR13), .A2(_01855__PTR0), .ZN(_02089__PTR13) );
  AND2_X1 U11901 ( .A1(_02088__PTR14), .A2(_01855__PTR0), .ZN(_02089__PTR14) );
  AND2_X1 U11902 ( .A1(P1_P1_InstQueueRd_Addr_PTR0), .A2(_02086__PTR1), .ZN(_02089__PTR5) );
  AND2_X1 U11903 ( .A1(_01890__PTR4), .A2(_02086__PTR1), .ZN(_02089__PTR6) );
  AND2_X1 U11904 ( .A1(_01890__PTR5), .A2(_02086__PTR1), .ZN(_02089__PTR7) );
  AND2_X1 U11905 ( .A1(_01890__PTR6), .A2(_02086__PTR1), .ZN(_02089__PTR8) );
  AND2_X1 U11906 ( .A1(_01884__PTR3), .A2(_02086__PTR0), .ZN(_02089__PTR0) );
  AND2_X1 U11907 ( .A1(_01884__PTR4), .A2(_02086__PTR0), .ZN(_02089__PTR1) );
  AND2_X1 U11908 ( .A1(_01884__PTR5), .A2(_02086__PTR0), .ZN(_02089__PTR2) );
  AND2_X1 U11909 ( .A1(_01884__PTR6), .A2(_02086__PTR0), .ZN(_02089__PTR3) );
  AND2_X1 U11910 ( .A1(P1_CodeFetch), .A2(_01863__PTR3), .ZN(_01873__PTR1) );
  AND2_X1 U11911 ( .A1(_01872__PTR0), .A2(_01874__PTR0), .ZN(_01873__PTR0) );
  AND2_X1 U11912 ( .A1(_01861__PTR0), .A2(_01863__PTR0), .ZN(_01862__PTR0) );
  AND2_X1 U11913 ( .A1(_01861__PTR1), .A2(_01855__PTR1), .ZN(_01862__PTR1) );
  AND2_X1 U11914 ( .A1(_01861__PTR2), .A2(_01863__PTR2), .ZN(_01862__PTR2) );
  AND2_X1 U11915 ( .A1(P1_RequestPending), .A2(_01863__PTR3), .ZN(_01862__PTR3) );
  AND2_X1 U11916 ( .A1(P1_MemoryFetch), .A2(_01863__PTR3), .ZN(_01869__PTR2) );
  AND2_X1 U11917 ( .A1(_01868__PTR1), .A2(_01870__PTR1), .ZN(_01869__PTR1) );
  AND2_X1 U11918 ( .A1(_01868__PTR0), .A2(_01870__PTR0), .ZN(_01869__PTR0) );
  AND2_X1 U11919 ( .A1(_01865__PTR0), .A2(_01855__PTR0), .ZN(_01866__PTR0) );
  AND2_X1 U11920 ( .A1(_01865__PTR1), .A2(_01855__PTR1), .ZN(_01866__PTR1) );
  AND2_X1 U11921 ( .A1(P1_ReadRequest), .A2(_01863__PTR3), .ZN(_01866__PTR2) );
  AND2_X1 U11922 ( .A1(_02104__PTR96), .A2(_02090__PTR4), .ZN(_02105__PTR96) );
  AND2_X1 U11923 ( .A1(_02104__PTR97), .A2(_02090__PTR4), .ZN(_02105__PTR97) );
  AND2_X1 U11924 ( .A1(_02104__PTR98), .A2(_02090__PTR4), .ZN(_02105__PTR98) );
  AND2_X1 U11925 ( .A1(_02104__PTR99), .A2(_02090__PTR4), .ZN(_02105__PTR99) );
  AND2_X1 U11926 ( .A1(_02104__PTR100), .A2(_02090__PTR4), .ZN(_02105__PTR100) );
  AND2_X1 U11927 ( .A1(_02104__PTR101), .A2(_02090__PTR4), .ZN(_02105__PTR101) );
  AND2_X1 U11928 ( .A1(_02104__PTR102), .A2(_02090__PTR4), .ZN(_02105__PTR102) );
  AND2_X1 U11929 ( .A1(_02104__PTR103), .A2(_02090__PTR4), .ZN(_02105__PTR103) );
  AND2_X1 U11930 ( .A1(_02104__PTR104), .A2(_02090__PTR4), .ZN(_02105__PTR104) );
  AND2_X1 U11931 ( .A1(_02104__PTR105), .A2(_02090__PTR4), .ZN(_02105__PTR105) );
  AND2_X1 U11932 ( .A1(_02104__PTR106), .A2(_02090__PTR4), .ZN(_02105__PTR106) );
  AND2_X1 U11933 ( .A1(_02104__PTR107), .A2(_02090__PTR4), .ZN(_02105__PTR107) );
  AND2_X1 U11934 ( .A1(_02104__PTR108), .A2(_02090__PTR4), .ZN(_02105__PTR108) );
  AND2_X1 U11935 ( .A1(_02104__PTR109), .A2(_02090__PTR4), .ZN(_02105__PTR109) );
  AND2_X1 U11936 ( .A1(_02104__PTR110), .A2(_02090__PTR4), .ZN(_02105__PTR110) );
  AND2_X1 U11937 ( .A1(_02104__PTR111), .A2(_02090__PTR4), .ZN(_02105__PTR111) );
  AND2_X1 U11938 ( .A1(_02104__PTR112), .A2(_02090__PTR4), .ZN(_02105__PTR112) );
  AND2_X1 U11939 ( .A1(_02104__PTR113), .A2(_02090__PTR4), .ZN(_02105__PTR113) );
  AND2_X1 U11940 ( .A1(_02104__PTR114), .A2(_02090__PTR4), .ZN(_02105__PTR114) );
  AND2_X1 U11941 ( .A1(_02104__PTR115), .A2(_02090__PTR4), .ZN(_02105__PTR115) );
  AND2_X1 U11942 ( .A1(_02104__PTR116), .A2(_02090__PTR4), .ZN(_02105__PTR116) );
  AND2_X1 U11943 ( .A1(_02104__PTR117), .A2(_02090__PTR4), .ZN(_02105__PTR117) );
  AND2_X1 U11944 ( .A1(_02104__PTR118), .A2(_02090__PTR4), .ZN(_02105__PTR118) );
  AND2_X1 U11945 ( .A1(_02104__PTR119), .A2(_02090__PTR4), .ZN(_02105__PTR119) );
  AND2_X1 U11946 ( .A1(_02104__PTR120), .A2(_02090__PTR4), .ZN(_02105__PTR120) );
  AND2_X1 U11947 ( .A1(_02104__PTR121), .A2(_02090__PTR4), .ZN(_02105__PTR121) );
  AND2_X1 U11948 ( .A1(_02104__PTR122), .A2(_02090__PTR4), .ZN(_02105__PTR122) );
  AND2_X1 U11949 ( .A1(_02104__PTR123), .A2(_02090__PTR4), .ZN(_02105__PTR123) );
  AND2_X1 U11950 ( .A1(_02104__PTR124), .A2(_02090__PTR4), .ZN(_02105__PTR124) );
  AND2_X1 U11951 ( .A1(_02104__PTR125), .A2(_02090__PTR4), .ZN(_02105__PTR125) );
  AND2_X1 U11952 ( .A1(_02104__PTR126), .A2(_02090__PTR4), .ZN(_02105__PTR126) );
  AND2_X1 U11953 ( .A1(_02104__PTR127), .A2(_02090__PTR4), .ZN(_02105__PTR127) );
  AND2_X1 U11954 ( .A1(_02104__PTR64), .A2(_01863__PTR2), .ZN(_02105__PTR64) );
  AND2_X1 U11955 ( .A1(_02104__PTR65), .A2(_01863__PTR2), .ZN(_02105__PTR65) );
  AND2_X1 U11956 ( .A1(_02104__PTR66), .A2(_01863__PTR2), .ZN(_02105__PTR66) );
  AND2_X1 U11957 ( .A1(_02104__PTR67), .A2(_01863__PTR2), .ZN(_02105__PTR67) );
  AND2_X1 U11958 ( .A1(_02104__PTR68), .A2(_01863__PTR2), .ZN(_02105__PTR68) );
  AND2_X1 U11959 ( .A1(_02104__PTR69), .A2(_01863__PTR2), .ZN(_02105__PTR69) );
  AND2_X1 U11960 ( .A1(_02104__PTR70), .A2(_01863__PTR2), .ZN(_02105__PTR70) );
  AND2_X1 U11961 ( .A1(_02104__PTR71), .A2(_01863__PTR2), .ZN(_02105__PTR71) );
  AND2_X1 U11962 ( .A1(_02104__PTR72), .A2(_01863__PTR2), .ZN(_02105__PTR72) );
  AND2_X1 U11963 ( .A1(_02104__PTR73), .A2(_01863__PTR2), .ZN(_02105__PTR73) );
  AND2_X1 U11964 ( .A1(_02104__PTR74), .A2(_01863__PTR2), .ZN(_02105__PTR74) );
  AND2_X1 U11965 ( .A1(_02104__PTR75), .A2(_01863__PTR2), .ZN(_02105__PTR75) );
  AND2_X1 U11966 ( .A1(_02104__PTR76), .A2(_01863__PTR2), .ZN(_02105__PTR76) );
  AND2_X1 U11967 ( .A1(_02104__PTR77), .A2(_01863__PTR2), .ZN(_02105__PTR77) );
  AND2_X1 U11968 ( .A1(_02104__PTR78), .A2(_01863__PTR2), .ZN(_02105__PTR78) );
  AND2_X1 U11969 ( .A1(_02104__PTR79), .A2(_01863__PTR2), .ZN(_02105__PTR79) );
  AND2_X1 U11970 ( .A1(_02104__PTR80), .A2(_01863__PTR2), .ZN(_02105__PTR80) );
  AND2_X1 U11971 ( .A1(_02104__PTR81), .A2(_01863__PTR2), .ZN(_02105__PTR81) );
  AND2_X1 U11972 ( .A1(_02104__PTR82), .A2(_01863__PTR2), .ZN(_02105__PTR82) );
  AND2_X1 U11973 ( .A1(_02104__PTR83), .A2(_01863__PTR2), .ZN(_02105__PTR83) );
  AND2_X1 U11974 ( .A1(_02104__PTR84), .A2(_01863__PTR2), .ZN(_02105__PTR84) );
  AND2_X1 U11975 ( .A1(_02104__PTR85), .A2(_01863__PTR2), .ZN(_02105__PTR85) );
  AND2_X1 U11976 ( .A1(_02104__PTR86), .A2(_01863__PTR2), .ZN(_02105__PTR86) );
  AND2_X1 U11977 ( .A1(_02104__PTR87), .A2(_01863__PTR2), .ZN(_02105__PTR87) );
  AND2_X1 U11978 ( .A1(_02104__PTR88), .A2(_01863__PTR2), .ZN(_02105__PTR88) );
  AND2_X1 U11979 ( .A1(_02104__PTR89), .A2(_01863__PTR2), .ZN(_02105__PTR89) );
  AND2_X1 U11980 ( .A1(_02104__PTR90), .A2(_01863__PTR2), .ZN(_02105__PTR90) );
  AND2_X1 U11981 ( .A1(_02104__PTR91), .A2(_01863__PTR2), .ZN(_02105__PTR91) );
  AND2_X1 U11982 ( .A1(_02104__PTR92), .A2(_01863__PTR2), .ZN(_02105__PTR92) );
  AND2_X1 U11983 ( .A1(_02104__PTR93), .A2(_01863__PTR2), .ZN(_02105__PTR93) );
  AND2_X1 U11984 ( .A1(_02104__PTR94), .A2(_01863__PTR2), .ZN(_02105__PTR94) );
  AND2_X1 U11985 ( .A1(_02104__PTR95), .A2(_01863__PTR2), .ZN(_02105__PTR95) );
  AND2_X1 U11986 ( .A1(_02104__PTR32), .A2(_01870__PTR0), .ZN(_02105__PTR32) );
  AND2_X1 U11987 ( .A1(_02104__PTR33), .A2(_01870__PTR0), .ZN(_02105__PTR33) );
  AND2_X1 U11988 ( .A1(_02104__PTR34), .A2(_01870__PTR0), .ZN(_02105__PTR34) );
  AND2_X1 U11989 ( .A1(_02104__PTR35), .A2(_01870__PTR0), .ZN(_02105__PTR35) );
  AND2_X1 U11990 ( .A1(_02104__PTR36), .A2(_01870__PTR0), .ZN(_02105__PTR36) );
  AND2_X1 U11991 ( .A1(_02104__PTR37), .A2(_01870__PTR0), .ZN(_02105__PTR37) );
  AND2_X1 U11992 ( .A1(_02104__PTR38), .A2(_01870__PTR0), .ZN(_02105__PTR38) );
  AND2_X1 U11993 ( .A1(_02104__PTR39), .A2(_01870__PTR0), .ZN(_02105__PTR39) );
  AND2_X1 U11994 ( .A1(_02104__PTR40), .A2(_01870__PTR0), .ZN(_02105__PTR40) );
  AND2_X1 U11995 ( .A1(_02104__PTR41), .A2(_01870__PTR0), .ZN(_02105__PTR41) );
  AND2_X1 U11996 ( .A1(_02104__PTR42), .A2(_01870__PTR0), .ZN(_02105__PTR42) );
  AND2_X1 U11997 ( .A1(_02104__PTR43), .A2(_01870__PTR0), .ZN(_02105__PTR43) );
  AND2_X1 U11998 ( .A1(_02104__PTR44), .A2(_01870__PTR0), .ZN(_02105__PTR44) );
  AND2_X1 U11999 ( .A1(_02104__PTR45), .A2(_01870__PTR0), .ZN(_02105__PTR45) );
  AND2_X1 U12000 ( .A1(_02104__PTR46), .A2(_01870__PTR0), .ZN(_02105__PTR46) );
  AND2_X1 U12001 ( .A1(_02104__PTR47), .A2(_01870__PTR0), .ZN(_02105__PTR47) );
  AND2_X1 U12002 ( .A1(_02104__PTR48), .A2(_01870__PTR0), .ZN(_02105__PTR48) );
  AND2_X1 U12003 ( .A1(_02104__PTR49), .A2(_01870__PTR0), .ZN(_02105__PTR49) );
  AND2_X1 U12004 ( .A1(_02104__PTR50), .A2(_01870__PTR0), .ZN(_02105__PTR50) );
  AND2_X1 U12005 ( .A1(_02104__PTR51), .A2(_01870__PTR0), .ZN(_02105__PTR51) );
  AND2_X1 U12006 ( .A1(_02104__PTR52), .A2(_01870__PTR0), .ZN(_02105__PTR52) );
  AND2_X1 U12007 ( .A1(_02104__PTR53), .A2(_01870__PTR0), .ZN(_02105__PTR53) );
  AND2_X1 U12008 ( .A1(_02104__PTR54), .A2(_01870__PTR0), .ZN(_02105__PTR54) );
  AND2_X1 U12009 ( .A1(_02104__PTR55), .A2(_01870__PTR0), .ZN(_02105__PTR55) );
  AND2_X1 U12010 ( .A1(_02104__PTR56), .A2(_01870__PTR0), .ZN(_02105__PTR56) );
  AND2_X1 U12011 ( .A1(_02104__PTR57), .A2(_01870__PTR0), .ZN(_02105__PTR57) );
  AND2_X1 U12012 ( .A1(_02104__PTR58), .A2(_01870__PTR0), .ZN(_02105__PTR58) );
  AND2_X1 U12013 ( .A1(_02104__PTR59), .A2(_01870__PTR0), .ZN(_02105__PTR59) );
  AND2_X1 U12014 ( .A1(_02104__PTR60), .A2(_01870__PTR0), .ZN(_02105__PTR60) );
  AND2_X1 U12015 ( .A1(_02104__PTR61), .A2(_01870__PTR0), .ZN(_02105__PTR61) );
  AND2_X1 U12016 ( .A1(_02104__PTR62), .A2(_01870__PTR0), .ZN(_02105__PTR62) );
  AND2_X1 U12017 ( .A1(_02104__PTR63), .A2(_01870__PTR0), .ZN(_02105__PTR63) );
  AND2_X1 U12018 ( .A1(P1_rEIP_PTR0), .A2(_01863__PTR3), .ZN(_02105__PTR0) );
  AND2_X1 U12019 ( .A1(P1_rEIP_PTR1), .A2(_01863__PTR3), .ZN(_02105__PTR1) );
  AND2_X1 U12020 ( .A1(P1_rEIP_PTR2), .A2(_01863__PTR3), .ZN(_02105__PTR2) );
  AND2_X1 U12021 ( .A1(P1_rEIP_PTR3), .A2(_01863__PTR3), .ZN(_02105__PTR3) );
  AND2_X1 U12022 ( .A1(P1_rEIP_PTR4), .A2(_01863__PTR3), .ZN(_02105__PTR4) );
  AND2_X1 U12023 ( .A1(P1_rEIP_PTR5), .A2(_01863__PTR3), .ZN(_02105__PTR5) );
  AND2_X1 U12024 ( .A1(P1_rEIP_PTR6), .A2(_01863__PTR3), .ZN(_02105__PTR6) );
  AND2_X1 U12025 ( .A1(P1_rEIP_PTR7), .A2(_01863__PTR3), .ZN(_02105__PTR7) );
  AND2_X1 U12026 ( .A1(P1_rEIP_PTR8), .A2(_01863__PTR3), .ZN(_02105__PTR8) );
  AND2_X1 U12027 ( .A1(P1_rEIP_PTR9), .A2(_01863__PTR3), .ZN(_02105__PTR9) );
  AND2_X1 U12028 ( .A1(P1_rEIP_PTR10), .A2(_01863__PTR3), .ZN(_02105__PTR10) );
  AND2_X1 U12029 ( .A1(P1_rEIP_PTR11), .A2(_01863__PTR3), .ZN(_02105__PTR11) );
  AND2_X1 U12030 ( .A1(P1_rEIP_PTR12), .A2(_01863__PTR3), .ZN(_02105__PTR12) );
  AND2_X1 U12031 ( .A1(P1_rEIP_PTR13), .A2(_01863__PTR3), .ZN(_02105__PTR13) );
  AND2_X1 U12032 ( .A1(P1_rEIP_PTR14), .A2(_01863__PTR3), .ZN(_02105__PTR14) );
  AND2_X1 U12033 ( .A1(P1_rEIP_PTR15), .A2(_01863__PTR3), .ZN(_02105__PTR15) );
  AND2_X1 U12034 ( .A1(P1_rEIP_PTR16), .A2(_01863__PTR3), .ZN(_02105__PTR16) );
  AND2_X1 U12035 ( .A1(P1_rEIP_PTR17), .A2(_01863__PTR3), .ZN(_02105__PTR17) );
  AND2_X1 U12036 ( .A1(P1_rEIP_PTR18), .A2(_01863__PTR3), .ZN(_02105__PTR18) );
  AND2_X1 U12037 ( .A1(P1_rEIP_PTR19), .A2(_01863__PTR3), .ZN(_02105__PTR19) );
  AND2_X1 U12038 ( .A1(P1_rEIP_PTR20), .A2(_01863__PTR3), .ZN(_02105__PTR20) );
  AND2_X1 U12039 ( .A1(P1_rEIP_PTR21), .A2(_01863__PTR3), .ZN(_02105__PTR21) );
  AND2_X1 U12040 ( .A1(P1_rEIP_PTR22), .A2(_01863__PTR3), .ZN(_02105__PTR22) );
  AND2_X1 U12041 ( .A1(P1_rEIP_PTR23), .A2(_01863__PTR3), .ZN(_02105__PTR23) );
  AND2_X1 U12042 ( .A1(P1_rEIP_PTR24), .A2(_01863__PTR3), .ZN(_02105__PTR24) );
  AND2_X1 U12043 ( .A1(P1_rEIP_PTR25), .A2(_01863__PTR3), .ZN(_02105__PTR25) );
  AND2_X1 U12044 ( .A1(P1_rEIP_PTR26), .A2(_01863__PTR3), .ZN(_02105__PTR26) );
  AND2_X1 U12045 ( .A1(P1_rEIP_PTR27), .A2(_01863__PTR3), .ZN(_02105__PTR27) );
  AND2_X1 U12046 ( .A1(P1_rEIP_PTR28), .A2(_01863__PTR3), .ZN(_02105__PTR28) );
  AND2_X1 U12047 ( .A1(P1_rEIP_PTR29), .A2(_01863__PTR3), .ZN(_02105__PTR29) );
  AND2_X1 U12048 ( .A1(P1_rEIP_PTR30), .A2(_01863__PTR3), .ZN(_02105__PTR30) );
  AND2_X1 U12049 ( .A1(P1_rEIP_PTR31), .A2(_01863__PTR3), .ZN(_02105__PTR31) );
  AND2_X1 U12050 ( .A1(_02084__PTR192), .A2(_01855__PTR3), .ZN(_02085__PTR192) );
  AND2_X1 U12051 ( .A1(_02084__PTR193), .A2(_01855__PTR3), .ZN(_02085__PTR193) );
  AND2_X1 U12052 ( .A1(_02084__PTR194), .A2(_01855__PTR3), .ZN(_02085__PTR194) );
  AND2_X1 U12053 ( .A1(_02084__PTR195), .A2(_01855__PTR3), .ZN(_02085__PTR195) );
  AND2_X1 U12054 ( .A1(_02084__PTR196), .A2(_01855__PTR3), .ZN(_02085__PTR196) );
  AND2_X1 U12055 ( .A1(_02084__PTR197), .A2(_01855__PTR3), .ZN(_02085__PTR197) );
  AND2_X1 U12056 ( .A1(_02084__PTR198), .A2(_01855__PTR3), .ZN(_02085__PTR198) );
  AND2_X1 U12057 ( .A1(_02084__PTR199), .A2(_01855__PTR3), .ZN(_02085__PTR199) );
  AND2_X1 U12058 ( .A1(_02084__PTR200), .A2(_01855__PTR3), .ZN(_02085__PTR200) );
  AND2_X1 U12059 ( .A1(_02084__PTR201), .A2(_01855__PTR3), .ZN(_02085__PTR201) );
  AND2_X1 U12060 ( .A1(_02084__PTR202), .A2(_01855__PTR3), .ZN(_02085__PTR202) );
  AND2_X1 U12061 ( .A1(_02084__PTR203), .A2(_01855__PTR3), .ZN(_02085__PTR203) );
  AND2_X1 U12062 ( .A1(_02084__PTR204), .A2(_01855__PTR3), .ZN(_02085__PTR204) );
  AND2_X1 U12063 ( .A1(_02084__PTR205), .A2(_01855__PTR3), .ZN(_02085__PTR205) );
  AND2_X1 U12064 ( .A1(_02084__PTR206), .A2(_01855__PTR3), .ZN(_02085__PTR206) );
  AND2_X1 U12065 ( .A1(_02084__PTR207), .A2(_01855__PTR3), .ZN(_02085__PTR207) );
  AND2_X1 U12066 ( .A1(_02084__PTR208), .A2(_01855__PTR3), .ZN(_02085__PTR208) );
  AND2_X1 U12067 ( .A1(_02084__PTR209), .A2(_01855__PTR3), .ZN(_02085__PTR209) );
  AND2_X1 U12068 ( .A1(_02084__PTR210), .A2(_01855__PTR3), .ZN(_02085__PTR210) );
  AND2_X1 U12069 ( .A1(_02084__PTR211), .A2(_01855__PTR3), .ZN(_02085__PTR211) );
  AND2_X1 U12070 ( .A1(_02084__PTR212), .A2(_01855__PTR3), .ZN(_02085__PTR212) );
  AND2_X1 U12071 ( .A1(_02084__PTR213), .A2(_01855__PTR3), .ZN(_02085__PTR213) );
  AND2_X1 U12072 ( .A1(_02084__PTR214), .A2(_01855__PTR3), .ZN(_02085__PTR214) );
  AND2_X1 U12073 ( .A1(_02084__PTR215), .A2(_01855__PTR3), .ZN(_02085__PTR215) );
  AND2_X1 U12074 ( .A1(_02084__PTR216), .A2(_01855__PTR3), .ZN(_02085__PTR216) );
  AND2_X1 U12075 ( .A1(_02084__PTR217), .A2(_01855__PTR3), .ZN(_02085__PTR217) );
  AND2_X1 U12076 ( .A1(_02084__PTR218), .A2(_01855__PTR3), .ZN(_02085__PTR218) );
  AND2_X1 U12077 ( .A1(_02084__PTR219), .A2(_01855__PTR3), .ZN(_02085__PTR219) );
  AND2_X1 U12078 ( .A1(_02084__PTR220), .A2(_01855__PTR3), .ZN(_02085__PTR220) );
  AND2_X1 U12079 ( .A1(_02084__PTR221), .A2(_01855__PTR3), .ZN(_02085__PTR221) );
  AND2_X1 U12080 ( .A1(_02084__PTR222), .A2(_01855__PTR3), .ZN(_02085__PTR222) );
  AND2_X1 U12081 ( .A1(_02084__PTR223), .A2(_01855__PTR3), .ZN(_02085__PTR223) );
  AND2_X1 U12082 ( .A1(_02084__PTR160), .A2(_01855__PTR2), .ZN(_02085__PTR160) );
  AND2_X1 U12083 ( .A1(_02084__PTR161), .A2(_01855__PTR2), .ZN(_02085__PTR161) );
  AND2_X1 U12084 ( .A1(_02084__PTR162), .A2(_01855__PTR2), .ZN(_02085__PTR162) );
  AND2_X1 U12085 ( .A1(_02084__PTR163), .A2(_01855__PTR2), .ZN(_02085__PTR163) );
  AND2_X1 U12086 ( .A1(_02084__PTR164), .A2(_01855__PTR2), .ZN(_02085__PTR164) );
  AND2_X1 U12087 ( .A1(_02084__PTR165), .A2(_01855__PTR2), .ZN(_02085__PTR165) );
  AND2_X1 U12088 ( .A1(_02084__PTR166), .A2(_01855__PTR2), .ZN(_02085__PTR166) );
  AND2_X1 U12089 ( .A1(_02084__PTR167), .A2(_01855__PTR2), .ZN(_02085__PTR167) );
  AND2_X1 U12090 ( .A1(_02084__PTR168), .A2(_01855__PTR2), .ZN(_02085__PTR168) );
  AND2_X1 U12091 ( .A1(_02084__PTR169), .A2(_01855__PTR2), .ZN(_02085__PTR169) );
  AND2_X1 U12092 ( .A1(_02084__PTR170), .A2(_01855__PTR2), .ZN(_02085__PTR170) );
  AND2_X1 U12093 ( .A1(_02084__PTR171), .A2(_01855__PTR2), .ZN(_02085__PTR171) );
  AND2_X1 U12094 ( .A1(_02084__PTR172), .A2(_01855__PTR2), .ZN(_02085__PTR172) );
  AND2_X1 U12095 ( .A1(_02084__PTR173), .A2(_01855__PTR2), .ZN(_02085__PTR173) );
  AND2_X1 U12096 ( .A1(_02084__PTR174), .A2(_01855__PTR2), .ZN(_02085__PTR174) );
  AND2_X1 U12097 ( .A1(_02084__PTR175), .A2(_01855__PTR2), .ZN(_02085__PTR175) );
  AND2_X1 U12098 ( .A1(_02084__PTR176), .A2(_01855__PTR2), .ZN(_02085__PTR176) );
  AND2_X1 U12099 ( .A1(_02084__PTR177), .A2(_01855__PTR2), .ZN(_02085__PTR177) );
  AND2_X1 U12100 ( .A1(_02084__PTR178), .A2(_01855__PTR2), .ZN(_02085__PTR178) );
  AND2_X1 U12101 ( .A1(_02084__PTR179), .A2(_01855__PTR2), .ZN(_02085__PTR179) );
  AND2_X1 U12102 ( .A1(_02084__PTR180), .A2(_01855__PTR2), .ZN(_02085__PTR180) );
  AND2_X1 U12103 ( .A1(_02084__PTR181), .A2(_01855__PTR2), .ZN(_02085__PTR181) );
  AND2_X1 U12104 ( .A1(_02084__PTR182), .A2(_01855__PTR2), .ZN(_02085__PTR182) );
  AND2_X1 U12105 ( .A1(_02084__PTR183), .A2(_01855__PTR2), .ZN(_02085__PTR183) );
  AND2_X1 U12106 ( .A1(_02084__PTR184), .A2(_01855__PTR2), .ZN(_02085__PTR184) );
  AND2_X1 U12107 ( .A1(_02084__PTR185), .A2(_01855__PTR2), .ZN(_02085__PTR185) );
  AND2_X1 U12108 ( .A1(_02084__PTR186), .A2(_01855__PTR2), .ZN(_02085__PTR186) );
  AND2_X1 U12109 ( .A1(_02084__PTR187), .A2(_01855__PTR2), .ZN(_02085__PTR187) );
  AND2_X1 U12110 ( .A1(_02084__PTR188), .A2(_01855__PTR2), .ZN(_02085__PTR188) );
  AND2_X1 U12111 ( .A1(_02084__PTR189), .A2(_01855__PTR2), .ZN(_02085__PTR189) );
  AND2_X1 U12112 ( .A1(_02084__PTR190), .A2(_01855__PTR2), .ZN(_02085__PTR190) );
  AND2_X1 U12113 ( .A1(_02084__PTR191), .A2(_01855__PTR2), .ZN(_02085__PTR191) );
  AND2_X1 U12114 ( .A1(_02084__PTR128), .A2(_02086__PTR4), .ZN(_02085__PTR128) );
  AND2_X1 U12115 ( .A1(_02084__PTR129), .A2(_02086__PTR4), .ZN(_02085__PTR129) );
  AND2_X1 U12116 ( .A1(_02084__PTR130), .A2(_02086__PTR4), .ZN(_02085__PTR130) );
  AND2_X1 U12117 ( .A1(_02084__PTR131), .A2(_02086__PTR4), .ZN(_02085__PTR131) );
  AND2_X1 U12118 ( .A1(_02084__PTR132), .A2(_02086__PTR4), .ZN(_02085__PTR132) );
  AND2_X1 U12119 ( .A1(_02084__PTR133), .A2(_02086__PTR4), .ZN(_02085__PTR133) );
  AND2_X1 U12120 ( .A1(_02084__PTR134), .A2(_02086__PTR4), .ZN(_02085__PTR134) );
  AND2_X1 U12121 ( .A1(_02084__PTR135), .A2(_02086__PTR4), .ZN(_02085__PTR135) );
  AND2_X1 U12122 ( .A1(_02084__PTR136), .A2(_02086__PTR4), .ZN(_02085__PTR136) );
  AND2_X1 U12123 ( .A1(_02084__PTR137), .A2(_02086__PTR4), .ZN(_02085__PTR137) );
  AND2_X1 U12124 ( .A1(_02084__PTR138), .A2(_02086__PTR4), .ZN(_02085__PTR138) );
  AND2_X1 U12125 ( .A1(_02084__PTR139), .A2(_02086__PTR4), .ZN(_02085__PTR139) );
  AND2_X1 U12126 ( .A1(_02084__PTR140), .A2(_02086__PTR4), .ZN(_02085__PTR140) );
  AND2_X1 U12127 ( .A1(_02084__PTR141), .A2(_02086__PTR4), .ZN(_02085__PTR141) );
  AND2_X1 U12128 ( .A1(_02084__PTR142), .A2(_02086__PTR4), .ZN(_02085__PTR142) );
  AND2_X1 U12129 ( .A1(_02084__PTR143), .A2(_02086__PTR4), .ZN(_02085__PTR143) );
  AND2_X1 U12130 ( .A1(_02084__PTR144), .A2(_02086__PTR4), .ZN(_02085__PTR144) );
  AND2_X1 U12131 ( .A1(_02084__PTR145), .A2(_02086__PTR4), .ZN(_02085__PTR145) );
  AND2_X1 U12132 ( .A1(_02084__PTR146), .A2(_02086__PTR4), .ZN(_02085__PTR146) );
  AND2_X1 U12133 ( .A1(_02084__PTR147), .A2(_02086__PTR4), .ZN(_02085__PTR147) );
  AND2_X1 U12134 ( .A1(_02084__PTR148), .A2(_02086__PTR4), .ZN(_02085__PTR148) );
  AND2_X1 U12135 ( .A1(_02084__PTR149), .A2(_02086__PTR4), .ZN(_02085__PTR149) );
  AND2_X1 U12136 ( .A1(_02084__PTR150), .A2(_02086__PTR4), .ZN(_02085__PTR150) );
  AND2_X1 U12137 ( .A1(_02084__PTR151), .A2(_02086__PTR4), .ZN(_02085__PTR151) );
  AND2_X1 U12138 ( .A1(_02084__PTR152), .A2(_02086__PTR4), .ZN(_02085__PTR152) );
  AND2_X1 U12139 ( .A1(_02084__PTR153), .A2(_02086__PTR4), .ZN(_02085__PTR153) );
  AND2_X1 U12140 ( .A1(_02084__PTR154), .A2(_02086__PTR4), .ZN(_02085__PTR154) );
  AND2_X1 U12141 ( .A1(_02084__PTR155), .A2(_02086__PTR4), .ZN(_02085__PTR155) );
  AND2_X1 U12142 ( .A1(_02084__PTR156), .A2(_02086__PTR4), .ZN(_02085__PTR156) );
  AND2_X1 U12143 ( .A1(_02084__PTR157), .A2(_02086__PTR4), .ZN(_02085__PTR157) );
  AND2_X1 U12144 ( .A1(_02084__PTR158), .A2(_02086__PTR4), .ZN(_02085__PTR158) );
  AND2_X1 U12145 ( .A1(_02084__PTR159), .A2(_02086__PTR4), .ZN(_02085__PTR159) );
  AND2_X1 U12146 ( .A1(P1_P1_InstAddrPointer_PTR0), .A2(_01855__PTR1), .ZN(_02085__PTR96) );
  AND2_X1 U12147 ( .A1(_02084__PTR97), .A2(_01855__PTR1), .ZN(_02085__PTR97) );
  AND2_X1 U12148 ( .A1(_02084__PTR98), .A2(_01855__PTR1), .ZN(_02085__PTR98) );
  AND2_X1 U12149 ( .A1(_02084__PTR99), .A2(_01855__PTR1), .ZN(_02085__PTR99) );
  AND2_X1 U12150 ( .A1(_02084__PTR100), .A2(_01855__PTR1), .ZN(_02085__PTR100) );
  AND2_X1 U12151 ( .A1(_02084__PTR101), .A2(_01855__PTR1), .ZN(_02085__PTR101) );
  AND2_X1 U12152 ( .A1(_02084__PTR102), .A2(_01855__PTR1), .ZN(_02085__PTR102) );
  AND2_X1 U12153 ( .A1(_02084__PTR103), .A2(_01855__PTR1), .ZN(_02085__PTR103) );
  AND2_X1 U12154 ( .A1(_02084__PTR104), .A2(_01855__PTR1), .ZN(_02085__PTR104) );
  AND2_X1 U12155 ( .A1(_02084__PTR105), .A2(_01855__PTR1), .ZN(_02085__PTR105) );
  AND2_X1 U12156 ( .A1(_02084__PTR106), .A2(_01855__PTR1), .ZN(_02085__PTR106) );
  AND2_X1 U12157 ( .A1(_02084__PTR107), .A2(_01855__PTR1), .ZN(_02085__PTR107) );
  AND2_X1 U12158 ( .A1(_02084__PTR108), .A2(_01855__PTR1), .ZN(_02085__PTR108) );
  AND2_X1 U12159 ( .A1(_02084__PTR109), .A2(_01855__PTR1), .ZN(_02085__PTR109) );
  AND2_X1 U12160 ( .A1(_02084__PTR110), .A2(_01855__PTR1), .ZN(_02085__PTR110) );
  AND2_X1 U12161 ( .A1(_02084__PTR111), .A2(_01855__PTR1), .ZN(_02085__PTR111) );
  AND2_X1 U12162 ( .A1(_02084__PTR112), .A2(_01855__PTR1), .ZN(_02085__PTR112) );
  AND2_X1 U12163 ( .A1(_02084__PTR113), .A2(_01855__PTR1), .ZN(_02085__PTR113) );
  AND2_X1 U12164 ( .A1(_02084__PTR114), .A2(_01855__PTR1), .ZN(_02085__PTR114) );
  AND2_X1 U12165 ( .A1(_02084__PTR115), .A2(_01855__PTR1), .ZN(_02085__PTR115) );
  AND2_X1 U12166 ( .A1(_02084__PTR116), .A2(_01855__PTR1), .ZN(_02085__PTR116) );
  AND2_X1 U12167 ( .A1(_02084__PTR117), .A2(_01855__PTR1), .ZN(_02085__PTR117) );
  AND2_X1 U12168 ( .A1(_02084__PTR118), .A2(_01855__PTR1), .ZN(_02085__PTR118) );
  AND2_X1 U12169 ( .A1(_02084__PTR119), .A2(_01855__PTR1), .ZN(_02085__PTR119) );
  AND2_X1 U12170 ( .A1(_02084__PTR120), .A2(_01855__PTR1), .ZN(_02085__PTR120) );
  AND2_X1 U12171 ( .A1(_02084__PTR121), .A2(_01855__PTR1), .ZN(_02085__PTR121) );
  AND2_X1 U12172 ( .A1(_02084__PTR122), .A2(_01855__PTR1), .ZN(_02085__PTR122) );
  AND2_X1 U12173 ( .A1(_02084__PTR123), .A2(_01855__PTR1), .ZN(_02085__PTR123) );
  AND2_X1 U12174 ( .A1(_02084__PTR124), .A2(_01855__PTR1), .ZN(_02085__PTR124) );
  AND2_X1 U12175 ( .A1(_02084__PTR125), .A2(_01855__PTR1), .ZN(_02085__PTR125) );
  AND2_X1 U12176 ( .A1(_02084__PTR126), .A2(_01855__PTR1), .ZN(_02085__PTR126) );
  AND2_X1 U12177 ( .A1(_02084__PTR127), .A2(_01855__PTR1), .ZN(_02085__PTR127) );
  AND2_X1 U12178 ( .A1(P1_P1_InstAddrPointer_PTR0), .A2(_01855__PTR0), .ZN(_02085__PTR64) );
  AND2_X1 U12179 ( .A1(_02084__PTR65), .A2(_01855__PTR0), .ZN(_02085__PTR65) );
  AND2_X1 U12180 ( .A1(_02084__PTR66), .A2(_01855__PTR0), .ZN(_02085__PTR66) );
  AND2_X1 U12181 ( .A1(_02084__PTR67), .A2(_01855__PTR0), .ZN(_02085__PTR67) );
  AND2_X1 U12182 ( .A1(_02084__PTR68), .A2(_01855__PTR0), .ZN(_02085__PTR68) );
  AND2_X1 U12183 ( .A1(_02084__PTR69), .A2(_01855__PTR0), .ZN(_02085__PTR69) );
  AND2_X1 U12184 ( .A1(_02084__PTR70), .A2(_01855__PTR0), .ZN(_02085__PTR70) );
  AND2_X1 U12185 ( .A1(_02084__PTR71), .A2(_01855__PTR0), .ZN(_02085__PTR71) );
  AND2_X1 U12186 ( .A1(_02084__PTR72), .A2(_01855__PTR0), .ZN(_02085__PTR72) );
  AND2_X1 U12187 ( .A1(_02084__PTR73), .A2(_01855__PTR0), .ZN(_02085__PTR73) );
  AND2_X1 U12188 ( .A1(_02084__PTR74), .A2(_01855__PTR0), .ZN(_02085__PTR74) );
  AND2_X1 U12189 ( .A1(_02084__PTR75), .A2(_01855__PTR0), .ZN(_02085__PTR75) );
  AND2_X1 U12190 ( .A1(_02084__PTR76), .A2(_01855__PTR0), .ZN(_02085__PTR76) );
  AND2_X1 U12191 ( .A1(_02084__PTR77), .A2(_01855__PTR0), .ZN(_02085__PTR77) );
  AND2_X1 U12192 ( .A1(_02084__PTR78), .A2(_01855__PTR0), .ZN(_02085__PTR78) );
  AND2_X1 U12193 ( .A1(_02084__PTR79), .A2(_01855__PTR0), .ZN(_02085__PTR79) );
  AND2_X1 U12194 ( .A1(_02084__PTR80), .A2(_01855__PTR0), .ZN(_02085__PTR80) );
  AND2_X1 U12195 ( .A1(_02084__PTR81), .A2(_01855__PTR0), .ZN(_02085__PTR81) );
  AND2_X1 U12196 ( .A1(_02084__PTR82), .A2(_01855__PTR0), .ZN(_02085__PTR82) );
  AND2_X1 U12197 ( .A1(_02084__PTR83), .A2(_01855__PTR0), .ZN(_02085__PTR83) );
  AND2_X1 U12198 ( .A1(_02084__PTR84), .A2(_01855__PTR0), .ZN(_02085__PTR84) );
  AND2_X1 U12199 ( .A1(_02084__PTR85), .A2(_01855__PTR0), .ZN(_02085__PTR85) );
  AND2_X1 U12200 ( .A1(_02084__PTR86), .A2(_01855__PTR0), .ZN(_02085__PTR86) );
  AND2_X1 U12201 ( .A1(_02084__PTR87), .A2(_01855__PTR0), .ZN(_02085__PTR87) );
  AND2_X1 U12202 ( .A1(_02084__PTR88), .A2(_01855__PTR0), .ZN(_02085__PTR88) );
  AND2_X1 U12203 ( .A1(_02084__PTR89), .A2(_01855__PTR0), .ZN(_02085__PTR89) );
  AND2_X1 U12204 ( .A1(_02084__PTR90), .A2(_01855__PTR0), .ZN(_02085__PTR90) );
  AND2_X1 U12205 ( .A1(_02084__PTR91), .A2(_01855__PTR0), .ZN(_02085__PTR91) );
  AND2_X1 U12206 ( .A1(_02084__PTR92), .A2(_01855__PTR0), .ZN(_02085__PTR92) );
  AND2_X1 U12207 ( .A1(_02084__PTR93), .A2(_01855__PTR0), .ZN(_02085__PTR93) );
  AND2_X1 U12208 ( .A1(_02084__PTR94), .A2(_01855__PTR0), .ZN(_02085__PTR94) );
  AND2_X1 U12209 ( .A1(_02084__PTR95), .A2(_01855__PTR0), .ZN(_02085__PTR95) );
  AND2_X1 U12210 ( .A1(P1_P1_InstAddrPointer_PTR0), .A2(_02086__PTR1), .ZN(_02085__PTR32) );
  AND2_X1 U12211 ( .A1(_02084__PTR33), .A2(_02086__PTR1), .ZN(_02085__PTR33) );
  AND2_X1 U12212 ( .A1(_02084__PTR34), .A2(_02086__PTR1), .ZN(_02085__PTR34) );
  AND2_X1 U12213 ( .A1(_02084__PTR35), .A2(_02086__PTR1), .ZN(_02085__PTR35) );
  AND2_X1 U12214 ( .A1(_02084__PTR36), .A2(_02086__PTR1), .ZN(_02085__PTR36) );
  AND2_X1 U12215 ( .A1(_02084__PTR37), .A2(_02086__PTR1), .ZN(_02085__PTR37) );
  AND2_X1 U12216 ( .A1(_02084__PTR38), .A2(_02086__PTR1), .ZN(_02085__PTR38) );
  AND2_X1 U12217 ( .A1(_02084__PTR39), .A2(_02086__PTR1), .ZN(_02085__PTR39) );
  AND2_X1 U12218 ( .A1(_02084__PTR40), .A2(_02086__PTR1), .ZN(_02085__PTR40) );
  AND2_X1 U12219 ( .A1(_02084__PTR41), .A2(_02086__PTR1), .ZN(_02085__PTR41) );
  AND2_X1 U12220 ( .A1(_02084__PTR42), .A2(_02086__PTR1), .ZN(_02085__PTR42) );
  AND2_X1 U12221 ( .A1(_02084__PTR43), .A2(_02086__PTR1), .ZN(_02085__PTR43) );
  AND2_X1 U12222 ( .A1(_02084__PTR44), .A2(_02086__PTR1), .ZN(_02085__PTR44) );
  AND2_X1 U12223 ( .A1(_02084__PTR45), .A2(_02086__PTR1), .ZN(_02085__PTR45) );
  AND2_X1 U12224 ( .A1(_02084__PTR46), .A2(_02086__PTR1), .ZN(_02085__PTR46) );
  AND2_X1 U12225 ( .A1(_02084__PTR47), .A2(_02086__PTR1), .ZN(_02085__PTR47) );
  AND2_X1 U12226 ( .A1(_02084__PTR48), .A2(_02086__PTR1), .ZN(_02085__PTR48) );
  AND2_X1 U12227 ( .A1(_02084__PTR49), .A2(_02086__PTR1), .ZN(_02085__PTR49) );
  AND2_X1 U12228 ( .A1(_02084__PTR50), .A2(_02086__PTR1), .ZN(_02085__PTR50) );
  AND2_X1 U12229 ( .A1(_02084__PTR51), .A2(_02086__PTR1), .ZN(_02085__PTR51) );
  AND2_X1 U12230 ( .A1(_02084__PTR52), .A2(_02086__PTR1), .ZN(_02085__PTR52) );
  AND2_X1 U12231 ( .A1(_02084__PTR53), .A2(_02086__PTR1), .ZN(_02085__PTR53) );
  AND2_X1 U12232 ( .A1(_02084__PTR54), .A2(_02086__PTR1), .ZN(_02085__PTR54) );
  AND2_X1 U12233 ( .A1(_02084__PTR55), .A2(_02086__PTR1), .ZN(_02085__PTR55) );
  AND2_X1 U12234 ( .A1(_02084__PTR56), .A2(_02086__PTR1), .ZN(_02085__PTR56) );
  AND2_X1 U12235 ( .A1(_02084__PTR57), .A2(_02086__PTR1), .ZN(_02085__PTR57) );
  AND2_X1 U12236 ( .A1(_02084__PTR58), .A2(_02086__PTR1), .ZN(_02085__PTR58) );
  AND2_X1 U12237 ( .A1(_02084__PTR59), .A2(_02086__PTR1), .ZN(_02085__PTR59) );
  AND2_X1 U12238 ( .A1(_02084__PTR60), .A2(_02086__PTR1), .ZN(_02085__PTR60) );
  AND2_X1 U12239 ( .A1(_02084__PTR61), .A2(_02086__PTR1), .ZN(_02085__PTR61) );
  AND2_X1 U12240 ( .A1(_02084__PTR62), .A2(_02086__PTR1), .ZN(_02085__PTR62) );
  AND2_X1 U12241 ( .A1(_02084__PTR63), .A2(_02086__PTR1), .ZN(_02085__PTR63) );
  AND2_X1 U12242 ( .A1(_02084__PTR0), .A2(_02086__PTR0), .ZN(_02085__PTR0) );
  AND2_X1 U12243 ( .A1(_02084__PTR1), .A2(_02086__PTR0), .ZN(_02085__PTR1) );
  AND2_X1 U12244 ( .A1(_02084__PTR2), .A2(_02086__PTR0), .ZN(_02085__PTR2) );
  AND2_X1 U12245 ( .A1(_02084__PTR3), .A2(_02086__PTR0), .ZN(_02085__PTR3) );
  AND2_X1 U12246 ( .A1(_02084__PTR4), .A2(_02086__PTR0), .ZN(_02085__PTR4) );
  AND2_X1 U12247 ( .A1(_02084__PTR5), .A2(_02086__PTR0), .ZN(_02085__PTR5) );
  AND2_X1 U12248 ( .A1(_02084__PTR6), .A2(_02086__PTR0), .ZN(_02085__PTR6) );
  AND2_X1 U12249 ( .A1(_02084__PTR7), .A2(_02086__PTR0), .ZN(_02085__PTR7) );
  AND2_X1 U12250 ( .A1(_02084__PTR8), .A2(_02086__PTR0), .ZN(_02085__PTR8) );
  AND2_X1 U12251 ( .A1(_02084__PTR9), .A2(_02086__PTR0), .ZN(_02085__PTR9) );
  AND2_X1 U12252 ( .A1(_02084__PTR10), .A2(_02086__PTR0), .ZN(_02085__PTR10) );
  AND2_X1 U12253 ( .A1(_02084__PTR11), .A2(_02086__PTR0), .ZN(_02085__PTR11) );
  AND2_X1 U12254 ( .A1(_02084__PTR12), .A2(_02086__PTR0), .ZN(_02085__PTR12) );
  AND2_X1 U12255 ( .A1(_02084__PTR13), .A2(_02086__PTR0), .ZN(_02085__PTR13) );
  AND2_X1 U12256 ( .A1(_02084__PTR14), .A2(_02086__PTR0), .ZN(_02085__PTR14) );
  AND2_X1 U12257 ( .A1(_02084__PTR15), .A2(_02086__PTR0), .ZN(_02085__PTR15) );
  AND2_X1 U12258 ( .A1(_02084__PTR16), .A2(_02086__PTR0), .ZN(_02085__PTR16) );
  AND2_X1 U12259 ( .A1(_02084__PTR17), .A2(_02086__PTR0), .ZN(_02085__PTR17) );
  AND2_X1 U12260 ( .A1(_02084__PTR18), .A2(_02086__PTR0), .ZN(_02085__PTR18) );
  AND2_X1 U12261 ( .A1(_02084__PTR19), .A2(_02086__PTR0), .ZN(_02085__PTR19) );
  AND2_X1 U12262 ( .A1(_02084__PTR20), .A2(_02086__PTR0), .ZN(_02085__PTR20) );
  AND2_X1 U12263 ( .A1(_02084__PTR21), .A2(_02086__PTR0), .ZN(_02085__PTR21) );
  AND2_X1 U12264 ( .A1(_02084__PTR22), .A2(_02086__PTR0), .ZN(_02085__PTR22) );
  AND2_X1 U12265 ( .A1(_02084__PTR23), .A2(_02086__PTR0), .ZN(_02085__PTR23) );
  AND2_X1 U12266 ( .A1(_02084__PTR24), .A2(_02086__PTR0), .ZN(_02085__PTR24) );
  AND2_X1 U12267 ( .A1(_02084__PTR25), .A2(_02086__PTR0), .ZN(_02085__PTR25) );
  AND2_X1 U12268 ( .A1(_02084__PTR26), .A2(_02086__PTR0), .ZN(_02085__PTR26) );
  AND2_X1 U12269 ( .A1(_02084__PTR27), .A2(_02086__PTR0), .ZN(_02085__PTR27) );
  AND2_X1 U12270 ( .A1(_02084__PTR28), .A2(_02086__PTR0), .ZN(_02085__PTR28) );
  AND2_X1 U12271 ( .A1(_02084__PTR29), .A2(_02086__PTR0), .ZN(_02085__PTR29) );
  AND2_X1 U12272 ( .A1(_02084__PTR30), .A2(_02086__PTR0), .ZN(_02085__PTR30) );
  AND2_X1 U12273 ( .A1(_02084__PTR31), .A2(_02086__PTR0), .ZN(_02085__PTR31) );
  AND2_X1 U12274 ( .A1(P1_P1_PhyAddrPointer_PTR0), .A2(_02094__PTR0), .ZN(_02093__PTR0) );
  AND2_X1 U12275 ( .A1(P1_P1_PhyAddrPointer_PTR1), .A2(_02094__PTR0), .ZN(_02093__PTR1) );
  AND2_X1 U12276 ( .A1(P1_P1_PhyAddrPointer_PTR2), .A2(_02094__PTR0), .ZN(_02093__PTR2) );
  AND2_X1 U12277 ( .A1(P1_P1_PhyAddrPointer_PTR3), .A2(_02094__PTR0), .ZN(_02093__PTR3) );
  AND2_X1 U12278 ( .A1(P1_P1_PhyAddrPointer_PTR4), .A2(_02094__PTR0), .ZN(_02093__PTR4) );
  AND2_X1 U12279 ( .A1(P1_P1_PhyAddrPointer_PTR5), .A2(_02094__PTR0), .ZN(_02093__PTR5) );
  AND2_X1 U12280 ( .A1(P1_P1_PhyAddrPointer_PTR6), .A2(_02094__PTR0), .ZN(_02093__PTR6) );
  AND2_X1 U12281 ( .A1(P1_P1_PhyAddrPointer_PTR7), .A2(_02094__PTR0), .ZN(_02093__PTR7) );
  AND2_X1 U12282 ( .A1(P1_P1_PhyAddrPointer_PTR8), .A2(_02094__PTR0), .ZN(_02093__PTR8) );
  AND2_X1 U12283 ( .A1(P1_P1_PhyAddrPointer_PTR9), .A2(_02094__PTR0), .ZN(_02093__PTR9) );
  AND2_X1 U12284 ( .A1(P1_P1_PhyAddrPointer_PTR10), .A2(_02094__PTR0), .ZN(_02093__PTR10) );
  AND2_X1 U12285 ( .A1(P1_P1_PhyAddrPointer_PTR11), .A2(_02094__PTR0), .ZN(_02093__PTR11) );
  AND2_X1 U12286 ( .A1(P1_P1_PhyAddrPointer_PTR12), .A2(_02094__PTR0), .ZN(_02093__PTR12) );
  AND2_X1 U12287 ( .A1(P1_P1_PhyAddrPointer_PTR13), .A2(_02094__PTR0), .ZN(_02093__PTR13) );
  AND2_X1 U12288 ( .A1(P1_P1_PhyAddrPointer_PTR14), .A2(_02094__PTR0), .ZN(_02093__PTR14) );
  AND2_X1 U12289 ( .A1(P1_P1_PhyAddrPointer_PTR15), .A2(_02094__PTR0), .ZN(_02093__PTR15) );
  AND2_X1 U12290 ( .A1(P1_P1_PhyAddrPointer_PTR16), .A2(_02094__PTR0), .ZN(_02093__PTR16) );
  AND2_X1 U12291 ( .A1(P1_P1_PhyAddrPointer_PTR17), .A2(_02094__PTR0), .ZN(_02093__PTR17) );
  AND2_X1 U12292 ( .A1(P1_P1_PhyAddrPointer_PTR18), .A2(_02094__PTR0), .ZN(_02093__PTR18) );
  AND2_X1 U12293 ( .A1(P1_P1_PhyAddrPointer_PTR19), .A2(_02094__PTR0), .ZN(_02093__PTR19) );
  AND2_X1 U12294 ( .A1(P1_P1_PhyAddrPointer_PTR20), .A2(_02094__PTR0), .ZN(_02093__PTR20) );
  AND2_X1 U12295 ( .A1(P1_P1_PhyAddrPointer_PTR21), .A2(_02094__PTR0), .ZN(_02093__PTR21) );
  AND2_X1 U12296 ( .A1(P1_P1_PhyAddrPointer_PTR22), .A2(_02094__PTR0), .ZN(_02093__PTR22) );
  AND2_X1 U12297 ( .A1(P1_P1_PhyAddrPointer_PTR23), .A2(_02094__PTR0), .ZN(_02093__PTR23) );
  AND2_X1 U12298 ( .A1(P1_P1_PhyAddrPointer_PTR24), .A2(_02094__PTR0), .ZN(_02093__PTR24) );
  AND2_X1 U12299 ( .A1(P1_P1_PhyAddrPointer_PTR25), .A2(_02094__PTR0), .ZN(_02093__PTR25) );
  AND2_X1 U12300 ( .A1(P1_P1_PhyAddrPointer_PTR26), .A2(_02094__PTR0), .ZN(_02093__PTR26) );
  AND2_X1 U12301 ( .A1(P1_P1_PhyAddrPointer_PTR27), .A2(_02094__PTR0), .ZN(_02093__PTR27) );
  AND2_X1 U12302 ( .A1(P1_P1_PhyAddrPointer_PTR28), .A2(_02094__PTR0), .ZN(_02093__PTR28) );
  AND2_X1 U12303 ( .A1(P1_P1_PhyAddrPointer_PTR29), .A2(_02094__PTR0), .ZN(_02093__PTR29) );
  AND2_X1 U12304 ( .A1(P1_P1_PhyAddrPointer_PTR30), .A2(_02094__PTR0), .ZN(_02093__PTR30) );
  AND2_X1 U12305 ( .A1(P1_P1_PhyAddrPointer_PTR31), .A2(_02094__PTR0), .ZN(_02093__PTR31) );
  AND2_X1 U12306 ( .A1(_02092__PTR32), .A2(_01855__PTR2), .ZN(_02093__PTR32) );
  AND2_X1 U12307 ( .A1(_02092__PTR33), .A2(_01855__PTR2), .ZN(_02093__PTR33) );
  AND2_X1 U12308 ( .A1(_02092__PTR34), .A2(_01855__PTR2), .ZN(_02093__PTR34) );
  AND2_X1 U12309 ( .A1(_02092__PTR35), .A2(_01855__PTR2), .ZN(_02093__PTR35) );
  AND2_X1 U12310 ( .A1(_02092__PTR36), .A2(_01855__PTR2), .ZN(_02093__PTR36) );
  AND2_X1 U12311 ( .A1(_02092__PTR37), .A2(_01855__PTR2), .ZN(_02093__PTR37) );
  AND2_X1 U12312 ( .A1(_02092__PTR38), .A2(_01855__PTR2), .ZN(_02093__PTR38) );
  AND2_X1 U12313 ( .A1(_02092__PTR39), .A2(_01855__PTR2), .ZN(_02093__PTR39) );
  AND2_X1 U12314 ( .A1(_02092__PTR40), .A2(_01855__PTR2), .ZN(_02093__PTR40) );
  AND2_X1 U12315 ( .A1(_02092__PTR41), .A2(_01855__PTR2), .ZN(_02093__PTR41) );
  AND2_X1 U12316 ( .A1(_02092__PTR42), .A2(_01855__PTR2), .ZN(_02093__PTR42) );
  AND2_X1 U12317 ( .A1(_02092__PTR43), .A2(_01855__PTR2), .ZN(_02093__PTR43) );
  AND2_X1 U12318 ( .A1(_02092__PTR44), .A2(_01855__PTR2), .ZN(_02093__PTR44) );
  AND2_X1 U12319 ( .A1(_02092__PTR45), .A2(_01855__PTR2), .ZN(_02093__PTR45) );
  AND2_X1 U12320 ( .A1(_02092__PTR46), .A2(_01855__PTR2), .ZN(_02093__PTR46) );
  AND2_X1 U12321 ( .A1(_02092__PTR47), .A2(_01855__PTR2), .ZN(_02093__PTR47) );
  AND2_X1 U12322 ( .A1(_02092__PTR48), .A2(_01855__PTR2), .ZN(_02093__PTR48) );
  AND2_X1 U12323 ( .A1(_02092__PTR49), .A2(_01855__PTR2), .ZN(_02093__PTR49) );
  AND2_X1 U12324 ( .A1(_02092__PTR50), .A2(_01855__PTR2), .ZN(_02093__PTR50) );
  AND2_X1 U12325 ( .A1(_02092__PTR51), .A2(_01855__PTR2), .ZN(_02093__PTR51) );
  AND2_X1 U12326 ( .A1(_02092__PTR52), .A2(_01855__PTR2), .ZN(_02093__PTR52) );
  AND2_X1 U12327 ( .A1(_02092__PTR53), .A2(_01855__PTR2), .ZN(_02093__PTR53) );
  AND2_X1 U12328 ( .A1(_02092__PTR54), .A2(_01855__PTR2), .ZN(_02093__PTR54) );
  AND2_X1 U12329 ( .A1(_02092__PTR55), .A2(_01855__PTR2), .ZN(_02093__PTR55) );
  AND2_X1 U12330 ( .A1(_02092__PTR56), .A2(_01855__PTR2), .ZN(_02093__PTR56) );
  AND2_X1 U12331 ( .A1(_02092__PTR57), .A2(_01855__PTR2), .ZN(_02093__PTR57) );
  AND2_X1 U12332 ( .A1(_02092__PTR58), .A2(_01855__PTR2), .ZN(_02093__PTR58) );
  AND2_X1 U12333 ( .A1(_02092__PTR59), .A2(_01855__PTR2), .ZN(_02093__PTR59) );
  AND2_X1 U12334 ( .A1(_02092__PTR60), .A2(_01855__PTR2), .ZN(_02093__PTR60) );
  AND2_X1 U12335 ( .A1(_02092__PTR61), .A2(_01855__PTR2), .ZN(_02093__PTR61) );
  AND2_X1 U12336 ( .A1(_02092__PTR62), .A2(_01855__PTR2), .ZN(_02093__PTR62) );
  AND2_X1 U12337 ( .A1(_02092__PTR63), .A2(_01855__PTR2), .ZN(_02093__PTR63) );
  AND2_X1 U12338 ( .A1(_02092__PTR64), .A2(_01855__PTR3), .ZN(_02093__PTR64) );
  AND2_X1 U12339 ( .A1(_02092__PTR65), .A2(_01855__PTR3), .ZN(_02093__PTR65) );
  AND2_X1 U12340 ( .A1(_02092__PTR66), .A2(_01855__PTR3), .ZN(_02093__PTR66) );
  AND2_X1 U12341 ( .A1(_02092__PTR67), .A2(_01855__PTR3), .ZN(_02093__PTR67) );
  AND2_X1 U12342 ( .A1(_02092__PTR68), .A2(_01855__PTR3), .ZN(_02093__PTR68) );
  AND2_X1 U12343 ( .A1(_02092__PTR69), .A2(_01855__PTR3), .ZN(_02093__PTR69) );
  AND2_X1 U12344 ( .A1(_02092__PTR70), .A2(_01855__PTR3), .ZN(_02093__PTR70) );
  AND2_X1 U12345 ( .A1(_02092__PTR71), .A2(_01855__PTR3), .ZN(_02093__PTR71) );
  AND2_X1 U12346 ( .A1(_02092__PTR72), .A2(_01855__PTR3), .ZN(_02093__PTR72) );
  AND2_X1 U12347 ( .A1(_02092__PTR73), .A2(_01855__PTR3), .ZN(_02093__PTR73) );
  AND2_X1 U12348 ( .A1(_02092__PTR74), .A2(_01855__PTR3), .ZN(_02093__PTR74) );
  AND2_X1 U12349 ( .A1(_02092__PTR75), .A2(_01855__PTR3), .ZN(_02093__PTR75) );
  AND2_X1 U12350 ( .A1(_02092__PTR76), .A2(_01855__PTR3), .ZN(_02093__PTR76) );
  AND2_X1 U12351 ( .A1(_02092__PTR77), .A2(_01855__PTR3), .ZN(_02093__PTR77) );
  AND2_X1 U12352 ( .A1(_02092__PTR78), .A2(_01855__PTR3), .ZN(_02093__PTR78) );
  AND2_X1 U12353 ( .A1(_02092__PTR79), .A2(_01855__PTR3), .ZN(_02093__PTR79) );
  AND2_X1 U12354 ( .A1(_02092__PTR80), .A2(_01855__PTR3), .ZN(_02093__PTR80) );
  AND2_X1 U12355 ( .A1(_02092__PTR81), .A2(_01855__PTR3), .ZN(_02093__PTR81) );
  AND2_X1 U12356 ( .A1(_02092__PTR82), .A2(_01855__PTR3), .ZN(_02093__PTR82) );
  AND2_X1 U12357 ( .A1(_02092__PTR83), .A2(_01855__PTR3), .ZN(_02093__PTR83) );
  AND2_X1 U12358 ( .A1(_02092__PTR84), .A2(_01855__PTR3), .ZN(_02093__PTR84) );
  AND2_X1 U12359 ( .A1(_02092__PTR85), .A2(_01855__PTR3), .ZN(_02093__PTR85) );
  AND2_X1 U12360 ( .A1(_02092__PTR86), .A2(_01855__PTR3), .ZN(_02093__PTR86) );
  AND2_X1 U12361 ( .A1(_02092__PTR87), .A2(_01855__PTR3), .ZN(_02093__PTR87) );
  AND2_X1 U12362 ( .A1(_02092__PTR88), .A2(_01855__PTR3), .ZN(_02093__PTR88) );
  AND2_X1 U12363 ( .A1(_02092__PTR89), .A2(_01855__PTR3), .ZN(_02093__PTR89) );
  AND2_X1 U12364 ( .A1(_02092__PTR90), .A2(_01855__PTR3), .ZN(_02093__PTR90) );
  AND2_X1 U12365 ( .A1(_02092__PTR91), .A2(_01855__PTR3), .ZN(_02093__PTR91) );
  AND2_X1 U12366 ( .A1(_02092__PTR92), .A2(_01855__PTR3), .ZN(_02093__PTR92) );
  AND2_X1 U12367 ( .A1(_02092__PTR93), .A2(_01855__PTR3), .ZN(_02093__PTR93) );
  AND2_X1 U12368 ( .A1(_02092__PTR94), .A2(_01855__PTR3), .ZN(_02093__PTR94) );
  AND2_X1 U12369 ( .A1(_02092__PTR95), .A2(_01855__PTR3), .ZN(_02093__PTR95) );
  AND2_X1 U12370 ( .A1(_02118__PTR4), .A2(_01863__PTR2), .ZN(_02119__PTR4) );
  AND2_X1 U12371 ( .A1(_02118__PTR5), .A2(_01863__PTR2), .ZN(_02119__PTR5) );
  AND2_X1 U12372 ( .A1(_02118__PTR6), .A2(_01863__PTR2), .ZN(_02119__PTR6) );
  AND2_X1 U12373 ( .A1(_02118__PTR7), .A2(_01863__PTR2), .ZN(_02119__PTR7) );
  AND2_X1 U12374 ( .A1(P1_P1_State2_PTR0), .A2(_02120__PTR0), .ZN(_02119__PTR0) );
  AND2_X1 U12375 ( .A1(P1_P1_State2_PTR1), .A2(_02120__PTR0), .ZN(_02119__PTR1) );
  AND2_X1 U12376 ( .A1(P1_P1_State2_PTR2), .A2(_02120__PTR0), .ZN(_02119__PTR2) );
  AND2_X1 U12377 ( .A1(P1_P1_State2_PTR3), .A2(_02120__PTR0), .ZN(_02119__PTR3) );
  AND2_X1 U12378 ( .A1(_02174__PTR8), .A2(_02413__PTR1), .ZN(_02412__PTR4) );
  AND2_X1 U12379 ( .A1(P2_rEIP_PTR1), .A2(_02413__PTR1), .ZN(_02412__PTR5) );
  AND2_X1 U12380 ( .A1(_02174__PTR2), .A2(_02413__PTR1), .ZN(_02412__PTR6) );
  AND2_X1 U12381 ( .A1(_02174__PTR8), .A2(_02413__PTR2), .ZN(_02412__PTR8) );
  AND2_X1 U12382 ( .A1(P2_rEIP_PTR1), .A2(_02413__PTR2), .ZN(_02412__PTR9) );
  AND2_X1 U12383 ( .A1(_02174__PTR6), .A2(_02413__PTR2), .ZN(_02412__PTR10) );
  AND2_X1 U12384 ( .A1(_02174__PTR7), .A2(_02413__PTR2), .ZN(_02412__PTR11) );
  AND2_X1 U12385 ( .A1(_02174__PTR8), .A2(_02413__PTR3), .ZN(_02412__PTR12) );
  AND2_X1 U12386 ( .A1(_02174__PTR9), .A2(_02413__PTR3), .ZN(_02412__PTR13) );
  AND2_X1 U12387 ( .A1(_02174__PTR10), .A2(_02413__PTR3), .ZN(_02412__PTR14) );
  AND2_X1 U12388 ( .A1(_02174__PTR11), .A2(_02413__PTR3), .ZN(_02412__PTR15) );
  AND2_X1 U12389 ( .A1(P2_Datao_PTR0), .A2(_02405__PTR0), .ZN(_02404__PTR0) );
  AND2_X1 U12390 ( .A1(P2_Datao_PTR1), .A2(_02405__PTR0), .ZN(_02404__PTR1) );
  AND2_X1 U12391 ( .A1(P2_Datao_PTR2), .A2(_02405__PTR0), .ZN(_02404__PTR2) );
  AND2_X1 U12392 ( .A1(P2_Datao_PTR3), .A2(_02405__PTR0), .ZN(_02404__PTR3) );
  AND2_X1 U12393 ( .A1(P2_Datao_PTR4), .A2(_02405__PTR0), .ZN(_02404__PTR4) );
  AND2_X1 U12394 ( .A1(P2_Datao_PTR5), .A2(_02405__PTR0), .ZN(_02404__PTR5) );
  AND2_X1 U12395 ( .A1(P2_Datao_PTR6), .A2(_02405__PTR0), .ZN(_02404__PTR6) );
  AND2_X1 U12396 ( .A1(P2_Datao_PTR7), .A2(_02405__PTR0), .ZN(_02404__PTR7) );
  AND2_X1 U12397 ( .A1(P2_Datao_PTR8), .A2(_02405__PTR0), .ZN(_02404__PTR8) );
  AND2_X1 U12398 ( .A1(P2_Datao_PTR9), .A2(_02405__PTR0), .ZN(_02404__PTR9) );
  AND2_X1 U12399 ( .A1(P2_Datao_PTR10), .A2(_02405__PTR0), .ZN(_02404__PTR10) );
  AND2_X1 U12400 ( .A1(P2_Datao_PTR11), .A2(_02405__PTR0), .ZN(_02404__PTR11) );
  AND2_X1 U12401 ( .A1(P2_Datao_PTR12), .A2(_02405__PTR0), .ZN(_02404__PTR12) );
  AND2_X1 U12402 ( .A1(P2_Datao_PTR13), .A2(_02405__PTR0), .ZN(_02404__PTR13) );
  AND2_X1 U12403 ( .A1(P2_Datao_PTR14), .A2(_02405__PTR0), .ZN(_02404__PTR14) );
  AND2_X1 U12404 ( .A1(P2_Datao_PTR15), .A2(_02405__PTR0), .ZN(_02404__PTR15) );
  AND2_X1 U12405 ( .A1(P2_Datao_PTR16), .A2(_02405__PTR0), .ZN(_02404__PTR16) );
  AND2_X1 U12406 ( .A1(P2_Datao_PTR17), .A2(_02405__PTR0), .ZN(_02404__PTR17) );
  AND2_X1 U12407 ( .A1(P2_Datao_PTR18), .A2(_02405__PTR0), .ZN(_02404__PTR18) );
  AND2_X1 U12408 ( .A1(P2_Datao_PTR19), .A2(_02405__PTR0), .ZN(_02404__PTR19) );
  AND2_X1 U12409 ( .A1(P2_Datao_PTR20), .A2(_02405__PTR0), .ZN(_02404__PTR20) );
  AND2_X1 U12410 ( .A1(P2_Datao_PTR21), .A2(_02405__PTR0), .ZN(_02404__PTR21) );
  AND2_X1 U12411 ( .A1(P2_Datao_PTR22), .A2(_02405__PTR0), .ZN(_02404__PTR22) );
  AND2_X1 U12412 ( .A1(P2_Datao_PTR23), .A2(_02405__PTR0), .ZN(_02404__PTR23) );
  AND2_X1 U12413 ( .A1(P2_Datao_PTR24), .A2(_02405__PTR0), .ZN(_02404__PTR24) );
  AND2_X1 U12414 ( .A1(P2_Datao_PTR25), .A2(_02405__PTR0), .ZN(_02404__PTR25) );
  AND2_X1 U12415 ( .A1(P2_Datao_PTR26), .A2(_02405__PTR0), .ZN(_02404__PTR26) );
  AND2_X1 U12416 ( .A1(P2_Datao_PTR27), .A2(_02405__PTR0), .ZN(_02404__PTR27) );
  AND2_X1 U12417 ( .A1(P2_Datao_PTR28), .A2(_02405__PTR0), .ZN(_02404__PTR28) );
  AND2_X1 U12418 ( .A1(P2_Datao_PTR29), .A2(_02405__PTR0), .ZN(_02404__PTR29) );
  AND2_X1 U12419 ( .A1(P2_Datao_PTR30), .A2(_02405__PTR0), .ZN(_02404__PTR30) );
  AND2_X1 U12420 ( .A1(P2_Datao_PTR31), .A2(_02405__PTR0), .ZN(_02404__PTR31) );
  AND2_X1 U12421 ( .A1(_02403__PTR64), .A2(_02156__PTR0), .ZN(_02404__PTR32) );
  AND2_X1 U12422 ( .A1(_02403__PTR65), .A2(_02156__PTR0), .ZN(_02404__PTR33) );
  AND2_X1 U12423 ( .A1(_02403__PTR66), .A2(_02156__PTR0), .ZN(_02404__PTR34) );
  AND2_X1 U12424 ( .A1(_02403__PTR67), .A2(_02156__PTR0), .ZN(_02404__PTR35) );
  AND2_X1 U12425 ( .A1(_02403__PTR68), .A2(_02156__PTR0), .ZN(_02404__PTR36) );
  AND2_X1 U12426 ( .A1(_02403__PTR69), .A2(_02156__PTR0), .ZN(_02404__PTR37) );
  AND2_X1 U12427 ( .A1(_02403__PTR70), .A2(_02156__PTR0), .ZN(_02404__PTR38) );
  AND2_X1 U12428 ( .A1(_02403__PTR71), .A2(_02156__PTR0), .ZN(_02404__PTR39) );
  AND2_X1 U12429 ( .A1(_02403__PTR72), .A2(_02156__PTR0), .ZN(_02404__PTR40) );
  AND2_X1 U12430 ( .A1(_02403__PTR73), .A2(_02156__PTR0), .ZN(_02404__PTR41) );
  AND2_X1 U12431 ( .A1(_02403__PTR74), .A2(_02156__PTR0), .ZN(_02404__PTR42) );
  AND2_X1 U12432 ( .A1(_02403__PTR75), .A2(_02156__PTR0), .ZN(_02404__PTR43) );
  AND2_X1 U12433 ( .A1(_02403__PTR76), .A2(_02156__PTR0), .ZN(_02404__PTR44) );
  AND2_X1 U12434 ( .A1(_02403__PTR77), .A2(_02156__PTR0), .ZN(_02404__PTR45) );
  AND2_X1 U12435 ( .A1(_02403__PTR78), .A2(_02156__PTR0), .ZN(_02404__PTR46) );
  AND2_X1 U12436 ( .A1(_02403__PTR79), .A2(_02156__PTR0), .ZN(_02404__PTR47) );
  AND2_X1 U12437 ( .A1(_02403__PTR48), .A2(_02156__PTR0), .ZN(_02404__PTR48) );
  AND2_X1 U12438 ( .A1(_02403__PTR49), .A2(_02156__PTR0), .ZN(_02404__PTR49) );
  AND2_X1 U12439 ( .A1(_02403__PTR50), .A2(_02156__PTR0), .ZN(_02404__PTR50) );
  AND2_X1 U12440 ( .A1(_02403__PTR51), .A2(_02156__PTR0), .ZN(_02404__PTR51) );
  AND2_X1 U12441 ( .A1(_02403__PTR52), .A2(_02156__PTR0), .ZN(_02404__PTR52) );
  AND2_X1 U12442 ( .A1(_02403__PTR53), .A2(_02156__PTR0), .ZN(_02404__PTR53) );
  AND2_X1 U12443 ( .A1(_02403__PTR54), .A2(_02156__PTR0), .ZN(_02404__PTR54) );
  AND2_X1 U12444 ( .A1(_02403__PTR55), .A2(_02156__PTR0), .ZN(_02404__PTR55) );
  AND2_X1 U12445 ( .A1(_02403__PTR56), .A2(_02156__PTR0), .ZN(_02404__PTR56) );
  AND2_X1 U12446 ( .A1(_02403__PTR57), .A2(_02156__PTR0), .ZN(_02404__PTR57) );
  AND2_X1 U12447 ( .A1(_02403__PTR58), .A2(_02156__PTR0), .ZN(_02404__PTR58) );
  AND2_X1 U12448 ( .A1(_02403__PTR59), .A2(_02156__PTR0), .ZN(_02404__PTR59) );
  AND2_X1 U12449 ( .A1(_02403__PTR60), .A2(_02156__PTR0), .ZN(_02404__PTR60) );
  AND2_X1 U12450 ( .A1(_02403__PTR61), .A2(_02156__PTR0), .ZN(_02404__PTR61) );
  AND2_X1 U12451 ( .A1(_02403__PTR62), .A2(_02156__PTR0), .ZN(_02404__PTR62) );
  AND2_X1 U12452 ( .A1(_02403__PTR95), .A2(_02156__PTR0), .ZN(_02404__PTR63) );
  AND2_X1 U12453 ( .A1(_02403__PTR64), .A2(_02156__PTR2), .ZN(_02404__PTR64) );
  AND2_X1 U12454 ( .A1(_02403__PTR65), .A2(_02156__PTR2), .ZN(_02404__PTR65) );
  AND2_X1 U12455 ( .A1(_02403__PTR66), .A2(_02156__PTR2), .ZN(_02404__PTR66) );
  AND2_X1 U12456 ( .A1(_02403__PTR67), .A2(_02156__PTR2), .ZN(_02404__PTR67) );
  AND2_X1 U12457 ( .A1(_02403__PTR68), .A2(_02156__PTR2), .ZN(_02404__PTR68) );
  AND2_X1 U12458 ( .A1(_02403__PTR69), .A2(_02156__PTR2), .ZN(_02404__PTR69) );
  AND2_X1 U12459 ( .A1(_02403__PTR70), .A2(_02156__PTR2), .ZN(_02404__PTR70) );
  AND2_X1 U12460 ( .A1(_02403__PTR71), .A2(_02156__PTR2), .ZN(_02404__PTR71) );
  AND2_X1 U12461 ( .A1(_02403__PTR72), .A2(_02156__PTR2), .ZN(_02404__PTR72) );
  AND2_X1 U12462 ( .A1(_02403__PTR73), .A2(_02156__PTR2), .ZN(_02404__PTR73) );
  AND2_X1 U12463 ( .A1(_02403__PTR74), .A2(_02156__PTR2), .ZN(_02404__PTR74) );
  AND2_X1 U12464 ( .A1(_02403__PTR75), .A2(_02156__PTR2), .ZN(_02404__PTR75) );
  AND2_X1 U12465 ( .A1(_02403__PTR76), .A2(_02156__PTR2), .ZN(_02404__PTR76) );
  AND2_X1 U12466 ( .A1(_02403__PTR77), .A2(_02156__PTR2), .ZN(_02404__PTR77) );
  AND2_X1 U12467 ( .A1(_02403__PTR78), .A2(_02156__PTR2), .ZN(_02404__PTR78) );
  AND2_X1 U12468 ( .A1(_02403__PTR79), .A2(_02156__PTR2), .ZN(_02404__PTR79) );
  AND2_X1 U12469 ( .A1(_02403__PTR80), .A2(_02156__PTR2), .ZN(_02404__PTR80) );
  AND2_X1 U12470 ( .A1(_02403__PTR81), .A2(_02156__PTR2), .ZN(_02404__PTR81) );
  AND2_X1 U12471 ( .A1(_02403__PTR82), .A2(_02156__PTR2), .ZN(_02404__PTR82) );
  AND2_X1 U12472 ( .A1(_02403__PTR83), .A2(_02156__PTR2), .ZN(_02404__PTR83) );
  AND2_X1 U12473 ( .A1(_02403__PTR84), .A2(_02156__PTR2), .ZN(_02404__PTR84) );
  AND2_X1 U12474 ( .A1(_02403__PTR85), .A2(_02156__PTR2), .ZN(_02404__PTR85) );
  AND2_X1 U12475 ( .A1(_02403__PTR86), .A2(_02156__PTR2), .ZN(_02404__PTR86) );
  AND2_X1 U12476 ( .A1(_02403__PTR87), .A2(_02156__PTR2), .ZN(_02404__PTR87) );
  AND2_X1 U12477 ( .A1(_02403__PTR88), .A2(_02156__PTR2), .ZN(_02404__PTR88) );
  AND2_X1 U12478 ( .A1(_02403__PTR89), .A2(_02156__PTR2), .ZN(_02404__PTR89) );
  AND2_X1 U12479 ( .A1(_02403__PTR90), .A2(_02156__PTR2), .ZN(_02404__PTR90) );
  AND2_X1 U12480 ( .A1(_02403__PTR91), .A2(_02156__PTR2), .ZN(_02404__PTR91) );
  AND2_X1 U12481 ( .A1(_02403__PTR92), .A2(_02156__PTR2), .ZN(_02404__PTR92) );
  AND2_X1 U12482 ( .A1(_02403__PTR93), .A2(_02156__PTR2), .ZN(_02404__PTR93) );
  AND2_X1 U12483 ( .A1(_02403__PTR94), .A2(_02156__PTR2), .ZN(_02404__PTR94) );
  AND2_X1 U12484 ( .A1(_02403__PTR95), .A2(_02156__PTR2), .ZN(_02404__PTR95) );
  AND2_X1 U12485 ( .A1(P2_P1_lWord_PTR0), .A2(_02398__PTR0), .ZN(_02401__PTR0) );
  AND2_X1 U12486 ( .A1(P2_P1_lWord_PTR1), .A2(_02398__PTR0), .ZN(_02401__PTR1) );
  AND2_X1 U12487 ( .A1(P2_P1_lWord_PTR2), .A2(_02398__PTR0), .ZN(_02401__PTR2) );
  AND2_X1 U12488 ( .A1(P2_P1_lWord_PTR3), .A2(_02398__PTR0), .ZN(_02401__PTR3) );
  AND2_X1 U12489 ( .A1(P2_P1_lWord_PTR4), .A2(_02398__PTR0), .ZN(_02401__PTR4) );
  AND2_X1 U12490 ( .A1(P2_P1_lWord_PTR5), .A2(_02398__PTR0), .ZN(_02401__PTR5) );
  AND2_X1 U12491 ( .A1(P2_P1_lWord_PTR6), .A2(_02398__PTR0), .ZN(_02401__PTR6) );
  AND2_X1 U12492 ( .A1(P2_P1_lWord_PTR7), .A2(_02398__PTR0), .ZN(_02401__PTR7) );
  AND2_X1 U12493 ( .A1(P2_P1_lWord_PTR8), .A2(_02398__PTR0), .ZN(_02401__PTR8) );
  AND2_X1 U12494 ( .A1(P2_P1_lWord_PTR9), .A2(_02398__PTR0), .ZN(_02401__PTR9) );
  AND2_X1 U12495 ( .A1(P2_P1_lWord_PTR10), .A2(_02398__PTR0), .ZN(_02401__PTR10) );
  AND2_X1 U12496 ( .A1(P2_P1_lWord_PTR11), .A2(_02398__PTR0), .ZN(_02401__PTR11) );
  AND2_X1 U12497 ( .A1(P2_P1_lWord_PTR12), .A2(_02398__PTR0), .ZN(_02401__PTR12) );
  AND2_X1 U12498 ( .A1(P2_P1_lWord_PTR13), .A2(_02398__PTR0), .ZN(_02401__PTR13) );
  AND2_X1 U12499 ( .A1(P2_P1_lWord_PTR14), .A2(_02398__PTR0), .ZN(_02401__PTR14) );
  AND2_X1 U12500 ( .A1(P2_P1_lWord_PTR15), .A2(_02398__PTR0), .ZN(_02401__PTR15) );
  AND2_X1 U12501 ( .A1(_02400__PTR16), .A2(_02156__PTR2), .ZN(_02401__PTR16) );
  AND2_X1 U12502 ( .A1(_02400__PTR17), .A2(_02156__PTR2), .ZN(_02401__PTR17) );
  AND2_X1 U12503 ( .A1(_02400__PTR18), .A2(_02156__PTR2), .ZN(_02401__PTR18) );
  AND2_X1 U12504 ( .A1(_02400__PTR19), .A2(_02156__PTR2), .ZN(_02401__PTR19) );
  AND2_X1 U12505 ( .A1(_02400__PTR20), .A2(_02156__PTR2), .ZN(_02401__PTR20) );
  AND2_X1 U12506 ( .A1(_02400__PTR21), .A2(_02156__PTR2), .ZN(_02401__PTR21) );
  AND2_X1 U12507 ( .A1(_02400__PTR22), .A2(_02156__PTR2), .ZN(_02401__PTR22) );
  AND2_X1 U12508 ( .A1(_02400__PTR23), .A2(_02156__PTR2), .ZN(_02401__PTR23) );
  AND2_X1 U12509 ( .A1(_02400__PTR24), .A2(_02156__PTR2), .ZN(_02401__PTR24) );
  AND2_X1 U12510 ( .A1(_02400__PTR25), .A2(_02156__PTR2), .ZN(_02401__PTR25) );
  AND2_X1 U12511 ( .A1(_02400__PTR26), .A2(_02156__PTR2), .ZN(_02401__PTR26) );
  AND2_X1 U12512 ( .A1(_02400__PTR27), .A2(_02156__PTR2), .ZN(_02401__PTR27) );
  AND2_X1 U12513 ( .A1(_02400__PTR28), .A2(_02156__PTR2), .ZN(_02401__PTR28) );
  AND2_X1 U12514 ( .A1(_02400__PTR29), .A2(_02156__PTR2), .ZN(_02401__PTR29) );
  AND2_X1 U12515 ( .A1(_02400__PTR30), .A2(_02156__PTR2), .ZN(_02401__PTR30) );
  AND2_X1 U12516 ( .A1(_02400__PTR31), .A2(_02156__PTR2), .ZN(_02401__PTR31) );
  AND2_X1 U12517 ( .A1(_02400__PTR32), .A2(_02379__PTR4), .ZN(_02401__PTR32) );
  AND2_X1 U12518 ( .A1(_02400__PTR33), .A2(_02379__PTR4), .ZN(_02401__PTR33) );
  AND2_X1 U12519 ( .A1(_02400__PTR34), .A2(_02379__PTR4), .ZN(_02401__PTR34) );
  AND2_X1 U12520 ( .A1(_02400__PTR35), .A2(_02379__PTR4), .ZN(_02401__PTR35) );
  AND2_X1 U12521 ( .A1(_02400__PTR36), .A2(_02379__PTR4), .ZN(_02401__PTR36) );
  AND2_X1 U12522 ( .A1(_02400__PTR37), .A2(_02379__PTR4), .ZN(_02401__PTR37) );
  AND2_X1 U12523 ( .A1(_02400__PTR38), .A2(_02379__PTR4), .ZN(_02401__PTR38) );
  AND2_X1 U12524 ( .A1(_02400__PTR39), .A2(_02379__PTR4), .ZN(_02401__PTR39) );
  AND2_X1 U12525 ( .A1(_02400__PTR40), .A2(_02379__PTR4), .ZN(_02401__PTR40) );
  AND2_X1 U12526 ( .A1(_02400__PTR41), .A2(_02379__PTR4), .ZN(_02401__PTR41) );
  AND2_X1 U12527 ( .A1(_02400__PTR42), .A2(_02379__PTR4), .ZN(_02401__PTR42) );
  AND2_X1 U12528 ( .A1(_02400__PTR43), .A2(_02379__PTR4), .ZN(_02401__PTR43) );
  AND2_X1 U12529 ( .A1(_02400__PTR44), .A2(_02379__PTR4), .ZN(_02401__PTR44) );
  AND2_X1 U12530 ( .A1(_02400__PTR45), .A2(_02379__PTR4), .ZN(_02401__PTR45) );
  AND2_X1 U12531 ( .A1(_02400__PTR46), .A2(_02379__PTR4), .ZN(_02401__PTR46) );
  AND2_X1 U12532 ( .A1(_02400__PTR47), .A2(_02379__PTR4), .ZN(_02401__PTR47) );
  AND2_X1 U12533 ( .A1(P2_P1_uWord_PTR0), .A2(_02398__PTR0), .ZN(_02397__PTR0) );
  AND2_X1 U12534 ( .A1(P2_P1_uWord_PTR1), .A2(_02398__PTR0), .ZN(_02397__PTR1) );
  AND2_X1 U12535 ( .A1(P2_P1_uWord_PTR2), .A2(_02398__PTR0), .ZN(_02397__PTR2) );
  AND2_X1 U12536 ( .A1(P2_P1_uWord_PTR3), .A2(_02398__PTR0), .ZN(_02397__PTR3) );
  AND2_X1 U12537 ( .A1(P2_P1_uWord_PTR4), .A2(_02398__PTR0), .ZN(_02397__PTR4) );
  AND2_X1 U12538 ( .A1(P2_P1_uWord_PTR5), .A2(_02398__PTR0), .ZN(_02397__PTR5) );
  AND2_X1 U12539 ( .A1(P2_P1_uWord_PTR6), .A2(_02398__PTR0), .ZN(_02397__PTR6) );
  AND2_X1 U12540 ( .A1(P2_P1_uWord_PTR7), .A2(_02398__PTR0), .ZN(_02397__PTR7) );
  AND2_X1 U12541 ( .A1(P2_P1_uWord_PTR8), .A2(_02398__PTR0), .ZN(_02397__PTR8) );
  AND2_X1 U12542 ( .A1(P2_P1_uWord_PTR9), .A2(_02398__PTR0), .ZN(_02397__PTR9) );
  AND2_X1 U12543 ( .A1(P2_P1_uWord_PTR10), .A2(_02398__PTR0), .ZN(_02397__PTR10) );
  AND2_X1 U12544 ( .A1(P2_P1_uWord_PTR11), .A2(_02398__PTR0), .ZN(_02397__PTR11) );
  AND2_X1 U12545 ( .A1(P2_P1_uWord_PTR12), .A2(_02398__PTR0), .ZN(_02397__PTR12) );
  AND2_X1 U12546 ( .A1(P2_P1_uWord_PTR13), .A2(_02398__PTR0), .ZN(_02397__PTR13) );
  AND2_X1 U12547 ( .A1(P2_P1_uWord_PTR14), .A2(_02398__PTR0), .ZN(_02397__PTR14) );
  AND2_X1 U12548 ( .A1(_02396__PTR15), .A2(_02156__PTR2), .ZN(_02397__PTR15) );
  AND2_X1 U12549 ( .A1(_02396__PTR16), .A2(_02156__PTR2), .ZN(_02397__PTR16) );
  AND2_X1 U12550 ( .A1(_02396__PTR17), .A2(_02156__PTR2), .ZN(_02397__PTR17) );
  AND2_X1 U12551 ( .A1(_02396__PTR18), .A2(_02156__PTR2), .ZN(_02397__PTR18) );
  AND2_X1 U12552 ( .A1(_02396__PTR19), .A2(_02156__PTR2), .ZN(_02397__PTR19) );
  AND2_X1 U12553 ( .A1(_02396__PTR20), .A2(_02156__PTR2), .ZN(_02397__PTR20) );
  AND2_X1 U12554 ( .A1(_02396__PTR21), .A2(_02156__PTR2), .ZN(_02397__PTR21) );
  AND2_X1 U12555 ( .A1(_02396__PTR22), .A2(_02156__PTR2), .ZN(_02397__PTR22) );
  AND2_X1 U12556 ( .A1(_02396__PTR23), .A2(_02156__PTR2), .ZN(_02397__PTR23) );
  AND2_X1 U12557 ( .A1(_02396__PTR24), .A2(_02156__PTR2), .ZN(_02397__PTR24) );
  AND2_X1 U12558 ( .A1(_02396__PTR25), .A2(_02156__PTR2), .ZN(_02397__PTR25) );
  AND2_X1 U12559 ( .A1(_02396__PTR26), .A2(_02156__PTR2), .ZN(_02397__PTR26) );
  AND2_X1 U12560 ( .A1(_02396__PTR27), .A2(_02156__PTR2), .ZN(_02397__PTR27) );
  AND2_X1 U12561 ( .A1(_02396__PTR28), .A2(_02156__PTR2), .ZN(_02397__PTR28) );
  AND2_X1 U12562 ( .A1(_02396__PTR29), .A2(_02156__PTR2), .ZN(_02397__PTR29) );
  AND2_X1 U12563 ( .A1(_02396__PTR30), .A2(_02379__PTR4), .ZN(_02397__PTR30) );
  AND2_X1 U12564 ( .A1(_02396__PTR31), .A2(_02379__PTR4), .ZN(_02397__PTR31) );
  AND2_X1 U12565 ( .A1(_02396__PTR32), .A2(_02379__PTR4), .ZN(_02397__PTR32) );
  AND2_X1 U12566 ( .A1(_02396__PTR33), .A2(_02379__PTR4), .ZN(_02397__PTR33) );
  AND2_X1 U12567 ( .A1(_02396__PTR34), .A2(_02379__PTR4), .ZN(_02397__PTR34) );
  AND2_X1 U12568 ( .A1(_02396__PTR35), .A2(_02379__PTR4), .ZN(_02397__PTR35) );
  AND2_X1 U12569 ( .A1(_02396__PTR36), .A2(_02379__PTR4), .ZN(_02397__PTR36) );
  AND2_X1 U12570 ( .A1(_02396__PTR37), .A2(_02379__PTR4), .ZN(_02397__PTR37) );
  AND2_X1 U12571 ( .A1(_02396__PTR38), .A2(_02379__PTR4), .ZN(_02397__PTR38) );
  AND2_X1 U12572 ( .A1(_02396__PTR39), .A2(_02379__PTR4), .ZN(_02397__PTR39) );
  AND2_X1 U12573 ( .A1(_02396__PTR40), .A2(_02379__PTR4), .ZN(_02397__PTR40) );
  AND2_X1 U12574 ( .A1(_02396__PTR41), .A2(_02379__PTR4), .ZN(_02397__PTR41) );
  AND2_X1 U12575 ( .A1(_02396__PTR42), .A2(_02379__PTR4), .ZN(_02397__PTR42) );
  AND2_X1 U12576 ( .A1(_02396__PTR43), .A2(_02379__PTR4), .ZN(_02397__PTR43) );
  AND2_X1 U12577 ( .A1(_02396__PTR44), .A2(_02379__PTR4), .ZN(_02397__PTR44) );
  AND2_X1 U12578 ( .A1(P2_EBX_PTR0), .A2(_02391__PTR0), .ZN(_02390__PTR0) );
  AND2_X1 U12579 ( .A1(P2_EBX_PTR1), .A2(_02391__PTR0), .ZN(_02390__PTR1) );
  AND2_X1 U12580 ( .A1(P2_EBX_PTR2), .A2(_02391__PTR0), .ZN(_02390__PTR2) );
  AND2_X1 U12581 ( .A1(P2_EBX_PTR3), .A2(_02391__PTR0), .ZN(_02390__PTR3) );
  AND2_X1 U12582 ( .A1(P2_EBX_PTR4), .A2(_02391__PTR0), .ZN(_02390__PTR4) );
  AND2_X1 U12583 ( .A1(P2_EBX_PTR5), .A2(_02391__PTR0), .ZN(_02390__PTR5) );
  AND2_X1 U12584 ( .A1(P2_EBX_PTR6), .A2(_02391__PTR0), .ZN(_02390__PTR6) );
  AND2_X1 U12585 ( .A1(P2_EBX_PTR7), .A2(_02391__PTR0), .ZN(_02390__PTR7) );
  AND2_X1 U12586 ( .A1(P2_EBX_PTR8), .A2(_02391__PTR0), .ZN(_02390__PTR8) );
  AND2_X1 U12587 ( .A1(P2_EBX_PTR9), .A2(_02391__PTR0), .ZN(_02390__PTR9) );
  AND2_X1 U12588 ( .A1(P2_EBX_PTR10), .A2(_02391__PTR0), .ZN(_02390__PTR10) );
  AND2_X1 U12589 ( .A1(P2_EBX_PTR11), .A2(_02391__PTR0), .ZN(_02390__PTR11) );
  AND2_X1 U12590 ( .A1(P2_EBX_PTR12), .A2(_02391__PTR0), .ZN(_02390__PTR12) );
  AND2_X1 U12591 ( .A1(P2_EBX_PTR13), .A2(_02391__PTR0), .ZN(_02390__PTR13) );
  AND2_X1 U12592 ( .A1(P2_EBX_PTR14), .A2(_02391__PTR0), .ZN(_02390__PTR14) );
  AND2_X1 U12593 ( .A1(P2_EBX_PTR15), .A2(_02391__PTR0), .ZN(_02390__PTR15) );
  AND2_X1 U12594 ( .A1(P2_EBX_PTR16), .A2(_02391__PTR0), .ZN(_02390__PTR16) );
  AND2_X1 U12595 ( .A1(P2_EBX_PTR17), .A2(_02391__PTR0), .ZN(_02390__PTR17) );
  AND2_X1 U12596 ( .A1(P2_EBX_PTR18), .A2(_02391__PTR0), .ZN(_02390__PTR18) );
  AND2_X1 U12597 ( .A1(P2_EBX_PTR19), .A2(_02391__PTR0), .ZN(_02390__PTR19) );
  AND2_X1 U12598 ( .A1(P2_EBX_PTR20), .A2(_02391__PTR0), .ZN(_02390__PTR20) );
  AND2_X1 U12599 ( .A1(P2_EBX_PTR21), .A2(_02391__PTR0), .ZN(_02390__PTR21) );
  AND2_X1 U12600 ( .A1(P2_EBX_PTR22), .A2(_02391__PTR0), .ZN(_02390__PTR22) );
  AND2_X1 U12601 ( .A1(P2_EBX_PTR23), .A2(_02391__PTR0), .ZN(_02390__PTR23) );
  AND2_X1 U12602 ( .A1(P2_EBX_PTR24), .A2(_02391__PTR0), .ZN(_02390__PTR24) );
  AND2_X1 U12603 ( .A1(P2_EBX_PTR25), .A2(_02391__PTR0), .ZN(_02390__PTR25) );
  AND2_X1 U12604 ( .A1(P2_EBX_PTR26), .A2(_02391__PTR0), .ZN(_02390__PTR26) );
  AND2_X1 U12605 ( .A1(P2_EBX_PTR27), .A2(_02391__PTR0), .ZN(_02390__PTR27) );
  AND2_X1 U12606 ( .A1(P2_EBX_PTR28), .A2(_02391__PTR0), .ZN(_02390__PTR28) );
  AND2_X1 U12607 ( .A1(P2_EBX_PTR29), .A2(_02391__PTR0), .ZN(_02390__PTR29) );
  AND2_X1 U12608 ( .A1(P2_EBX_PTR30), .A2(_02391__PTR0), .ZN(_02390__PTR30) );
  AND2_X1 U12609 ( .A1(P2_EBX_PTR31), .A2(_02391__PTR0), .ZN(_02390__PTR31) );
  AND2_X1 U12610 ( .A1(_02389__PTR32), .A2(_02391__PTR1), .ZN(_02390__PTR32) );
  AND2_X1 U12611 ( .A1(_02389__PTR33), .A2(_02391__PTR1), .ZN(_02390__PTR33) );
  AND2_X1 U12612 ( .A1(_02389__PTR34), .A2(_02391__PTR1), .ZN(_02390__PTR34) );
  AND2_X1 U12613 ( .A1(_02389__PTR35), .A2(_02391__PTR1), .ZN(_02390__PTR35) );
  AND2_X1 U12614 ( .A1(_02389__PTR36), .A2(_02391__PTR1), .ZN(_02390__PTR36) );
  AND2_X1 U12615 ( .A1(_02389__PTR37), .A2(_02391__PTR1), .ZN(_02390__PTR37) );
  AND2_X1 U12616 ( .A1(_02389__PTR38), .A2(_02391__PTR1), .ZN(_02390__PTR38) );
  AND2_X1 U12617 ( .A1(_02389__PTR39), .A2(_02391__PTR1), .ZN(_02390__PTR39) );
  AND2_X1 U12618 ( .A1(_02389__PTR40), .A2(_02391__PTR1), .ZN(_02390__PTR40) );
  AND2_X1 U12619 ( .A1(_02389__PTR41), .A2(_02391__PTR1), .ZN(_02390__PTR41) );
  AND2_X1 U12620 ( .A1(_02389__PTR42), .A2(_02391__PTR1), .ZN(_02390__PTR42) );
  AND2_X1 U12621 ( .A1(_02389__PTR43), .A2(_02391__PTR1), .ZN(_02390__PTR43) );
  AND2_X1 U12622 ( .A1(_02389__PTR44), .A2(_02391__PTR1), .ZN(_02390__PTR44) );
  AND2_X1 U12623 ( .A1(_02389__PTR45), .A2(_02391__PTR1), .ZN(_02390__PTR45) );
  AND2_X1 U12624 ( .A1(_02389__PTR46), .A2(_02391__PTR1), .ZN(_02390__PTR46) );
  AND2_X1 U12625 ( .A1(_02389__PTR47), .A2(_02391__PTR1), .ZN(_02390__PTR47) );
  AND2_X1 U12626 ( .A1(_02389__PTR48), .A2(_02391__PTR1), .ZN(_02390__PTR48) );
  AND2_X1 U12627 ( .A1(_02389__PTR49), .A2(_02391__PTR1), .ZN(_02390__PTR49) );
  AND2_X1 U12628 ( .A1(_02389__PTR50), .A2(_02391__PTR1), .ZN(_02390__PTR50) );
  AND2_X1 U12629 ( .A1(_02389__PTR51), .A2(_02391__PTR1), .ZN(_02390__PTR51) );
  AND2_X1 U12630 ( .A1(_02389__PTR52), .A2(_02391__PTR1), .ZN(_02390__PTR52) );
  AND2_X1 U12631 ( .A1(_02389__PTR53), .A2(_02391__PTR1), .ZN(_02390__PTR53) );
  AND2_X1 U12632 ( .A1(_02389__PTR54), .A2(_02391__PTR1), .ZN(_02390__PTR54) );
  AND2_X1 U12633 ( .A1(_02389__PTR55), .A2(_02391__PTR1), .ZN(_02390__PTR55) );
  AND2_X1 U12634 ( .A1(_02389__PTR56), .A2(_02391__PTR1), .ZN(_02390__PTR56) );
  AND2_X1 U12635 ( .A1(_02389__PTR57), .A2(_02391__PTR1), .ZN(_02390__PTR57) );
  AND2_X1 U12636 ( .A1(_02389__PTR58), .A2(_02391__PTR1), .ZN(_02390__PTR58) );
  AND2_X1 U12637 ( .A1(_02389__PTR59), .A2(_02391__PTR1), .ZN(_02390__PTR59) );
  AND2_X1 U12638 ( .A1(_02389__PTR60), .A2(_02391__PTR1), .ZN(_02390__PTR60) );
  AND2_X1 U12639 ( .A1(_02389__PTR61), .A2(_02391__PTR1), .ZN(_02390__PTR61) );
  AND2_X1 U12640 ( .A1(_02389__PTR62), .A2(_02391__PTR1), .ZN(_02390__PTR62) );
  AND2_X1 U12641 ( .A1(_02389__PTR63), .A2(_02391__PTR1), .ZN(_02390__PTR63) );
  AND2_X1 U12642 ( .A1(_02389__PTR64), .A2(_02391__PTR2), .ZN(_02390__PTR64) );
  AND2_X1 U12643 ( .A1(_02389__PTR65), .A2(_02391__PTR2), .ZN(_02390__PTR65) );
  AND2_X1 U12644 ( .A1(_02389__PTR66), .A2(_02391__PTR2), .ZN(_02390__PTR66) );
  AND2_X1 U12645 ( .A1(_02389__PTR67), .A2(_02391__PTR2), .ZN(_02390__PTR67) );
  AND2_X1 U12646 ( .A1(_02389__PTR68), .A2(_02391__PTR2), .ZN(_02390__PTR68) );
  AND2_X1 U12647 ( .A1(_02389__PTR69), .A2(_02391__PTR2), .ZN(_02390__PTR69) );
  AND2_X1 U12648 ( .A1(_02389__PTR70), .A2(_02391__PTR2), .ZN(_02390__PTR70) );
  AND2_X1 U12649 ( .A1(_02389__PTR71), .A2(_02391__PTR2), .ZN(_02390__PTR71) );
  AND2_X1 U12650 ( .A1(_02389__PTR72), .A2(_02391__PTR2), .ZN(_02390__PTR72) );
  AND2_X1 U12651 ( .A1(_02389__PTR73), .A2(_02391__PTR2), .ZN(_02390__PTR73) );
  AND2_X1 U12652 ( .A1(_02389__PTR74), .A2(_02391__PTR2), .ZN(_02390__PTR74) );
  AND2_X1 U12653 ( .A1(_02389__PTR75), .A2(_02391__PTR2), .ZN(_02390__PTR75) );
  AND2_X1 U12654 ( .A1(_02389__PTR76), .A2(_02391__PTR2), .ZN(_02390__PTR76) );
  AND2_X1 U12655 ( .A1(_02389__PTR77), .A2(_02391__PTR2), .ZN(_02390__PTR77) );
  AND2_X1 U12656 ( .A1(_02389__PTR78), .A2(_02391__PTR2), .ZN(_02390__PTR78) );
  AND2_X1 U12657 ( .A1(_02389__PTR79), .A2(_02391__PTR2), .ZN(_02390__PTR79) );
  AND2_X1 U12658 ( .A1(_02389__PTR80), .A2(_02391__PTR2), .ZN(_02390__PTR80) );
  AND2_X1 U12659 ( .A1(_02389__PTR81), .A2(_02391__PTR2), .ZN(_02390__PTR81) );
  AND2_X1 U12660 ( .A1(_02389__PTR82), .A2(_02391__PTR2), .ZN(_02390__PTR82) );
  AND2_X1 U12661 ( .A1(_02389__PTR83), .A2(_02391__PTR2), .ZN(_02390__PTR83) );
  AND2_X1 U12662 ( .A1(_02389__PTR84), .A2(_02391__PTR2), .ZN(_02390__PTR84) );
  AND2_X1 U12663 ( .A1(_02389__PTR85), .A2(_02391__PTR2), .ZN(_02390__PTR85) );
  AND2_X1 U12664 ( .A1(_02389__PTR86), .A2(_02391__PTR2), .ZN(_02390__PTR86) );
  AND2_X1 U12665 ( .A1(_02389__PTR87), .A2(_02391__PTR2), .ZN(_02390__PTR87) );
  AND2_X1 U12666 ( .A1(_02389__PTR88), .A2(_02391__PTR2), .ZN(_02390__PTR88) );
  AND2_X1 U12667 ( .A1(_02389__PTR89), .A2(_02391__PTR2), .ZN(_02390__PTR89) );
  AND2_X1 U12668 ( .A1(_02389__PTR90), .A2(_02391__PTR2), .ZN(_02390__PTR90) );
  AND2_X1 U12669 ( .A1(_02389__PTR91), .A2(_02391__PTR2), .ZN(_02390__PTR91) );
  AND2_X1 U12670 ( .A1(_02389__PTR92), .A2(_02391__PTR2), .ZN(_02390__PTR92) );
  AND2_X1 U12671 ( .A1(_02389__PTR93), .A2(_02391__PTR2), .ZN(_02390__PTR93) );
  AND2_X1 U12672 ( .A1(_02389__PTR94), .A2(_02391__PTR2), .ZN(_02390__PTR94) );
  AND2_X1 U12673 ( .A1(_02389__PTR95), .A2(_02391__PTR2), .ZN(_02390__PTR95) );
  AND2_X1 U12674 ( .A1(P2_EAX_PTR0), .A2(_02387__PTR0), .ZN(_02386__PTR0) );
  AND2_X1 U12675 ( .A1(P2_EAX_PTR1), .A2(_02387__PTR0), .ZN(_02386__PTR1) );
  AND2_X1 U12676 ( .A1(P2_EAX_PTR2), .A2(_02387__PTR0), .ZN(_02386__PTR2) );
  AND2_X1 U12677 ( .A1(P2_EAX_PTR3), .A2(_02387__PTR0), .ZN(_02386__PTR3) );
  AND2_X1 U12678 ( .A1(P2_EAX_PTR4), .A2(_02387__PTR0), .ZN(_02386__PTR4) );
  AND2_X1 U12679 ( .A1(P2_EAX_PTR5), .A2(_02387__PTR0), .ZN(_02386__PTR5) );
  AND2_X1 U12680 ( .A1(P2_EAX_PTR6), .A2(_02387__PTR0), .ZN(_02386__PTR6) );
  AND2_X1 U12681 ( .A1(P2_EAX_PTR7), .A2(_02387__PTR0), .ZN(_02386__PTR7) );
  AND2_X1 U12682 ( .A1(P2_EAX_PTR8), .A2(_02387__PTR0), .ZN(_02386__PTR8) );
  AND2_X1 U12683 ( .A1(P2_EAX_PTR9), .A2(_02387__PTR0), .ZN(_02386__PTR9) );
  AND2_X1 U12684 ( .A1(P2_EAX_PTR10), .A2(_02387__PTR0), .ZN(_02386__PTR10) );
  AND2_X1 U12685 ( .A1(P2_EAX_PTR11), .A2(_02387__PTR0), .ZN(_02386__PTR11) );
  AND2_X1 U12686 ( .A1(P2_EAX_PTR12), .A2(_02387__PTR0), .ZN(_02386__PTR12) );
  AND2_X1 U12687 ( .A1(P2_EAX_PTR13), .A2(_02387__PTR0), .ZN(_02386__PTR13) );
  AND2_X1 U12688 ( .A1(P2_EAX_PTR14), .A2(_02387__PTR0), .ZN(_02386__PTR14) );
  AND2_X1 U12689 ( .A1(P2_EAX_PTR15), .A2(_02387__PTR0), .ZN(_02386__PTR15) );
  AND2_X1 U12690 ( .A1(P2_EAX_PTR16), .A2(_02387__PTR0), .ZN(_02386__PTR16) );
  AND2_X1 U12691 ( .A1(P2_EAX_PTR17), .A2(_02387__PTR0), .ZN(_02386__PTR17) );
  AND2_X1 U12692 ( .A1(P2_EAX_PTR18), .A2(_02387__PTR0), .ZN(_02386__PTR18) );
  AND2_X1 U12693 ( .A1(P2_EAX_PTR19), .A2(_02387__PTR0), .ZN(_02386__PTR19) );
  AND2_X1 U12694 ( .A1(P2_EAX_PTR20), .A2(_02387__PTR0), .ZN(_02386__PTR20) );
  AND2_X1 U12695 ( .A1(P2_EAX_PTR21), .A2(_02387__PTR0), .ZN(_02386__PTR21) );
  AND2_X1 U12696 ( .A1(P2_EAX_PTR22), .A2(_02387__PTR0), .ZN(_02386__PTR22) );
  AND2_X1 U12697 ( .A1(P2_EAX_PTR23), .A2(_02387__PTR0), .ZN(_02386__PTR23) );
  AND2_X1 U12698 ( .A1(P2_EAX_PTR24), .A2(_02387__PTR0), .ZN(_02386__PTR24) );
  AND2_X1 U12699 ( .A1(P2_EAX_PTR25), .A2(_02387__PTR0), .ZN(_02386__PTR25) );
  AND2_X1 U12700 ( .A1(P2_EAX_PTR26), .A2(_02387__PTR0), .ZN(_02386__PTR26) );
  AND2_X1 U12701 ( .A1(P2_EAX_PTR27), .A2(_02387__PTR0), .ZN(_02386__PTR27) );
  AND2_X1 U12702 ( .A1(P2_EAX_PTR28), .A2(_02387__PTR0), .ZN(_02386__PTR28) );
  AND2_X1 U12703 ( .A1(P2_EAX_PTR29), .A2(_02387__PTR0), .ZN(_02386__PTR29) );
  AND2_X1 U12704 ( .A1(P2_EAX_PTR30), .A2(_02387__PTR0), .ZN(_02386__PTR30) );
  AND2_X1 U12705 ( .A1(P2_EAX_PTR31), .A2(_02387__PTR0), .ZN(_02386__PTR31) );
  AND2_X1 U12706 ( .A1(_02385__PTR32), .A2(_02387__PTR1), .ZN(_02386__PTR32) );
  AND2_X1 U12707 ( .A1(_02385__PTR33), .A2(_02387__PTR1), .ZN(_02386__PTR33) );
  AND2_X1 U12708 ( .A1(_02385__PTR34), .A2(_02387__PTR1), .ZN(_02386__PTR34) );
  AND2_X1 U12709 ( .A1(_02385__PTR35), .A2(_02387__PTR1), .ZN(_02386__PTR35) );
  AND2_X1 U12710 ( .A1(_02385__PTR36), .A2(_02387__PTR1), .ZN(_02386__PTR36) );
  AND2_X1 U12711 ( .A1(_02385__PTR37), .A2(_02387__PTR1), .ZN(_02386__PTR37) );
  AND2_X1 U12712 ( .A1(_02385__PTR38), .A2(_02387__PTR1), .ZN(_02386__PTR38) );
  AND2_X1 U12713 ( .A1(_02385__PTR39), .A2(_02387__PTR1), .ZN(_02386__PTR39) );
  AND2_X1 U12714 ( .A1(_02385__PTR40), .A2(_02387__PTR1), .ZN(_02386__PTR40) );
  AND2_X1 U12715 ( .A1(_02385__PTR41), .A2(_02387__PTR1), .ZN(_02386__PTR41) );
  AND2_X1 U12716 ( .A1(_02385__PTR42), .A2(_02387__PTR1), .ZN(_02386__PTR42) );
  AND2_X1 U12717 ( .A1(_02385__PTR43), .A2(_02387__PTR1), .ZN(_02386__PTR43) );
  AND2_X1 U12718 ( .A1(_02385__PTR44), .A2(_02387__PTR1), .ZN(_02386__PTR44) );
  AND2_X1 U12719 ( .A1(_02385__PTR45), .A2(_02387__PTR1), .ZN(_02386__PTR45) );
  AND2_X1 U12720 ( .A1(_02385__PTR46), .A2(_02387__PTR1), .ZN(_02386__PTR46) );
  AND2_X1 U12721 ( .A1(_02385__PTR47), .A2(_02387__PTR1), .ZN(_02386__PTR47) );
  AND2_X1 U12722 ( .A1(_02385__PTR48), .A2(_02387__PTR1), .ZN(_02386__PTR48) );
  AND2_X1 U12723 ( .A1(_02385__PTR49), .A2(_02387__PTR1), .ZN(_02386__PTR49) );
  AND2_X1 U12724 ( .A1(_02385__PTR50), .A2(_02387__PTR1), .ZN(_02386__PTR50) );
  AND2_X1 U12725 ( .A1(_02385__PTR51), .A2(_02387__PTR1), .ZN(_02386__PTR51) );
  AND2_X1 U12726 ( .A1(_02385__PTR52), .A2(_02387__PTR1), .ZN(_02386__PTR52) );
  AND2_X1 U12727 ( .A1(_02385__PTR53), .A2(_02387__PTR1), .ZN(_02386__PTR53) );
  AND2_X1 U12728 ( .A1(_02385__PTR54), .A2(_02387__PTR1), .ZN(_02386__PTR54) );
  AND2_X1 U12729 ( .A1(_02385__PTR55), .A2(_02387__PTR1), .ZN(_02386__PTR55) );
  AND2_X1 U12730 ( .A1(_02385__PTR56), .A2(_02387__PTR1), .ZN(_02386__PTR56) );
  AND2_X1 U12731 ( .A1(_02385__PTR57), .A2(_02387__PTR1), .ZN(_02386__PTR57) );
  AND2_X1 U12732 ( .A1(_02385__PTR58), .A2(_02387__PTR1), .ZN(_02386__PTR58) );
  AND2_X1 U12733 ( .A1(_02385__PTR59), .A2(_02387__PTR1), .ZN(_02386__PTR59) );
  AND2_X1 U12734 ( .A1(_02385__PTR60), .A2(_02387__PTR1), .ZN(_02386__PTR60) );
  AND2_X1 U12735 ( .A1(_02385__PTR61), .A2(_02387__PTR1), .ZN(_02386__PTR61) );
  AND2_X1 U12736 ( .A1(_02385__PTR62), .A2(_02387__PTR1), .ZN(_02386__PTR62) );
  AND2_X1 U12737 ( .A1(_02385__PTR63), .A2(_02387__PTR1), .ZN(_02386__PTR63) );
  AND2_X1 U12738 ( .A1(_02385__PTR96), .A2(_02379__PTR3), .ZN(_02386__PTR64) );
  AND2_X1 U12739 ( .A1(_02385__PTR97), .A2(_02379__PTR3), .ZN(_02386__PTR65) );
  AND2_X1 U12740 ( .A1(_02385__PTR98), .A2(_02379__PTR3), .ZN(_02386__PTR66) );
  AND2_X1 U12741 ( .A1(_02385__PTR99), .A2(_02379__PTR3), .ZN(_02386__PTR67) );
  AND2_X1 U12742 ( .A1(_02385__PTR100), .A2(_02379__PTR3), .ZN(_02386__PTR68) );
  AND2_X1 U12743 ( .A1(_02385__PTR101), .A2(_02379__PTR3), .ZN(_02386__PTR69) );
  AND2_X1 U12744 ( .A1(_02385__PTR102), .A2(_02379__PTR3), .ZN(_02386__PTR70) );
  AND2_X1 U12745 ( .A1(_02385__PTR103), .A2(_02379__PTR3), .ZN(_02386__PTR71) );
  AND2_X1 U12746 ( .A1(_02385__PTR104), .A2(_02379__PTR3), .ZN(_02386__PTR72) );
  AND2_X1 U12747 ( .A1(_02385__PTR105), .A2(_02379__PTR3), .ZN(_02386__PTR73) );
  AND2_X1 U12748 ( .A1(_02385__PTR106), .A2(_02379__PTR3), .ZN(_02386__PTR74) );
  AND2_X1 U12749 ( .A1(_02385__PTR107), .A2(_02379__PTR3), .ZN(_02386__PTR75) );
  AND2_X1 U12750 ( .A1(_02385__PTR108), .A2(_02379__PTR3), .ZN(_02386__PTR76) );
  AND2_X1 U12751 ( .A1(_02385__PTR109), .A2(_02379__PTR3), .ZN(_02386__PTR77) );
  AND2_X1 U12752 ( .A1(_02385__PTR110), .A2(_02379__PTR3), .ZN(_02386__PTR78) );
  AND2_X1 U12753 ( .A1(_02385__PTR111), .A2(_02379__PTR3), .ZN(_02386__PTR79) );
  AND2_X1 U12754 ( .A1(_02385__PTR80), .A2(_02379__PTR3), .ZN(_02386__PTR80) );
  AND2_X1 U12755 ( .A1(_02385__PTR81), .A2(_02379__PTR3), .ZN(_02386__PTR81) );
  AND2_X1 U12756 ( .A1(_02385__PTR82), .A2(_02379__PTR3), .ZN(_02386__PTR82) );
  AND2_X1 U12757 ( .A1(_02385__PTR83), .A2(_02379__PTR3), .ZN(_02386__PTR83) );
  AND2_X1 U12758 ( .A1(_02385__PTR84), .A2(_02379__PTR3), .ZN(_02386__PTR84) );
  AND2_X1 U12759 ( .A1(_02385__PTR85), .A2(_02379__PTR3), .ZN(_02386__PTR85) );
  AND2_X1 U12760 ( .A1(_02385__PTR86), .A2(_02379__PTR3), .ZN(_02386__PTR86) );
  AND2_X1 U12761 ( .A1(_02385__PTR87), .A2(_02379__PTR3), .ZN(_02386__PTR87) );
  AND2_X1 U12762 ( .A1(_02385__PTR88), .A2(_02379__PTR3), .ZN(_02386__PTR88) );
  AND2_X1 U12763 ( .A1(_02385__PTR89), .A2(_02379__PTR3), .ZN(_02386__PTR89) );
  AND2_X1 U12764 ( .A1(_02385__PTR90), .A2(_02379__PTR3), .ZN(_02386__PTR90) );
  AND2_X1 U12765 ( .A1(_02385__PTR91), .A2(_02379__PTR3), .ZN(_02386__PTR91) );
  AND2_X1 U12766 ( .A1(_02385__PTR92), .A2(_02379__PTR3), .ZN(_02386__PTR92) );
  AND2_X1 U12767 ( .A1(_02385__PTR93), .A2(_02379__PTR3), .ZN(_02386__PTR93) );
  AND2_X1 U12768 ( .A1(_02385__PTR94), .A2(_02379__PTR3), .ZN(_02386__PTR94) );
  AND2_X1 U12769 ( .A1(_02385__PTR95), .A2(_02379__PTR3), .ZN(_02386__PTR95) );
  AND2_X1 U12770 ( .A1(_02385__PTR96), .A2(_02379__PTR4), .ZN(_02386__PTR96) );
  AND2_X1 U12771 ( .A1(_02385__PTR97), .A2(_02379__PTR4), .ZN(_02386__PTR97) );
  AND2_X1 U12772 ( .A1(_02385__PTR98), .A2(_02379__PTR4), .ZN(_02386__PTR98) );
  AND2_X1 U12773 ( .A1(_02385__PTR99), .A2(_02379__PTR4), .ZN(_02386__PTR99) );
  AND2_X1 U12774 ( .A1(_02385__PTR100), .A2(_02379__PTR4), .ZN(_02386__PTR100) );
  AND2_X1 U12775 ( .A1(_02385__PTR101), .A2(_02379__PTR4), .ZN(_02386__PTR101) );
  AND2_X1 U12776 ( .A1(_02385__PTR102), .A2(_02379__PTR4), .ZN(_02386__PTR102) );
  AND2_X1 U12777 ( .A1(_02385__PTR103), .A2(_02379__PTR4), .ZN(_02386__PTR103) );
  AND2_X1 U12778 ( .A1(_02385__PTR104), .A2(_02379__PTR4), .ZN(_02386__PTR104) );
  AND2_X1 U12779 ( .A1(_02385__PTR105), .A2(_02379__PTR4), .ZN(_02386__PTR105) );
  AND2_X1 U12780 ( .A1(_02385__PTR106), .A2(_02379__PTR4), .ZN(_02386__PTR106) );
  AND2_X1 U12781 ( .A1(_02385__PTR107), .A2(_02379__PTR4), .ZN(_02386__PTR107) );
  AND2_X1 U12782 ( .A1(_02385__PTR108), .A2(_02379__PTR4), .ZN(_02386__PTR108) );
  AND2_X1 U12783 ( .A1(_02385__PTR109), .A2(_02379__PTR4), .ZN(_02386__PTR109) );
  AND2_X1 U12784 ( .A1(_02385__PTR110), .A2(_02379__PTR4), .ZN(_02386__PTR110) );
  AND2_X1 U12785 ( .A1(_02385__PTR111), .A2(_02379__PTR4), .ZN(_02386__PTR111) );
  AND2_X1 U12786 ( .A1(_02385__PTR112), .A2(_02379__PTR4), .ZN(_02386__PTR112) );
  AND2_X1 U12787 ( .A1(_02385__PTR113), .A2(_02379__PTR4), .ZN(_02386__PTR113) );
  AND2_X1 U12788 ( .A1(_02385__PTR114), .A2(_02379__PTR4), .ZN(_02386__PTR114) );
  AND2_X1 U12789 ( .A1(_02385__PTR115), .A2(_02379__PTR4), .ZN(_02386__PTR115) );
  AND2_X1 U12790 ( .A1(_02385__PTR116), .A2(_02379__PTR4), .ZN(_02386__PTR116) );
  AND2_X1 U12791 ( .A1(_02385__PTR117), .A2(_02379__PTR4), .ZN(_02386__PTR117) );
  AND2_X1 U12792 ( .A1(_02385__PTR118), .A2(_02379__PTR4), .ZN(_02386__PTR118) );
  AND2_X1 U12793 ( .A1(_02385__PTR119), .A2(_02379__PTR4), .ZN(_02386__PTR119) );
  AND2_X1 U12794 ( .A1(_02385__PTR120), .A2(_02379__PTR4), .ZN(_02386__PTR120) );
  AND2_X1 U12795 ( .A1(_02385__PTR121), .A2(_02379__PTR4), .ZN(_02386__PTR121) );
  AND2_X1 U12796 ( .A1(_02385__PTR122), .A2(_02379__PTR4), .ZN(_02386__PTR122) );
  AND2_X1 U12797 ( .A1(_02385__PTR123), .A2(_02379__PTR4), .ZN(_02386__PTR123) );
  AND2_X1 U12798 ( .A1(_02385__PTR124), .A2(_02379__PTR4), .ZN(_02386__PTR124) );
  AND2_X1 U12799 ( .A1(_02385__PTR125), .A2(_02379__PTR4), .ZN(_02386__PTR125) );
  AND2_X1 U12800 ( .A1(_02385__PTR126), .A2(_02379__PTR4), .ZN(_02386__PTR126) );
  AND2_X1 U12801 ( .A1(_02385__PTR127), .A2(_02379__PTR4), .ZN(_02386__PTR127) );
  AND2_X1 U12802 ( .A1(_02385__PTR128), .A2(_02387__PTR4), .ZN(_02386__PTR128) );
  AND2_X1 U12803 ( .A1(_02385__PTR129), .A2(_02387__PTR4), .ZN(_02386__PTR129) );
  AND2_X1 U12804 ( .A1(_02385__PTR130), .A2(_02387__PTR4), .ZN(_02386__PTR130) );
  AND2_X1 U12805 ( .A1(_02385__PTR131), .A2(_02387__PTR4), .ZN(_02386__PTR131) );
  AND2_X1 U12806 ( .A1(_02385__PTR132), .A2(_02387__PTR4), .ZN(_02386__PTR132) );
  AND2_X1 U12807 ( .A1(_02385__PTR133), .A2(_02387__PTR4), .ZN(_02386__PTR133) );
  AND2_X1 U12808 ( .A1(_02385__PTR134), .A2(_02387__PTR4), .ZN(_02386__PTR134) );
  AND2_X1 U12809 ( .A1(_02385__PTR135), .A2(_02387__PTR4), .ZN(_02386__PTR135) );
  AND2_X1 U12810 ( .A1(_02385__PTR136), .A2(_02387__PTR4), .ZN(_02386__PTR136) );
  AND2_X1 U12811 ( .A1(_02385__PTR137), .A2(_02387__PTR4), .ZN(_02386__PTR137) );
  AND2_X1 U12812 ( .A1(_02385__PTR138), .A2(_02387__PTR4), .ZN(_02386__PTR138) );
  AND2_X1 U12813 ( .A1(_02385__PTR139), .A2(_02387__PTR4), .ZN(_02386__PTR139) );
  AND2_X1 U12814 ( .A1(_02385__PTR140), .A2(_02387__PTR4), .ZN(_02386__PTR140) );
  AND2_X1 U12815 ( .A1(_02385__PTR141), .A2(_02387__PTR4), .ZN(_02386__PTR141) );
  AND2_X1 U12816 ( .A1(_02385__PTR142), .A2(_02387__PTR4), .ZN(_02386__PTR142) );
  AND2_X1 U12817 ( .A1(_02385__PTR143), .A2(_02387__PTR4), .ZN(_02386__PTR143) );
  AND2_X1 U12818 ( .A1(_02385__PTR144), .A2(_02387__PTR4), .ZN(_02386__PTR144) );
  AND2_X1 U12819 ( .A1(_02385__PTR145), .A2(_02387__PTR4), .ZN(_02386__PTR145) );
  AND2_X1 U12820 ( .A1(_02385__PTR146), .A2(_02387__PTR4), .ZN(_02386__PTR146) );
  AND2_X1 U12821 ( .A1(_02385__PTR147), .A2(_02387__PTR4), .ZN(_02386__PTR147) );
  AND2_X1 U12822 ( .A1(_02385__PTR148), .A2(_02387__PTR4), .ZN(_02386__PTR148) );
  AND2_X1 U12823 ( .A1(_02385__PTR149), .A2(_02387__PTR4), .ZN(_02386__PTR149) );
  AND2_X1 U12824 ( .A1(_02385__PTR150), .A2(_02387__PTR4), .ZN(_02386__PTR150) );
  AND2_X1 U12825 ( .A1(_02385__PTR151), .A2(_02387__PTR4), .ZN(_02386__PTR151) );
  AND2_X1 U12826 ( .A1(_02385__PTR152), .A2(_02387__PTR4), .ZN(_02386__PTR152) );
  AND2_X1 U12827 ( .A1(_02385__PTR153), .A2(_02387__PTR4), .ZN(_02386__PTR153) );
  AND2_X1 U12828 ( .A1(_02385__PTR154), .A2(_02387__PTR4), .ZN(_02386__PTR154) );
  AND2_X1 U12829 ( .A1(_02385__PTR155), .A2(_02387__PTR4), .ZN(_02386__PTR155) );
  AND2_X1 U12830 ( .A1(_02385__PTR156), .A2(_02387__PTR4), .ZN(_02386__PTR156) );
  AND2_X1 U12831 ( .A1(_02385__PTR157), .A2(_02387__PTR4), .ZN(_02386__PTR157) );
  AND2_X1 U12832 ( .A1(_02385__PTR158), .A2(_02387__PTR4), .ZN(_02386__PTR158) );
  AND2_X1 U12833 ( .A1(_02385__PTR159), .A2(_02387__PTR4), .ZN(_02386__PTR159) );
  AND2_X1 U12834 ( .A1(_02150__PTR0), .A2(_02148__PTR0), .ZN(_02151__PTR0) );
  AND2_X1 U12835 ( .A1(_02150__PTR1), .A2(_02148__PTR1), .ZN(_02151__PTR1) );
  AND2_X1 U12836 ( .A1(_02150__PTR2), .A2(_02152__PTR2), .ZN(_02151__PTR2) );
  AND2_X1 U12837 ( .A1(_02150__PTR3), .A2(_02148__PTR3), .ZN(_02151__PTR3) );
  AND2_X1 U12838 ( .A1(_02146__PTR0), .A2(_02148__PTR0), .ZN(_02147__PTR0) );
  AND2_X1 U12839 ( .A1(_02146__PTR1), .A2(_02148__PTR1), .ZN(_02147__PTR1) );
  AND2_X1 U12840 ( .A1(_02146__PTR2), .A2(_02148__PTR2), .ZN(_02147__PTR2) );
  AND2_X1 U12841 ( .A1(_02146__PTR3), .A2(_02148__PTR3), .ZN(_02147__PTR3) );
  AND2_X1 U12842 ( .A1(_02176__PTR3), .A2(_02375__PTR0), .ZN(_02378__PTR0) );
  AND2_X1 U12843 ( .A1(_02176__PTR4), .A2(_02375__PTR0), .ZN(_02378__PTR1) );
  AND2_X1 U12844 ( .A1(_02176__PTR5), .A2(_02375__PTR0), .ZN(_02378__PTR2) );
  AND2_X1 U12845 ( .A1(_02176__PTR6), .A2(_02375__PTR0), .ZN(_02378__PTR3) );
  AND2_X1 U12846 ( .A1(P2_P1_InstQueueRd_Addr_PTR0), .A2(_02375__PTR1), .ZN(_02378__PTR5) );
  AND2_X1 U12847 ( .A1(_02182__PTR4), .A2(_02375__PTR1), .ZN(_02378__PTR6) );
  AND2_X1 U12848 ( .A1(_02182__PTR5), .A2(_02375__PTR1), .ZN(_02378__PTR7) );
  AND2_X1 U12849 ( .A1(_02182__PTR6), .A2(_02375__PTR1), .ZN(_02378__PTR8) );
  AND2_X1 U12850 ( .A1(P2_P1_InstQueueRd_Addr_PTR0), .A2(_02148__PTR0), .ZN(_02378__PTR10) );
  AND2_X1 U12851 ( .A1(_02377__PTR11), .A2(_02148__PTR0), .ZN(_02378__PTR11) );
  AND2_X1 U12852 ( .A1(_02377__PTR12), .A2(_02148__PTR0), .ZN(_02378__PTR12) );
  AND2_X1 U12853 ( .A1(_02377__PTR13), .A2(_02148__PTR0), .ZN(_02378__PTR13) );
  AND2_X1 U12854 ( .A1(_02377__PTR14), .A2(_02148__PTR0), .ZN(_02378__PTR14) );
  AND2_X1 U12855 ( .A1(P2_P1_InstQueueRd_Addr_PTR0), .A2(_02379__PTR3), .ZN(_02378__PTR15) );
  AND2_X1 U12856 ( .A1(_02377__PTR21), .A2(_02379__PTR3), .ZN(_02378__PTR16) );
  AND2_X1 U12857 ( .A1(_02377__PTR22), .A2(_02379__PTR3), .ZN(_02378__PTR17) );
  AND2_X1 U12858 ( .A1(_02377__PTR23), .A2(_02379__PTR3), .ZN(_02378__PTR18) );
  AND2_X1 U12859 ( .A1(_02377__PTR19), .A2(_02379__PTR3), .ZN(_02378__PTR19) );
  AND2_X1 U12860 ( .A1(P2_P1_InstQueueRd_Addr_PTR0), .A2(_02379__PTR4), .ZN(_02378__PTR20) );
  AND2_X1 U12861 ( .A1(_02377__PTR21), .A2(_02379__PTR4), .ZN(_02378__PTR21) );
  AND2_X1 U12862 ( .A1(_02377__PTR22), .A2(_02379__PTR4), .ZN(_02378__PTR22) );
  AND2_X1 U12863 ( .A1(_02377__PTR23), .A2(_02379__PTR4), .ZN(_02378__PTR23) );
  AND2_X1 U12864 ( .A1(_02377__PTR24), .A2(_02379__PTR4), .ZN(_02378__PTR24) );
  AND2_X1 U12865 ( .A1(_02377__PTR25), .A2(_02375__PTR4), .ZN(_02378__PTR25) );
  AND2_X1 U12866 ( .A1(_02377__PTR26), .A2(_02375__PTR4), .ZN(_02378__PTR26) );
  AND2_X1 U12867 ( .A1(_02377__PTR27), .A2(_02375__PTR4), .ZN(_02378__PTR27) );
  AND2_X1 U12868 ( .A1(_02377__PTR28), .A2(_02375__PTR4), .ZN(_02378__PTR28) );
  AND2_X1 U12869 ( .A1(_02377__PTR29), .A2(_02375__PTR4), .ZN(_02378__PTR29) );
  AND2_X1 U12870 ( .A1(P2_P1_InstQueueRd_Addr_PTR0), .A2(_02379__PTR6), .ZN(_02378__PTR30) );
  AND2_X1 U12871 ( .A1(P2_P1_InstQueueRd_Addr_PTR1), .A2(_02379__PTR6), .ZN(_02378__PTR31) );
  AND2_X1 U12872 ( .A1(P2_P1_InstQueueRd_Addr_PTR2), .A2(_02379__PTR6), .ZN(_02378__PTR32) );
  AND2_X1 U12873 ( .A1(P2_P1_InstQueueRd_Addr_PTR3), .A2(_02379__PTR6), .ZN(_02378__PTR33) );
  AND2_X1 U12874 ( .A1(P2_P1_InstQueueRd_Addr_PTR4), .A2(_02379__PTR6), .ZN(_02378__PTR34) );
  AND2_X1 U12875 ( .A1(_02165__PTR0), .A2(_02167__PTR0), .ZN(_02166__PTR0) );
  AND2_X1 U12876 ( .A1(P2_CodeFetch), .A2(_02156__PTR3), .ZN(_02166__PTR1) );
  AND2_X1 U12877 ( .A1(_02154__PTR0), .A2(_02156__PTR0), .ZN(_02155__PTR0) );
  AND2_X1 U12878 ( .A1(_02154__PTR1), .A2(_02148__PTR1), .ZN(_02155__PTR1) );
  AND2_X1 U12879 ( .A1(_02154__PTR2), .A2(_02156__PTR2), .ZN(_02155__PTR2) );
  AND2_X1 U12880 ( .A1(P2_RequestPending), .A2(_02156__PTR3), .ZN(_02155__PTR3) );
  AND2_X1 U12881 ( .A1(_02161__PTR0), .A2(_02163__PTR0), .ZN(_02162__PTR0) );
  AND2_X1 U12882 ( .A1(_02161__PTR1), .A2(_02163__PTR1), .ZN(_02162__PTR1) );
  AND2_X1 U12883 ( .A1(P2_MemoryFetch), .A2(_02156__PTR3), .ZN(_02162__PTR2) );
  AND2_X1 U12884 ( .A1(_02158__PTR0), .A2(_02148__PTR0), .ZN(_02159__PTR0) );
  AND2_X1 U12885 ( .A1(_02158__PTR1), .A2(_02148__PTR1), .ZN(_02159__PTR1) );
  AND2_X1 U12886 ( .A1(P2_ReadRequest), .A2(_02156__PTR3), .ZN(_02159__PTR2) );
  AND2_X1 U12887 ( .A1(P2_rEIP_PTR0), .A2(_02156__PTR3), .ZN(_02394__PTR0) );
  AND2_X1 U12888 ( .A1(P2_rEIP_PTR1), .A2(_02156__PTR3), .ZN(_02394__PTR1) );
  AND2_X1 U12889 ( .A1(P2_rEIP_PTR2), .A2(_02156__PTR3), .ZN(_02394__PTR2) );
  AND2_X1 U12890 ( .A1(P2_rEIP_PTR3), .A2(_02156__PTR3), .ZN(_02394__PTR3) );
  AND2_X1 U12891 ( .A1(P2_rEIP_PTR4), .A2(_02156__PTR3), .ZN(_02394__PTR4) );
  AND2_X1 U12892 ( .A1(P2_rEIP_PTR5), .A2(_02156__PTR3), .ZN(_02394__PTR5) );
  AND2_X1 U12893 ( .A1(P2_rEIP_PTR6), .A2(_02156__PTR3), .ZN(_02394__PTR6) );
  AND2_X1 U12894 ( .A1(P2_rEIP_PTR7), .A2(_02156__PTR3), .ZN(_02394__PTR7) );
  AND2_X1 U12895 ( .A1(P2_rEIP_PTR8), .A2(_02156__PTR3), .ZN(_02394__PTR8) );
  AND2_X1 U12896 ( .A1(P2_rEIP_PTR9), .A2(_02156__PTR3), .ZN(_02394__PTR9) );
  AND2_X1 U12897 ( .A1(P2_rEIP_PTR10), .A2(_02156__PTR3), .ZN(_02394__PTR10) );
  AND2_X1 U12898 ( .A1(P2_rEIP_PTR11), .A2(_02156__PTR3), .ZN(_02394__PTR11) );
  AND2_X1 U12899 ( .A1(P2_rEIP_PTR12), .A2(_02156__PTR3), .ZN(_02394__PTR12) );
  AND2_X1 U12900 ( .A1(P2_rEIP_PTR13), .A2(_02156__PTR3), .ZN(_02394__PTR13) );
  AND2_X1 U12901 ( .A1(P2_rEIP_PTR14), .A2(_02156__PTR3), .ZN(_02394__PTR14) );
  AND2_X1 U12902 ( .A1(P2_rEIP_PTR15), .A2(_02156__PTR3), .ZN(_02394__PTR15) );
  AND2_X1 U12903 ( .A1(P2_rEIP_PTR16), .A2(_02156__PTR3), .ZN(_02394__PTR16) );
  AND2_X1 U12904 ( .A1(P2_rEIP_PTR17), .A2(_02156__PTR3), .ZN(_02394__PTR17) );
  AND2_X1 U12905 ( .A1(P2_rEIP_PTR18), .A2(_02156__PTR3), .ZN(_02394__PTR18) );
  AND2_X1 U12906 ( .A1(P2_rEIP_PTR19), .A2(_02156__PTR3), .ZN(_02394__PTR19) );
  AND2_X1 U12907 ( .A1(P2_rEIP_PTR20), .A2(_02156__PTR3), .ZN(_02394__PTR20) );
  AND2_X1 U12908 ( .A1(P2_rEIP_PTR21), .A2(_02156__PTR3), .ZN(_02394__PTR21) );
  AND2_X1 U12909 ( .A1(P2_rEIP_PTR22), .A2(_02156__PTR3), .ZN(_02394__PTR22) );
  AND2_X1 U12910 ( .A1(P2_rEIP_PTR23), .A2(_02156__PTR3), .ZN(_02394__PTR23) );
  AND2_X1 U12911 ( .A1(P2_rEIP_PTR24), .A2(_02156__PTR3), .ZN(_02394__PTR24) );
  AND2_X1 U12912 ( .A1(P2_rEIP_PTR25), .A2(_02156__PTR3), .ZN(_02394__PTR25) );
  AND2_X1 U12913 ( .A1(P2_rEIP_PTR26), .A2(_02156__PTR3), .ZN(_02394__PTR26) );
  AND2_X1 U12914 ( .A1(P2_rEIP_PTR27), .A2(_02156__PTR3), .ZN(_02394__PTR27) );
  AND2_X1 U12915 ( .A1(P2_rEIP_PTR28), .A2(_02156__PTR3), .ZN(_02394__PTR28) );
  AND2_X1 U12916 ( .A1(P2_rEIP_PTR29), .A2(_02156__PTR3), .ZN(_02394__PTR29) );
  AND2_X1 U12917 ( .A1(P2_rEIP_PTR30), .A2(_02156__PTR3), .ZN(_02394__PTR30) );
  AND2_X1 U12918 ( .A1(P2_rEIP_PTR31), .A2(_02156__PTR3), .ZN(_02394__PTR31) );
  AND2_X1 U12919 ( .A1(_02393__PTR32), .A2(_02163__PTR0), .ZN(_02394__PTR32) );
  AND2_X1 U12920 ( .A1(_02393__PTR33), .A2(_02163__PTR0), .ZN(_02394__PTR33) );
  AND2_X1 U12921 ( .A1(_02393__PTR34), .A2(_02163__PTR0), .ZN(_02394__PTR34) );
  AND2_X1 U12922 ( .A1(_02393__PTR35), .A2(_02163__PTR0), .ZN(_02394__PTR35) );
  AND2_X1 U12923 ( .A1(_02393__PTR36), .A2(_02163__PTR0), .ZN(_02394__PTR36) );
  AND2_X1 U12924 ( .A1(_02393__PTR37), .A2(_02163__PTR0), .ZN(_02394__PTR37) );
  AND2_X1 U12925 ( .A1(_02393__PTR38), .A2(_02163__PTR0), .ZN(_02394__PTR38) );
  AND2_X1 U12926 ( .A1(_02393__PTR39), .A2(_02163__PTR0), .ZN(_02394__PTR39) );
  AND2_X1 U12927 ( .A1(_02393__PTR40), .A2(_02163__PTR0), .ZN(_02394__PTR40) );
  AND2_X1 U12928 ( .A1(_02393__PTR41), .A2(_02163__PTR0), .ZN(_02394__PTR41) );
  AND2_X1 U12929 ( .A1(_02393__PTR42), .A2(_02163__PTR0), .ZN(_02394__PTR42) );
  AND2_X1 U12930 ( .A1(_02393__PTR43), .A2(_02163__PTR0), .ZN(_02394__PTR43) );
  AND2_X1 U12931 ( .A1(_02393__PTR44), .A2(_02163__PTR0), .ZN(_02394__PTR44) );
  AND2_X1 U12932 ( .A1(_02393__PTR45), .A2(_02163__PTR0), .ZN(_02394__PTR45) );
  AND2_X1 U12933 ( .A1(_02393__PTR46), .A2(_02163__PTR0), .ZN(_02394__PTR46) );
  AND2_X1 U12934 ( .A1(_02393__PTR47), .A2(_02163__PTR0), .ZN(_02394__PTR47) );
  AND2_X1 U12935 ( .A1(_02393__PTR48), .A2(_02163__PTR0), .ZN(_02394__PTR48) );
  AND2_X1 U12936 ( .A1(_02393__PTR49), .A2(_02163__PTR0), .ZN(_02394__PTR49) );
  AND2_X1 U12937 ( .A1(_02393__PTR50), .A2(_02163__PTR0), .ZN(_02394__PTR50) );
  AND2_X1 U12938 ( .A1(_02393__PTR51), .A2(_02163__PTR0), .ZN(_02394__PTR51) );
  AND2_X1 U12939 ( .A1(_02393__PTR52), .A2(_02163__PTR0), .ZN(_02394__PTR52) );
  AND2_X1 U12940 ( .A1(_02393__PTR53), .A2(_02163__PTR0), .ZN(_02394__PTR53) );
  AND2_X1 U12941 ( .A1(_02393__PTR54), .A2(_02163__PTR0), .ZN(_02394__PTR54) );
  AND2_X1 U12942 ( .A1(_02393__PTR55), .A2(_02163__PTR0), .ZN(_02394__PTR55) );
  AND2_X1 U12943 ( .A1(_02393__PTR56), .A2(_02163__PTR0), .ZN(_02394__PTR56) );
  AND2_X1 U12944 ( .A1(_02393__PTR57), .A2(_02163__PTR0), .ZN(_02394__PTR57) );
  AND2_X1 U12945 ( .A1(_02393__PTR58), .A2(_02163__PTR0), .ZN(_02394__PTR58) );
  AND2_X1 U12946 ( .A1(_02393__PTR59), .A2(_02163__PTR0), .ZN(_02394__PTR59) );
  AND2_X1 U12947 ( .A1(_02393__PTR60), .A2(_02163__PTR0), .ZN(_02394__PTR60) );
  AND2_X1 U12948 ( .A1(_02393__PTR61), .A2(_02163__PTR0), .ZN(_02394__PTR61) );
  AND2_X1 U12949 ( .A1(_02393__PTR62), .A2(_02163__PTR0), .ZN(_02394__PTR62) );
  AND2_X1 U12950 ( .A1(_02393__PTR63), .A2(_02163__PTR0), .ZN(_02394__PTR63) );
  AND2_X1 U12951 ( .A1(_02393__PTR64), .A2(_02156__PTR2), .ZN(_02394__PTR64) );
  AND2_X1 U12952 ( .A1(_02393__PTR65), .A2(_02156__PTR2), .ZN(_02394__PTR65) );
  AND2_X1 U12953 ( .A1(_02393__PTR66), .A2(_02156__PTR2), .ZN(_02394__PTR66) );
  AND2_X1 U12954 ( .A1(_02393__PTR67), .A2(_02156__PTR2), .ZN(_02394__PTR67) );
  AND2_X1 U12955 ( .A1(_02393__PTR68), .A2(_02156__PTR2), .ZN(_02394__PTR68) );
  AND2_X1 U12956 ( .A1(_02393__PTR69), .A2(_02156__PTR2), .ZN(_02394__PTR69) );
  AND2_X1 U12957 ( .A1(_02393__PTR70), .A2(_02156__PTR2), .ZN(_02394__PTR70) );
  AND2_X1 U12958 ( .A1(_02393__PTR71), .A2(_02156__PTR2), .ZN(_02394__PTR71) );
  AND2_X1 U12959 ( .A1(_02393__PTR72), .A2(_02156__PTR2), .ZN(_02394__PTR72) );
  AND2_X1 U12960 ( .A1(_02393__PTR73), .A2(_02156__PTR2), .ZN(_02394__PTR73) );
  AND2_X1 U12961 ( .A1(_02393__PTR74), .A2(_02156__PTR2), .ZN(_02394__PTR74) );
  AND2_X1 U12962 ( .A1(_02393__PTR75), .A2(_02156__PTR2), .ZN(_02394__PTR75) );
  AND2_X1 U12963 ( .A1(_02393__PTR76), .A2(_02156__PTR2), .ZN(_02394__PTR76) );
  AND2_X1 U12964 ( .A1(_02393__PTR77), .A2(_02156__PTR2), .ZN(_02394__PTR77) );
  AND2_X1 U12965 ( .A1(_02393__PTR78), .A2(_02156__PTR2), .ZN(_02394__PTR78) );
  AND2_X1 U12966 ( .A1(_02393__PTR79), .A2(_02156__PTR2), .ZN(_02394__PTR79) );
  AND2_X1 U12967 ( .A1(_02393__PTR80), .A2(_02156__PTR2), .ZN(_02394__PTR80) );
  AND2_X1 U12968 ( .A1(_02393__PTR81), .A2(_02156__PTR2), .ZN(_02394__PTR81) );
  AND2_X1 U12969 ( .A1(_02393__PTR82), .A2(_02156__PTR2), .ZN(_02394__PTR82) );
  AND2_X1 U12970 ( .A1(_02393__PTR83), .A2(_02156__PTR2), .ZN(_02394__PTR83) );
  AND2_X1 U12971 ( .A1(_02393__PTR84), .A2(_02156__PTR2), .ZN(_02394__PTR84) );
  AND2_X1 U12972 ( .A1(_02393__PTR85), .A2(_02156__PTR2), .ZN(_02394__PTR85) );
  AND2_X1 U12973 ( .A1(_02393__PTR86), .A2(_02156__PTR2), .ZN(_02394__PTR86) );
  AND2_X1 U12974 ( .A1(_02393__PTR87), .A2(_02156__PTR2), .ZN(_02394__PTR87) );
  AND2_X1 U12975 ( .A1(_02393__PTR88), .A2(_02156__PTR2), .ZN(_02394__PTR88) );
  AND2_X1 U12976 ( .A1(_02393__PTR89), .A2(_02156__PTR2), .ZN(_02394__PTR89) );
  AND2_X1 U12977 ( .A1(_02393__PTR90), .A2(_02156__PTR2), .ZN(_02394__PTR90) );
  AND2_X1 U12978 ( .A1(_02393__PTR91), .A2(_02156__PTR2), .ZN(_02394__PTR91) );
  AND2_X1 U12979 ( .A1(_02393__PTR92), .A2(_02156__PTR2), .ZN(_02394__PTR92) );
  AND2_X1 U12980 ( .A1(_02393__PTR93), .A2(_02156__PTR2), .ZN(_02394__PTR93) );
  AND2_X1 U12981 ( .A1(_02393__PTR94), .A2(_02156__PTR2), .ZN(_02394__PTR94) );
  AND2_X1 U12982 ( .A1(_02393__PTR95), .A2(_02156__PTR2), .ZN(_02394__PTR95) );
  AND2_X1 U12983 ( .A1(_02393__PTR96), .A2(_02379__PTR4), .ZN(_02394__PTR96) );
  AND2_X1 U12984 ( .A1(_02393__PTR97), .A2(_02379__PTR4), .ZN(_02394__PTR97) );
  AND2_X1 U12985 ( .A1(_02393__PTR98), .A2(_02379__PTR4), .ZN(_02394__PTR98) );
  AND2_X1 U12986 ( .A1(_02393__PTR99), .A2(_02379__PTR4), .ZN(_02394__PTR99) );
  AND2_X1 U12987 ( .A1(_02393__PTR100), .A2(_02379__PTR4), .ZN(_02394__PTR100) );
  AND2_X1 U12988 ( .A1(_02393__PTR101), .A2(_02379__PTR4), .ZN(_02394__PTR101) );
  AND2_X1 U12989 ( .A1(_02393__PTR102), .A2(_02379__PTR4), .ZN(_02394__PTR102) );
  AND2_X1 U12990 ( .A1(_02393__PTR103), .A2(_02379__PTR4), .ZN(_02394__PTR103) );
  AND2_X1 U12991 ( .A1(_02393__PTR104), .A2(_02379__PTR4), .ZN(_02394__PTR104) );
  AND2_X1 U12992 ( .A1(_02393__PTR105), .A2(_02379__PTR4), .ZN(_02394__PTR105) );
  AND2_X1 U12993 ( .A1(_02393__PTR106), .A2(_02379__PTR4), .ZN(_02394__PTR106) );
  AND2_X1 U12994 ( .A1(_02393__PTR107), .A2(_02379__PTR4), .ZN(_02394__PTR107) );
  AND2_X1 U12995 ( .A1(_02393__PTR108), .A2(_02379__PTR4), .ZN(_02394__PTR108) );
  AND2_X1 U12996 ( .A1(_02393__PTR109), .A2(_02379__PTR4), .ZN(_02394__PTR109) );
  AND2_X1 U12997 ( .A1(_02393__PTR110), .A2(_02379__PTR4), .ZN(_02394__PTR110) );
  AND2_X1 U12998 ( .A1(_02393__PTR111), .A2(_02379__PTR4), .ZN(_02394__PTR111) );
  AND2_X1 U12999 ( .A1(_02393__PTR112), .A2(_02379__PTR4), .ZN(_02394__PTR112) );
  AND2_X1 U13000 ( .A1(_02393__PTR113), .A2(_02379__PTR4), .ZN(_02394__PTR113) );
  AND2_X1 U13001 ( .A1(_02393__PTR114), .A2(_02379__PTR4), .ZN(_02394__PTR114) );
  AND2_X1 U13002 ( .A1(_02393__PTR115), .A2(_02379__PTR4), .ZN(_02394__PTR115) );
  AND2_X1 U13003 ( .A1(_02393__PTR116), .A2(_02379__PTR4), .ZN(_02394__PTR116) );
  AND2_X1 U13004 ( .A1(_02393__PTR117), .A2(_02379__PTR4), .ZN(_02394__PTR117) );
  AND2_X1 U13005 ( .A1(_02393__PTR118), .A2(_02379__PTR4), .ZN(_02394__PTR118) );
  AND2_X1 U13006 ( .A1(_02393__PTR119), .A2(_02379__PTR4), .ZN(_02394__PTR119) );
  AND2_X1 U13007 ( .A1(_02393__PTR120), .A2(_02379__PTR4), .ZN(_02394__PTR120) );
  AND2_X1 U13008 ( .A1(_02393__PTR121), .A2(_02379__PTR4), .ZN(_02394__PTR121) );
  AND2_X1 U13009 ( .A1(_02393__PTR122), .A2(_02379__PTR4), .ZN(_02394__PTR122) );
  AND2_X1 U13010 ( .A1(_02393__PTR123), .A2(_02379__PTR4), .ZN(_02394__PTR123) );
  AND2_X1 U13011 ( .A1(_02393__PTR124), .A2(_02379__PTR4), .ZN(_02394__PTR124) );
  AND2_X1 U13012 ( .A1(_02393__PTR125), .A2(_02379__PTR4), .ZN(_02394__PTR125) );
  AND2_X1 U13013 ( .A1(_02393__PTR126), .A2(_02379__PTR4), .ZN(_02394__PTR126) );
  AND2_X1 U13014 ( .A1(_02393__PTR127), .A2(_02379__PTR4), .ZN(_02394__PTR127) );
  AND2_X1 U13015 ( .A1(_02373__PTR0), .A2(_02375__PTR0), .ZN(_02374__PTR0) );
  AND2_X1 U13016 ( .A1(_02373__PTR1), .A2(_02375__PTR0), .ZN(_02374__PTR1) );
  AND2_X1 U13017 ( .A1(_02373__PTR2), .A2(_02375__PTR0), .ZN(_02374__PTR2) );
  AND2_X1 U13018 ( .A1(_02373__PTR3), .A2(_02375__PTR0), .ZN(_02374__PTR3) );
  AND2_X1 U13019 ( .A1(_02373__PTR4), .A2(_02375__PTR0), .ZN(_02374__PTR4) );
  AND2_X1 U13020 ( .A1(_02373__PTR5), .A2(_02375__PTR0), .ZN(_02374__PTR5) );
  AND2_X1 U13021 ( .A1(_02373__PTR6), .A2(_02375__PTR0), .ZN(_02374__PTR6) );
  AND2_X1 U13022 ( .A1(_02373__PTR7), .A2(_02375__PTR0), .ZN(_02374__PTR7) );
  AND2_X1 U13023 ( .A1(_02373__PTR8), .A2(_02375__PTR0), .ZN(_02374__PTR8) );
  AND2_X1 U13024 ( .A1(_02373__PTR9), .A2(_02375__PTR0), .ZN(_02374__PTR9) );
  AND2_X1 U13025 ( .A1(_02373__PTR10), .A2(_02375__PTR0), .ZN(_02374__PTR10) );
  AND2_X1 U13026 ( .A1(_02373__PTR11), .A2(_02375__PTR0), .ZN(_02374__PTR11) );
  AND2_X1 U13027 ( .A1(_02373__PTR12), .A2(_02375__PTR0), .ZN(_02374__PTR12) );
  AND2_X1 U13028 ( .A1(_02373__PTR13), .A2(_02375__PTR0), .ZN(_02374__PTR13) );
  AND2_X1 U13029 ( .A1(_02373__PTR14), .A2(_02375__PTR0), .ZN(_02374__PTR14) );
  AND2_X1 U13030 ( .A1(_02373__PTR15), .A2(_02375__PTR0), .ZN(_02374__PTR15) );
  AND2_X1 U13031 ( .A1(_02373__PTR16), .A2(_02375__PTR0), .ZN(_02374__PTR16) );
  AND2_X1 U13032 ( .A1(_02373__PTR17), .A2(_02375__PTR0), .ZN(_02374__PTR17) );
  AND2_X1 U13033 ( .A1(_02373__PTR18), .A2(_02375__PTR0), .ZN(_02374__PTR18) );
  AND2_X1 U13034 ( .A1(_02373__PTR19), .A2(_02375__PTR0), .ZN(_02374__PTR19) );
  AND2_X1 U13035 ( .A1(_02373__PTR20), .A2(_02375__PTR0), .ZN(_02374__PTR20) );
  AND2_X1 U13036 ( .A1(_02373__PTR21), .A2(_02375__PTR0), .ZN(_02374__PTR21) );
  AND2_X1 U13037 ( .A1(_02373__PTR22), .A2(_02375__PTR0), .ZN(_02374__PTR22) );
  AND2_X1 U13038 ( .A1(_02373__PTR23), .A2(_02375__PTR0), .ZN(_02374__PTR23) );
  AND2_X1 U13039 ( .A1(_02373__PTR24), .A2(_02375__PTR0), .ZN(_02374__PTR24) );
  AND2_X1 U13040 ( .A1(_02373__PTR25), .A2(_02375__PTR0), .ZN(_02374__PTR25) );
  AND2_X1 U13041 ( .A1(_02373__PTR26), .A2(_02375__PTR0), .ZN(_02374__PTR26) );
  AND2_X1 U13042 ( .A1(_02373__PTR27), .A2(_02375__PTR0), .ZN(_02374__PTR27) );
  AND2_X1 U13043 ( .A1(_02373__PTR28), .A2(_02375__PTR0), .ZN(_02374__PTR28) );
  AND2_X1 U13044 ( .A1(_02373__PTR29), .A2(_02375__PTR0), .ZN(_02374__PTR29) );
  AND2_X1 U13045 ( .A1(_02373__PTR30), .A2(_02375__PTR0), .ZN(_02374__PTR30) );
  AND2_X1 U13046 ( .A1(_02373__PTR31), .A2(_02375__PTR0), .ZN(_02374__PTR31) );
  AND2_X1 U13047 ( .A1(P2_P1_InstAddrPointer_PTR0), .A2(_02375__PTR1), .ZN(_02374__PTR32) );
  AND2_X1 U13048 ( .A1(_02373__PTR33), .A2(_02375__PTR1), .ZN(_02374__PTR33) );
  AND2_X1 U13049 ( .A1(_02373__PTR34), .A2(_02375__PTR1), .ZN(_02374__PTR34) );
  AND2_X1 U13050 ( .A1(_02373__PTR35), .A2(_02375__PTR1), .ZN(_02374__PTR35) );
  AND2_X1 U13051 ( .A1(_02373__PTR36), .A2(_02375__PTR1), .ZN(_02374__PTR36) );
  AND2_X1 U13052 ( .A1(_02373__PTR37), .A2(_02375__PTR1), .ZN(_02374__PTR37) );
  AND2_X1 U13053 ( .A1(_02373__PTR38), .A2(_02375__PTR1), .ZN(_02374__PTR38) );
  AND2_X1 U13054 ( .A1(_02373__PTR39), .A2(_02375__PTR1), .ZN(_02374__PTR39) );
  AND2_X1 U13055 ( .A1(_02373__PTR40), .A2(_02375__PTR1), .ZN(_02374__PTR40) );
  AND2_X1 U13056 ( .A1(_02373__PTR41), .A2(_02375__PTR1), .ZN(_02374__PTR41) );
  AND2_X1 U13057 ( .A1(_02373__PTR42), .A2(_02375__PTR1), .ZN(_02374__PTR42) );
  AND2_X1 U13058 ( .A1(_02373__PTR43), .A2(_02375__PTR1), .ZN(_02374__PTR43) );
  AND2_X1 U13059 ( .A1(_02373__PTR44), .A2(_02375__PTR1), .ZN(_02374__PTR44) );
  AND2_X1 U13060 ( .A1(_02373__PTR45), .A2(_02375__PTR1), .ZN(_02374__PTR45) );
  AND2_X1 U13061 ( .A1(_02373__PTR46), .A2(_02375__PTR1), .ZN(_02374__PTR46) );
  AND2_X1 U13062 ( .A1(_02373__PTR47), .A2(_02375__PTR1), .ZN(_02374__PTR47) );
  AND2_X1 U13063 ( .A1(_02373__PTR48), .A2(_02375__PTR1), .ZN(_02374__PTR48) );
  AND2_X1 U13064 ( .A1(_02373__PTR49), .A2(_02375__PTR1), .ZN(_02374__PTR49) );
  AND2_X1 U13065 ( .A1(_02373__PTR50), .A2(_02375__PTR1), .ZN(_02374__PTR50) );
  AND2_X1 U13066 ( .A1(_02373__PTR51), .A2(_02375__PTR1), .ZN(_02374__PTR51) );
  AND2_X1 U13067 ( .A1(_02373__PTR52), .A2(_02375__PTR1), .ZN(_02374__PTR52) );
  AND2_X1 U13068 ( .A1(_02373__PTR53), .A2(_02375__PTR1), .ZN(_02374__PTR53) );
  AND2_X1 U13069 ( .A1(_02373__PTR54), .A2(_02375__PTR1), .ZN(_02374__PTR54) );
  AND2_X1 U13070 ( .A1(_02373__PTR55), .A2(_02375__PTR1), .ZN(_02374__PTR55) );
  AND2_X1 U13071 ( .A1(_02373__PTR56), .A2(_02375__PTR1), .ZN(_02374__PTR56) );
  AND2_X1 U13072 ( .A1(_02373__PTR57), .A2(_02375__PTR1), .ZN(_02374__PTR57) );
  AND2_X1 U13073 ( .A1(_02373__PTR58), .A2(_02375__PTR1), .ZN(_02374__PTR58) );
  AND2_X1 U13074 ( .A1(_02373__PTR59), .A2(_02375__PTR1), .ZN(_02374__PTR59) );
  AND2_X1 U13075 ( .A1(_02373__PTR60), .A2(_02375__PTR1), .ZN(_02374__PTR60) );
  AND2_X1 U13076 ( .A1(_02373__PTR61), .A2(_02375__PTR1), .ZN(_02374__PTR61) );
  AND2_X1 U13077 ( .A1(_02373__PTR62), .A2(_02375__PTR1), .ZN(_02374__PTR62) );
  AND2_X1 U13078 ( .A1(_02373__PTR63), .A2(_02375__PTR1), .ZN(_02374__PTR63) );
  AND2_X1 U13079 ( .A1(P2_P1_InstAddrPointer_PTR0), .A2(_02148__PTR0), .ZN(_02374__PTR64) );
  AND2_X1 U13080 ( .A1(_02373__PTR65), .A2(_02148__PTR0), .ZN(_02374__PTR65) );
  AND2_X1 U13081 ( .A1(_02373__PTR66), .A2(_02148__PTR0), .ZN(_02374__PTR66) );
  AND2_X1 U13082 ( .A1(_02373__PTR67), .A2(_02148__PTR0), .ZN(_02374__PTR67) );
  AND2_X1 U13083 ( .A1(_02373__PTR68), .A2(_02148__PTR0), .ZN(_02374__PTR68) );
  AND2_X1 U13084 ( .A1(_02373__PTR69), .A2(_02148__PTR0), .ZN(_02374__PTR69) );
  AND2_X1 U13085 ( .A1(_02373__PTR70), .A2(_02148__PTR0), .ZN(_02374__PTR70) );
  AND2_X1 U13086 ( .A1(_02373__PTR71), .A2(_02148__PTR0), .ZN(_02374__PTR71) );
  AND2_X1 U13087 ( .A1(_02373__PTR72), .A2(_02148__PTR0), .ZN(_02374__PTR72) );
  AND2_X1 U13088 ( .A1(_02373__PTR73), .A2(_02148__PTR0), .ZN(_02374__PTR73) );
  AND2_X1 U13089 ( .A1(_02373__PTR74), .A2(_02148__PTR0), .ZN(_02374__PTR74) );
  AND2_X1 U13090 ( .A1(_02373__PTR75), .A2(_02148__PTR0), .ZN(_02374__PTR75) );
  AND2_X1 U13091 ( .A1(_02373__PTR76), .A2(_02148__PTR0), .ZN(_02374__PTR76) );
  AND2_X1 U13092 ( .A1(_02373__PTR77), .A2(_02148__PTR0), .ZN(_02374__PTR77) );
  AND2_X1 U13093 ( .A1(_02373__PTR78), .A2(_02148__PTR0), .ZN(_02374__PTR78) );
  AND2_X1 U13094 ( .A1(_02373__PTR79), .A2(_02148__PTR0), .ZN(_02374__PTR79) );
  AND2_X1 U13095 ( .A1(_02373__PTR80), .A2(_02148__PTR0), .ZN(_02374__PTR80) );
  AND2_X1 U13096 ( .A1(_02373__PTR81), .A2(_02148__PTR0), .ZN(_02374__PTR81) );
  AND2_X1 U13097 ( .A1(_02373__PTR82), .A2(_02148__PTR0), .ZN(_02374__PTR82) );
  AND2_X1 U13098 ( .A1(_02373__PTR83), .A2(_02148__PTR0), .ZN(_02374__PTR83) );
  AND2_X1 U13099 ( .A1(_02373__PTR84), .A2(_02148__PTR0), .ZN(_02374__PTR84) );
  AND2_X1 U13100 ( .A1(_02373__PTR85), .A2(_02148__PTR0), .ZN(_02374__PTR85) );
  AND2_X1 U13101 ( .A1(_02373__PTR86), .A2(_02148__PTR0), .ZN(_02374__PTR86) );
  AND2_X1 U13102 ( .A1(_02373__PTR87), .A2(_02148__PTR0), .ZN(_02374__PTR87) );
  AND2_X1 U13103 ( .A1(_02373__PTR88), .A2(_02148__PTR0), .ZN(_02374__PTR88) );
  AND2_X1 U13104 ( .A1(_02373__PTR89), .A2(_02148__PTR0), .ZN(_02374__PTR89) );
  AND2_X1 U13105 ( .A1(_02373__PTR90), .A2(_02148__PTR0), .ZN(_02374__PTR90) );
  AND2_X1 U13106 ( .A1(_02373__PTR91), .A2(_02148__PTR0), .ZN(_02374__PTR91) );
  AND2_X1 U13107 ( .A1(_02373__PTR92), .A2(_02148__PTR0), .ZN(_02374__PTR92) );
  AND2_X1 U13108 ( .A1(_02373__PTR93), .A2(_02148__PTR0), .ZN(_02374__PTR93) );
  AND2_X1 U13109 ( .A1(_02373__PTR94), .A2(_02148__PTR0), .ZN(_02374__PTR94) );
  AND2_X1 U13110 ( .A1(_02373__PTR95), .A2(_02148__PTR0), .ZN(_02374__PTR95) );
  AND2_X1 U13111 ( .A1(P2_P1_InstAddrPointer_PTR0), .A2(_02148__PTR1), .ZN(_02374__PTR96) );
  AND2_X1 U13112 ( .A1(_02373__PTR97), .A2(_02148__PTR1), .ZN(_02374__PTR97) );
  AND2_X1 U13113 ( .A1(_02373__PTR98), .A2(_02148__PTR1), .ZN(_02374__PTR98) );
  AND2_X1 U13114 ( .A1(_02373__PTR99), .A2(_02148__PTR1), .ZN(_02374__PTR99) );
  AND2_X1 U13115 ( .A1(_02373__PTR100), .A2(_02148__PTR1), .ZN(_02374__PTR100) );
  AND2_X1 U13116 ( .A1(_02373__PTR101), .A2(_02148__PTR1), .ZN(_02374__PTR101) );
  AND2_X1 U13117 ( .A1(_02373__PTR102), .A2(_02148__PTR1), .ZN(_02374__PTR102) );
  AND2_X1 U13118 ( .A1(_02373__PTR103), .A2(_02148__PTR1), .ZN(_02374__PTR103) );
  AND2_X1 U13119 ( .A1(_02373__PTR104), .A2(_02148__PTR1), .ZN(_02374__PTR104) );
  AND2_X1 U13120 ( .A1(_02373__PTR105), .A2(_02148__PTR1), .ZN(_02374__PTR105) );
  AND2_X1 U13121 ( .A1(_02373__PTR106), .A2(_02148__PTR1), .ZN(_02374__PTR106) );
  AND2_X1 U13122 ( .A1(_02373__PTR107), .A2(_02148__PTR1), .ZN(_02374__PTR107) );
  AND2_X1 U13123 ( .A1(_02373__PTR108), .A2(_02148__PTR1), .ZN(_02374__PTR108) );
  AND2_X1 U13124 ( .A1(_02373__PTR109), .A2(_02148__PTR1), .ZN(_02374__PTR109) );
  AND2_X1 U13125 ( .A1(_02373__PTR110), .A2(_02148__PTR1), .ZN(_02374__PTR110) );
  AND2_X1 U13126 ( .A1(_02373__PTR111), .A2(_02148__PTR1), .ZN(_02374__PTR111) );
  AND2_X1 U13127 ( .A1(_02373__PTR112), .A2(_02148__PTR1), .ZN(_02374__PTR112) );
  AND2_X1 U13128 ( .A1(_02373__PTR113), .A2(_02148__PTR1), .ZN(_02374__PTR113) );
  AND2_X1 U13129 ( .A1(_02373__PTR114), .A2(_02148__PTR1), .ZN(_02374__PTR114) );
  AND2_X1 U13130 ( .A1(_02373__PTR115), .A2(_02148__PTR1), .ZN(_02374__PTR115) );
  AND2_X1 U13131 ( .A1(_02373__PTR116), .A2(_02148__PTR1), .ZN(_02374__PTR116) );
  AND2_X1 U13132 ( .A1(_02373__PTR117), .A2(_02148__PTR1), .ZN(_02374__PTR117) );
  AND2_X1 U13133 ( .A1(_02373__PTR118), .A2(_02148__PTR1), .ZN(_02374__PTR118) );
  AND2_X1 U13134 ( .A1(_02373__PTR119), .A2(_02148__PTR1), .ZN(_02374__PTR119) );
  AND2_X1 U13135 ( .A1(_02373__PTR120), .A2(_02148__PTR1), .ZN(_02374__PTR120) );
  AND2_X1 U13136 ( .A1(_02373__PTR121), .A2(_02148__PTR1), .ZN(_02374__PTR121) );
  AND2_X1 U13137 ( .A1(_02373__PTR122), .A2(_02148__PTR1), .ZN(_02374__PTR122) );
  AND2_X1 U13138 ( .A1(_02373__PTR123), .A2(_02148__PTR1), .ZN(_02374__PTR123) );
  AND2_X1 U13139 ( .A1(_02373__PTR124), .A2(_02148__PTR1), .ZN(_02374__PTR124) );
  AND2_X1 U13140 ( .A1(_02373__PTR125), .A2(_02148__PTR1), .ZN(_02374__PTR125) );
  AND2_X1 U13141 ( .A1(_02373__PTR126), .A2(_02148__PTR1), .ZN(_02374__PTR126) );
  AND2_X1 U13142 ( .A1(_02373__PTR127), .A2(_02148__PTR1), .ZN(_02374__PTR127) );
  AND2_X1 U13143 ( .A1(_02373__PTR128), .A2(_02375__PTR4), .ZN(_02374__PTR128) );
  AND2_X1 U13144 ( .A1(_02373__PTR129), .A2(_02375__PTR4), .ZN(_02374__PTR129) );
  AND2_X1 U13145 ( .A1(_02373__PTR130), .A2(_02375__PTR4), .ZN(_02374__PTR130) );
  AND2_X1 U13146 ( .A1(_02373__PTR131), .A2(_02375__PTR4), .ZN(_02374__PTR131) );
  AND2_X1 U13147 ( .A1(_02373__PTR132), .A2(_02375__PTR4), .ZN(_02374__PTR132) );
  AND2_X1 U13148 ( .A1(_02373__PTR133), .A2(_02375__PTR4), .ZN(_02374__PTR133) );
  AND2_X1 U13149 ( .A1(_02373__PTR134), .A2(_02375__PTR4), .ZN(_02374__PTR134) );
  AND2_X1 U13150 ( .A1(_02373__PTR135), .A2(_02375__PTR4), .ZN(_02374__PTR135) );
  AND2_X1 U13151 ( .A1(_02373__PTR136), .A2(_02375__PTR4), .ZN(_02374__PTR136) );
  AND2_X1 U13152 ( .A1(_02373__PTR137), .A2(_02375__PTR4), .ZN(_02374__PTR137) );
  AND2_X1 U13153 ( .A1(_02373__PTR138), .A2(_02375__PTR4), .ZN(_02374__PTR138) );
  AND2_X1 U13154 ( .A1(_02373__PTR139), .A2(_02375__PTR4), .ZN(_02374__PTR139) );
  AND2_X1 U13155 ( .A1(_02373__PTR140), .A2(_02375__PTR4), .ZN(_02374__PTR140) );
  AND2_X1 U13156 ( .A1(_02373__PTR141), .A2(_02375__PTR4), .ZN(_02374__PTR141) );
  AND2_X1 U13157 ( .A1(_02373__PTR142), .A2(_02375__PTR4), .ZN(_02374__PTR142) );
  AND2_X1 U13158 ( .A1(_02373__PTR143), .A2(_02375__PTR4), .ZN(_02374__PTR143) );
  AND2_X1 U13159 ( .A1(_02373__PTR144), .A2(_02375__PTR4), .ZN(_02374__PTR144) );
  AND2_X1 U13160 ( .A1(_02373__PTR145), .A2(_02375__PTR4), .ZN(_02374__PTR145) );
  AND2_X1 U13161 ( .A1(_02373__PTR146), .A2(_02375__PTR4), .ZN(_02374__PTR146) );
  AND2_X1 U13162 ( .A1(_02373__PTR147), .A2(_02375__PTR4), .ZN(_02374__PTR147) );
  AND2_X1 U13163 ( .A1(_02373__PTR148), .A2(_02375__PTR4), .ZN(_02374__PTR148) );
  AND2_X1 U13164 ( .A1(_02373__PTR149), .A2(_02375__PTR4), .ZN(_02374__PTR149) );
  AND2_X1 U13165 ( .A1(_02373__PTR150), .A2(_02375__PTR4), .ZN(_02374__PTR150) );
  AND2_X1 U13166 ( .A1(_02373__PTR151), .A2(_02375__PTR4), .ZN(_02374__PTR151) );
  AND2_X1 U13167 ( .A1(_02373__PTR152), .A2(_02375__PTR4), .ZN(_02374__PTR152) );
  AND2_X1 U13168 ( .A1(_02373__PTR153), .A2(_02375__PTR4), .ZN(_02374__PTR153) );
  AND2_X1 U13169 ( .A1(_02373__PTR154), .A2(_02375__PTR4), .ZN(_02374__PTR154) );
  AND2_X1 U13170 ( .A1(_02373__PTR155), .A2(_02375__PTR4), .ZN(_02374__PTR155) );
  AND2_X1 U13171 ( .A1(_02373__PTR156), .A2(_02375__PTR4), .ZN(_02374__PTR156) );
  AND2_X1 U13172 ( .A1(_02373__PTR157), .A2(_02375__PTR4), .ZN(_02374__PTR157) );
  AND2_X1 U13173 ( .A1(_02373__PTR158), .A2(_02375__PTR4), .ZN(_02374__PTR158) );
  AND2_X1 U13174 ( .A1(_02373__PTR159), .A2(_02375__PTR4), .ZN(_02374__PTR159) );
  AND2_X1 U13175 ( .A1(_02373__PTR160), .A2(_02148__PTR2), .ZN(_02374__PTR160) );
  AND2_X1 U13176 ( .A1(_02373__PTR161), .A2(_02148__PTR2), .ZN(_02374__PTR161) );
  AND2_X1 U13177 ( .A1(_02373__PTR162), .A2(_02148__PTR2), .ZN(_02374__PTR162) );
  AND2_X1 U13178 ( .A1(_02373__PTR163), .A2(_02148__PTR2), .ZN(_02374__PTR163) );
  AND2_X1 U13179 ( .A1(_02373__PTR164), .A2(_02148__PTR2), .ZN(_02374__PTR164) );
  AND2_X1 U13180 ( .A1(_02373__PTR165), .A2(_02148__PTR2), .ZN(_02374__PTR165) );
  AND2_X1 U13181 ( .A1(_02373__PTR166), .A2(_02148__PTR2), .ZN(_02374__PTR166) );
  AND2_X1 U13182 ( .A1(_02373__PTR167), .A2(_02148__PTR2), .ZN(_02374__PTR167) );
  AND2_X1 U13183 ( .A1(_02373__PTR168), .A2(_02148__PTR2), .ZN(_02374__PTR168) );
  AND2_X1 U13184 ( .A1(_02373__PTR169), .A2(_02148__PTR2), .ZN(_02374__PTR169) );
  AND2_X1 U13185 ( .A1(_02373__PTR170), .A2(_02148__PTR2), .ZN(_02374__PTR170) );
  AND2_X1 U13186 ( .A1(_02373__PTR171), .A2(_02148__PTR2), .ZN(_02374__PTR171) );
  AND2_X1 U13187 ( .A1(_02373__PTR172), .A2(_02148__PTR2), .ZN(_02374__PTR172) );
  AND2_X1 U13188 ( .A1(_02373__PTR173), .A2(_02148__PTR2), .ZN(_02374__PTR173) );
  AND2_X1 U13189 ( .A1(_02373__PTR174), .A2(_02148__PTR2), .ZN(_02374__PTR174) );
  AND2_X1 U13190 ( .A1(_02373__PTR175), .A2(_02148__PTR2), .ZN(_02374__PTR175) );
  AND2_X1 U13191 ( .A1(_02373__PTR176), .A2(_02148__PTR2), .ZN(_02374__PTR176) );
  AND2_X1 U13192 ( .A1(_02373__PTR177), .A2(_02148__PTR2), .ZN(_02374__PTR177) );
  AND2_X1 U13193 ( .A1(_02373__PTR178), .A2(_02148__PTR2), .ZN(_02374__PTR178) );
  AND2_X1 U13194 ( .A1(_02373__PTR179), .A2(_02148__PTR2), .ZN(_02374__PTR179) );
  AND2_X1 U13195 ( .A1(_02373__PTR180), .A2(_02148__PTR2), .ZN(_02374__PTR180) );
  AND2_X1 U13196 ( .A1(_02373__PTR181), .A2(_02148__PTR2), .ZN(_02374__PTR181) );
  AND2_X1 U13197 ( .A1(_02373__PTR182), .A2(_02148__PTR2), .ZN(_02374__PTR182) );
  AND2_X1 U13198 ( .A1(_02373__PTR183), .A2(_02148__PTR2), .ZN(_02374__PTR183) );
  AND2_X1 U13199 ( .A1(_02373__PTR184), .A2(_02148__PTR2), .ZN(_02374__PTR184) );
  AND2_X1 U13200 ( .A1(_02373__PTR185), .A2(_02148__PTR2), .ZN(_02374__PTR185) );
  AND2_X1 U13201 ( .A1(_02373__PTR186), .A2(_02148__PTR2), .ZN(_02374__PTR186) );
  AND2_X1 U13202 ( .A1(_02373__PTR187), .A2(_02148__PTR2), .ZN(_02374__PTR187) );
  AND2_X1 U13203 ( .A1(_02373__PTR188), .A2(_02148__PTR2), .ZN(_02374__PTR188) );
  AND2_X1 U13204 ( .A1(_02373__PTR189), .A2(_02148__PTR2), .ZN(_02374__PTR189) );
  AND2_X1 U13205 ( .A1(_02373__PTR190), .A2(_02148__PTR2), .ZN(_02374__PTR190) );
  AND2_X1 U13206 ( .A1(_02373__PTR191), .A2(_02148__PTR2), .ZN(_02374__PTR191) );
  AND2_X1 U13207 ( .A1(_02373__PTR192), .A2(_02148__PTR3), .ZN(_02374__PTR192) );
  AND2_X1 U13208 ( .A1(_02373__PTR193), .A2(_02148__PTR3), .ZN(_02374__PTR193) );
  AND2_X1 U13209 ( .A1(_02373__PTR194), .A2(_02148__PTR3), .ZN(_02374__PTR194) );
  AND2_X1 U13210 ( .A1(_02373__PTR195), .A2(_02148__PTR3), .ZN(_02374__PTR195) );
  AND2_X1 U13211 ( .A1(_02373__PTR196), .A2(_02148__PTR3), .ZN(_02374__PTR196) );
  AND2_X1 U13212 ( .A1(_02373__PTR197), .A2(_02148__PTR3), .ZN(_02374__PTR197) );
  AND2_X1 U13213 ( .A1(_02373__PTR198), .A2(_02148__PTR3), .ZN(_02374__PTR198) );
  AND2_X1 U13214 ( .A1(_02373__PTR199), .A2(_02148__PTR3), .ZN(_02374__PTR199) );
  AND2_X1 U13215 ( .A1(_02373__PTR200), .A2(_02148__PTR3), .ZN(_02374__PTR200) );
  AND2_X1 U13216 ( .A1(_02373__PTR201), .A2(_02148__PTR3), .ZN(_02374__PTR201) );
  AND2_X1 U13217 ( .A1(_02373__PTR202), .A2(_02148__PTR3), .ZN(_02374__PTR202) );
  AND2_X1 U13218 ( .A1(_02373__PTR203), .A2(_02148__PTR3), .ZN(_02374__PTR203) );
  AND2_X1 U13219 ( .A1(_02373__PTR204), .A2(_02148__PTR3), .ZN(_02374__PTR204) );
  AND2_X1 U13220 ( .A1(_02373__PTR205), .A2(_02148__PTR3), .ZN(_02374__PTR205) );
  AND2_X1 U13221 ( .A1(_02373__PTR206), .A2(_02148__PTR3), .ZN(_02374__PTR206) );
  AND2_X1 U13222 ( .A1(_02373__PTR207), .A2(_02148__PTR3), .ZN(_02374__PTR207) );
  AND2_X1 U13223 ( .A1(_02373__PTR208), .A2(_02148__PTR3), .ZN(_02374__PTR208) );
  AND2_X1 U13224 ( .A1(_02373__PTR209), .A2(_02148__PTR3), .ZN(_02374__PTR209) );
  AND2_X1 U13225 ( .A1(_02373__PTR210), .A2(_02148__PTR3), .ZN(_02374__PTR210) );
  AND2_X1 U13226 ( .A1(_02373__PTR211), .A2(_02148__PTR3), .ZN(_02374__PTR211) );
  AND2_X1 U13227 ( .A1(_02373__PTR212), .A2(_02148__PTR3), .ZN(_02374__PTR212) );
  AND2_X1 U13228 ( .A1(_02373__PTR213), .A2(_02148__PTR3), .ZN(_02374__PTR213) );
  AND2_X1 U13229 ( .A1(_02373__PTR214), .A2(_02148__PTR3), .ZN(_02374__PTR214) );
  AND2_X1 U13230 ( .A1(_02373__PTR215), .A2(_02148__PTR3), .ZN(_02374__PTR215) );
  AND2_X1 U13231 ( .A1(_02373__PTR216), .A2(_02148__PTR3), .ZN(_02374__PTR216) );
  AND2_X1 U13232 ( .A1(_02373__PTR217), .A2(_02148__PTR3), .ZN(_02374__PTR217) );
  AND2_X1 U13233 ( .A1(_02373__PTR218), .A2(_02148__PTR3), .ZN(_02374__PTR218) );
  AND2_X1 U13234 ( .A1(_02373__PTR219), .A2(_02148__PTR3), .ZN(_02374__PTR219) );
  AND2_X1 U13235 ( .A1(_02373__PTR220), .A2(_02148__PTR3), .ZN(_02374__PTR220) );
  AND2_X1 U13236 ( .A1(_02373__PTR221), .A2(_02148__PTR3), .ZN(_02374__PTR221) );
  AND2_X1 U13237 ( .A1(_02373__PTR222), .A2(_02148__PTR3), .ZN(_02374__PTR222) );
  AND2_X1 U13238 ( .A1(_02373__PTR223), .A2(_02148__PTR3), .ZN(_02374__PTR223) );
  AND2_X1 U13239 ( .A1(P2_P1_PhyAddrPointer_PTR0), .A2(_02383__PTR0), .ZN(_02382__PTR0) );
  AND2_X1 U13240 ( .A1(P2_P1_PhyAddrPointer_PTR1), .A2(_02383__PTR0), .ZN(_02382__PTR1) );
  AND2_X1 U13241 ( .A1(P2_P1_PhyAddrPointer_PTR2), .A2(_02383__PTR0), .ZN(_02382__PTR2) );
  AND2_X1 U13242 ( .A1(P2_P1_PhyAddrPointer_PTR3), .A2(_02383__PTR0), .ZN(_02382__PTR3) );
  AND2_X1 U13243 ( .A1(P2_P1_PhyAddrPointer_PTR4), .A2(_02383__PTR0), .ZN(_02382__PTR4) );
  AND2_X1 U13244 ( .A1(P2_P1_PhyAddrPointer_PTR5), .A2(_02383__PTR0), .ZN(_02382__PTR5) );
  AND2_X1 U13245 ( .A1(P2_P1_PhyAddrPointer_PTR6), .A2(_02383__PTR0), .ZN(_02382__PTR6) );
  AND2_X1 U13246 ( .A1(P2_P1_PhyAddrPointer_PTR7), .A2(_02383__PTR0), .ZN(_02382__PTR7) );
  AND2_X1 U13247 ( .A1(P2_P1_PhyAddrPointer_PTR8), .A2(_02383__PTR0), .ZN(_02382__PTR8) );
  AND2_X1 U13248 ( .A1(P2_P1_PhyAddrPointer_PTR9), .A2(_02383__PTR0), .ZN(_02382__PTR9) );
  AND2_X1 U13249 ( .A1(P2_P1_PhyAddrPointer_PTR10), .A2(_02383__PTR0), .ZN(_02382__PTR10) );
  AND2_X1 U13250 ( .A1(P2_P1_PhyAddrPointer_PTR11), .A2(_02383__PTR0), .ZN(_02382__PTR11) );
  AND2_X1 U13251 ( .A1(P2_P1_PhyAddrPointer_PTR12), .A2(_02383__PTR0), .ZN(_02382__PTR12) );
  AND2_X1 U13252 ( .A1(P2_P1_PhyAddrPointer_PTR13), .A2(_02383__PTR0), .ZN(_02382__PTR13) );
  AND2_X1 U13253 ( .A1(P2_P1_PhyAddrPointer_PTR14), .A2(_02383__PTR0), .ZN(_02382__PTR14) );
  AND2_X1 U13254 ( .A1(P2_P1_PhyAddrPointer_PTR15), .A2(_02383__PTR0), .ZN(_02382__PTR15) );
  AND2_X1 U13255 ( .A1(P2_P1_PhyAddrPointer_PTR16), .A2(_02383__PTR0), .ZN(_02382__PTR16) );
  AND2_X1 U13256 ( .A1(P2_P1_PhyAddrPointer_PTR17), .A2(_02383__PTR0), .ZN(_02382__PTR17) );
  AND2_X1 U13257 ( .A1(P2_P1_PhyAddrPointer_PTR18), .A2(_02383__PTR0), .ZN(_02382__PTR18) );
  AND2_X1 U13258 ( .A1(P2_P1_PhyAddrPointer_PTR19), .A2(_02383__PTR0), .ZN(_02382__PTR19) );
  AND2_X1 U13259 ( .A1(P2_P1_PhyAddrPointer_PTR20), .A2(_02383__PTR0), .ZN(_02382__PTR20) );
  AND2_X1 U13260 ( .A1(P2_P1_PhyAddrPointer_PTR21), .A2(_02383__PTR0), .ZN(_02382__PTR21) );
  AND2_X1 U13261 ( .A1(P2_P1_PhyAddrPointer_PTR22), .A2(_02383__PTR0), .ZN(_02382__PTR22) );
  AND2_X1 U13262 ( .A1(P2_P1_PhyAddrPointer_PTR23), .A2(_02383__PTR0), .ZN(_02382__PTR23) );
  AND2_X1 U13263 ( .A1(P2_P1_PhyAddrPointer_PTR24), .A2(_02383__PTR0), .ZN(_02382__PTR24) );
  AND2_X1 U13264 ( .A1(P2_P1_PhyAddrPointer_PTR25), .A2(_02383__PTR0), .ZN(_02382__PTR25) );
  AND2_X1 U13265 ( .A1(P2_P1_PhyAddrPointer_PTR26), .A2(_02383__PTR0), .ZN(_02382__PTR26) );
  AND2_X1 U13266 ( .A1(P2_P1_PhyAddrPointer_PTR27), .A2(_02383__PTR0), .ZN(_02382__PTR27) );
  AND2_X1 U13267 ( .A1(P2_P1_PhyAddrPointer_PTR28), .A2(_02383__PTR0), .ZN(_02382__PTR28) );
  AND2_X1 U13268 ( .A1(P2_P1_PhyAddrPointer_PTR29), .A2(_02383__PTR0), .ZN(_02382__PTR29) );
  AND2_X1 U13269 ( .A1(P2_P1_PhyAddrPointer_PTR30), .A2(_02383__PTR0), .ZN(_02382__PTR30) );
  AND2_X1 U13270 ( .A1(P2_P1_PhyAddrPointer_PTR31), .A2(_02383__PTR0), .ZN(_02382__PTR31) );
  AND2_X1 U13271 ( .A1(_02381__PTR32), .A2(_02148__PTR2), .ZN(_02382__PTR32) );
  AND2_X1 U13272 ( .A1(_02381__PTR33), .A2(_02148__PTR2), .ZN(_02382__PTR33) );
  AND2_X1 U13273 ( .A1(_02381__PTR34), .A2(_02148__PTR2), .ZN(_02382__PTR34) );
  AND2_X1 U13274 ( .A1(_02381__PTR35), .A2(_02148__PTR2), .ZN(_02382__PTR35) );
  AND2_X1 U13275 ( .A1(_02381__PTR36), .A2(_02148__PTR2), .ZN(_02382__PTR36) );
  AND2_X1 U13276 ( .A1(_02381__PTR37), .A2(_02148__PTR2), .ZN(_02382__PTR37) );
  AND2_X1 U13277 ( .A1(_02381__PTR38), .A2(_02148__PTR2), .ZN(_02382__PTR38) );
  AND2_X1 U13278 ( .A1(_02381__PTR39), .A2(_02148__PTR2), .ZN(_02382__PTR39) );
  AND2_X1 U13279 ( .A1(_02381__PTR40), .A2(_02148__PTR2), .ZN(_02382__PTR40) );
  AND2_X1 U13280 ( .A1(_02381__PTR41), .A2(_02148__PTR2), .ZN(_02382__PTR41) );
  AND2_X1 U13281 ( .A1(_02381__PTR42), .A2(_02148__PTR2), .ZN(_02382__PTR42) );
  AND2_X1 U13282 ( .A1(_02381__PTR43), .A2(_02148__PTR2), .ZN(_02382__PTR43) );
  AND2_X1 U13283 ( .A1(_02381__PTR44), .A2(_02148__PTR2), .ZN(_02382__PTR44) );
  AND2_X1 U13284 ( .A1(_02381__PTR45), .A2(_02148__PTR2), .ZN(_02382__PTR45) );
  AND2_X1 U13285 ( .A1(_02381__PTR46), .A2(_02148__PTR2), .ZN(_02382__PTR46) );
  AND2_X1 U13286 ( .A1(_02381__PTR47), .A2(_02148__PTR2), .ZN(_02382__PTR47) );
  AND2_X1 U13287 ( .A1(_02381__PTR48), .A2(_02148__PTR2), .ZN(_02382__PTR48) );
  AND2_X1 U13288 ( .A1(_02381__PTR49), .A2(_02148__PTR2), .ZN(_02382__PTR49) );
  AND2_X1 U13289 ( .A1(_02381__PTR50), .A2(_02148__PTR2), .ZN(_02382__PTR50) );
  AND2_X1 U13290 ( .A1(_02381__PTR51), .A2(_02148__PTR2), .ZN(_02382__PTR51) );
  AND2_X1 U13291 ( .A1(_02381__PTR52), .A2(_02148__PTR2), .ZN(_02382__PTR52) );
  AND2_X1 U13292 ( .A1(_02381__PTR53), .A2(_02148__PTR2), .ZN(_02382__PTR53) );
  AND2_X1 U13293 ( .A1(_02381__PTR54), .A2(_02148__PTR2), .ZN(_02382__PTR54) );
  AND2_X1 U13294 ( .A1(_02381__PTR55), .A2(_02148__PTR2), .ZN(_02382__PTR55) );
  AND2_X1 U13295 ( .A1(_02381__PTR56), .A2(_02148__PTR2), .ZN(_02382__PTR56) );
  AND2_X1 U13296 ( .A1(_02381__PTR57), .A2(_02148__PTR2), .ZN(_02382__PTR57) );
  AND2_X1 U13297 ( .A1(_02381__PTR58), .A2(_02148__PTR2), .ZN(_02382__PTR58) );
  AND2_X1 U13298 ( .A1(_02381__PTR59), .A2(_02148__PTR2), .ZN(_02382__PTR59) );
  AND2_X1 U13299 ( .A1(_02381__PTR60), .A2(_02148__PTR2), .ZN(_02382__PTR60) );
  AND2_X1 U13300 ( .A1(_02381__PTR61), .A2(_02148__PTR2), .ZN(_02382__PTR61) );
  AND2_X1 U13301 ( .A1(_02381__PTR62), .A2(_02148__PTR2), .ZN(_02382__PTR62) );
  AND2_X1 U13302 ( .A1(_02381__PTR63), .A2(_02148__PTR2), .ZN(_02382__PTR63) );
  AND2_X1 U13303 ( .A1(_02381__PTR64), .A2(_02148__PTR3), .ZN(_02382__PTR64) );
  AND2_X1 U13304 ( .A1(_02381__PTR65), .A2(_02148__PTR3), .ZN(_02382__PTR65) );
  AND2_X1 U13305 ( .A1(_02381__PTR66), .A2(_02148__PTR3), .ZN(_02382__PTR66) );
  AND2_X1 U13306 ( .A1(_02381__PTR67), .A2(_02148__PTR3), .ZN(_02382__PTR67) );
  AND2_X1 U13307 ( .A1(_02381__PTR68), .A2(_02148__PTR3), .ZN(_02382__PTR68) );
  AND2_X1 U13308 ( .A1(_02381__PTR69), .A2(_02148__PTR3), .ZN(_02382__PTR69) );
  AND2_X1 U13309 ( .A1(_02381__PTR70), .A2(_02148__PTR3), .ZN(_02382__PTR70) );
  AND2_X1 U13310 ( .A1(_02381__PTR71), .A2(_02148__PTR3), .ZN(_02382__PTR71) );
  AND2_X1 U13311 ( .A1(_02381__PTR72), .A2(_02148__PTR3), .ZN(_02382__PTR72) );
  AND2_X1 U13312 ( .A1(_02381__PTR73), .A2(_02148__PTR3), .ZN(_02382__PTR73) );
  AND2_X1 U13313 ( .A1(_02381__PTR74), .A2(_02148__PTR3), .ZN(_02382__PTR74) );
  AND2_X1 U13314 ( .A1(_02381__PTR75), .A2(_02148__PTR3), .ZN(_02382__PTR75) );
  AND2_X1 U13315 ( .A1(_02381__PTR76), .A2(_02148__PTR3), .ZN(_02382__PTR76) );
  AND2_X1 U13316 ( .A1(_02381__PTR77), .A2(_02148__PTR3), .ZN(_02382__PTR77) );
  AND2_X1 U13317 ( .A1(_02381__PTR78), .A2(_02148__PTR3), .ZN(_02382__PTR78) );
  AND2_X1 U13318 ( .A1(_02381__PTR79), .A2(_02148__PTR3), .ZN(_02382__PTR79) );
  AND2_X1 U13319 ( .A1(_02381__PTR80), .A2(_02148__PTR3), .ZN(_02382__PTR80) );
  AND2_X1 U13320 ( .A1(_02381__PTR81), .A2(_02148__PTR3), .ZN(_02382__PTR81) );
  AND2_X1 U13321 ( .A1(_02381__PTR82), .A2(_02148__PTR3), .ZN(_02382__PTR82) );
  AND2_X1 U13322 ( .A1(_02381__PTR83), .A2(_02148__PTR3), .ZN(_02382__PTR83) );
  AND2_X1 U13323 ( .A1(_02381__PTR84), .A2(_02148__PTR3), .ZN(_02382__PTR84) );
  AND2_X1 U13324 ( .A1(_02381__PTR85), .A2(_02148__PTR3), .ZN(_02382__PTR85) );
  AND2_X1 U13325 ( .A1(_02381__PTR86), .A2(_02148__PTR3), .ZN(_02382__PTR86) );
  AND2_X1 U13326 ( .A1(_02381__PTR87), .A2(_02148__PTR3), .ZN(_02382__PTR87) );
  AND2_X1 U13327 ( .A1(_02381__PTR88), .A2(_02148__PTR3), .ZN(_02382__PTR88) );
  AND2_X1 U13328 ( .A1(_02381__PTR89), .A2(_02148__PTR3), .ZN(_02382__PTR89) );
  AND2_X1 U13329 ( .A1(_02381__PTR90), .A2(_02148__PTR3), .ZN(_02382__PTR90) );
  AND2_X1 U13330 ( .A1(_02381__PTR91), .A2(_02148__PTR3), .ZN(_02382__PTR91) );
  AND2_X1 U13331 ( .A1(_02381__PTR92), .A2(_02148__PTR3), .ZN(_02382__PTR92) );
  AND2_X1 U13332 ( .A1(_02381__PTR93), .A2(_02148__PTR3), .ZN(_02382__PTR93) );
  AND2_X1 U13333 ( .A1(_02381__PTR94), .A2(_02148__PTR3), .ZN(_02382__PTR94) );
  AND2_X1 U13334 ( .A1(_02381__PTR95), .A2(_02148__PTR3), .ZN(_02382__PTR95) );
  AND2_X1 U13335 ( .A1(P2_P1_State2_PTR0), .A2(_02409__PTR0), .ZN(_02408__PTR0) );
  AND2_X1 U13336 ( .A1(P2_P1_State2_PTR1), .A2(_02409__PTR0), .ZN(_02408__PTR1) );
  AND2_X1 U13337 ( .A1(P2_P1_State2_PTR2), .A2(_02409__PTR0), .ZN(_02408__PTR2) );
  AND2_X1 U13338 ( .A1(P2_P1_State2_PTR3), .A2(_02409__PTR0), .ZN(_02408__PTR3) );
  AND2_X1 U13339 ( .A1(_02407__PTR4), .A2(_02156__PTR2), .ZN(_02408__PTR4) );
  AND2_X1 U13340 ( .A1(_02407__PTR5), .A2(_02156__PTR2), .ZN(_02408__PTR5) );
  AND2_X1 U13341 ( .A1(_02407__PTR6), .A2(_02156__PTR2), .ZN(_02408__PTR6) );
  AND2_X1 U13342 ( .A1(_02407__PTR7), .A2(_02156__PTR2), .ZN(_02408__PTR7) );
  AND2_X1 U13343 ( .A1(_02463__PTR8), .A2(_02702__PTR1), .ZN(_02701__PTR4) );
  AND2_X1 U13344 ( .A1(P3_rEIP_PTR1), .A2(_02702__PTR1), .ZN(_02701__PTR5) );
  AND2_X1 U13345 ( .A1(_02463__PTR2), .A2(_02702__PTR1), .ZN(_02701__PTR6) );
  AND2_X1 U13346 ( .A1(_02463__PTR8), .A2(_02702__PTR2), .ZN(_02701__PTR8) );
  AND2_X1 U13347 ( .A1(P3_rEIP_PTR1), .A2(_02702__PTR2), .ZN(_02701__PTR9) );
  AND2_X1 U13348 ( .A1(_02463__PTR6), .A2(_02702__PTR2), .ZN(_02701__PTR10) );
  AND2_X1 U13349 ( .A1(_02463__PTR7), .A2(_02702__PTR2), .ZN(_02701__PTR11) );
  AND2_X1 U13350 ( .A1(_02463__PTR8), .A2(_02702__PTR3), .ZN(_02701__PTR12) );
  AND2_X1 U13351 ( .A1(_02463__PTR9), .A2(_02702__PTR3), .ZN(_02701__PTR13) );
  AND2_X1 U13352 ( .A1(_02463__PTR10), .A2(_02702__PTR3), .ZN(_02701__PTR14) );
  AND2_X1 U13353 ( .A1(_02463__PTR11), .A2(_02702__PTR3), .ZN(_02701__PTR15) );
  AND2_X1 U13354 ( .A1(P3_Datao_PTR0), .A2(_02694__PTR0), .ZN(_02693__PTR0) );
  AND2_X1 U13355 ( .A1(P3_Datao_PTR1), .A2(_02694__PTR0), .ZN(_02693__PTR1) );
  AND2_X1 U13356 ( .A1(P3_Datao_PTR2), .A2(_02694__PTR0), .ZN(_02693__PTR2) );
  AND2_X1 U13357 ( .A1(P3_Datao_PTR3), .A2(_02694__PTR0), .ZN(_02693__PTR3) );
  AND2_X1 U13358 ( .A1(P3_Datao_PTR4), .A2(_02694__PTR0), .ZN(_02693__PTR4) );
  AND2_X1 U13359 ( .A1(P3_Datao_PTR5), .A2(_02694__PTR0), .ZN(_02693__PTR5) );
  AND2_X1 U13360 ( .A1(P3_Datao_PTR6), .A2(_02694__PTR0), .ZN(_02693__PTR6) );
  AND2_X1 U13361 ( .A1(P3_Datao_PTR7), .A2(_02694__PTR0), .ZN(_02693__PTR7) );
  AND2_X1 U13362 ( .A1(P3_Datao_PTR8), .A2(_02694__PTR0), .ZN(_02693__PTR8) );
  AND2_X1 U13363 ( .A1(P3_Datao_PTR9), .A2(_02694__PTR0), .ZN(_02693__PTR9) );
  AND2_X1 U13364 ( .A1(P3_Datao_PTR10), .A2(_02694__PTR0), .ZN(_02693__PTR10) );
  AND2_X1 U13365 ( .A1(P3_Datao_PTR11), .A2(_02694__PTR0), .ZN(_02693__PTR11) );
  AND2_X1 U13366 ( .A1(P3_Datao_PTR12), .A2(_02694__PTR0), .ZN(_02693__PTR12) );
  AND2_X1 U13367 ( .A1(P3_Datao_PTR13), .A2(_02694__PTR0), .ZN(_02693__PTR13) );
  AND2_X1 U13368 ( .A1(P3_Datao_PTR14), .A2(_02694__PTR0), .ZN(_02693__PTR14) );
  AND2_X1 U13369 ( .A1(P3_Datao_PTR15), .A2(_02694__PTR0), .ZN(_02693__PTR15) );
  AND2_X1 U13370 ( .A1(P3_Datao_PTR16), .A2(_02694__PTR0), .ZN(_02693__PTR16) );
  AND2_X1 U13371 ( .A1(P3_Datao_PTR17), .A2(_02694__PTR0), .ZN(_02693__PTR17) );
  AND2_X1 U13372 ( .A1(P3_Datao_PTR18), .A2(_02694__PTR0), .ZN(_02693__PTR18) );
  AND2_X1 U13373 ( .A1(P3_Datao_PTR19), .A2(_02694__PTR0), .ZN(_02693__PTR19) );
  AND2_X1 U13374 ( .A1(P3_Datao_PTR20), .A2(_02694__PTR0), .ZN(_02693__PTR20) );
  AND2_X1 U13375 ( .A1(P3_Datao_PTR21), .A2(_02694__PTR0), .ZN(_02693__PTR21) );
  AND2_X1 U13376 ( .A1(P3_Datao_PTR22), .A2(_02694__PTR0), .ZN(_02693__PTR22) );
  AND2_X1 U13377 ( .A1(P3_Datao_PTR23), .A2(_02694__PTR0), .ZN(_02693__PTR23) );
  AND2_X1 U13378 ( .A1(P3_Datao_PTR24), .A2(_02694__PTR0), .ZN(_02693__PTR24) );
  AND2_X1 U13379 ( .A1(P3_Datao_PTR25), .A2(_02694__PTR0), .ZN(_02693__PTR25) );
  AND2_X1 U13380 ( .A1(P3_Datao_PTR26), .A2(_02694__PTR0), .ZN(_02693__PTR26) );
  AND2_X1 U13381 ( .A1(P3_Datao_PTR27), .A2(_02694__PTR0), .ZN(_02693__PTR27) );
  AND2_X1 U13382 ( .A1(P3_Datao_PTR28), .A2(_02694__PTR0), .ZN(_02693__PTR28) );
  AND2_X1 U13383 ( .A1(P3_Datao_PTR29), .A2(_02694__PTR0), .ZN(_02693__PTR29) );
  AND2_X1 U13384 ( .A1(P3_Datao_PTR30), .A2(_02694__PTR0), .ZN(_02693__PTR30) );
  AND2_X1 U13385 ( .A1(P3_Datao_PTR31), .A2(_02694__PTR0), .ZN(_02693__PTR31) );
  AND2_X1 U13386 ( .A1(_02692__PTR64), .A2(_02445__PTR0), .ZN(_02693__PTR32) );
  AND2_X1 U13387 ( .A1(_02692__PTR65), .A2(_02445__PTR0), .ZN(_02693__PTR33) );
  AND2_X1 U13388 ( .A1(_02692__PTR66), .A2(_02445__PTR0), .ZN(_02693__PTR34) );
  AND2_X1 U13389 ( .A1(_02692__PTR67), .A2(_02445__PTR0), .ZN(_02693__PTR35) );
  AND2_X1 U13390 ( .A1(_02692__PTR68), .A2(_02445__PTR0), .ZN(_02693__PTR36) );
  AND2_X1 U13391 ( .A1(_02692__PTR69), .A2(_02445__PTR0), .ZN(_02693__PTR37) );
  AND2_X1 U13392 ( .A1(_02692__PTR70), .A2(_02445__PTR0), .ZN(_02693__PTR38) );
  AND2_X1 U13393 ( .A1(_02692__PTR71), .A2(_02445__PTR0), .ZN(_02693__PTR39) );
  AND2_X1 U13394 ( .A1(_02692__PTR72), .A2(_02445__PTR0), .ZN(_02693__PTR40) );
  AND2_X1 U13395 ( .A1(_02692__PTR73), .A2(_02445__PTR0), .ZN(_02693__PTR41) );
  AND2_X1 U13396 ( .A1(_02692__PTR74), .A2(_02445__PTR0), .ZN(_02693__PTR42) );
  AND2_X1 U13397 ( .A1(_02692__PTR75), .A2(_02445__PTR0), .ZN(_02693__PTR43) );
  AND2_X1 U13398 ( .A1(_02692__PTR76), .A2(_02445__PTR0), .ZN(_02693__PTR44) );
  AND2_X1 U13399 ( .A1(_02692__PTR77), .A2(_02445__PTR0), .ZN(_02693__PTR45) );
  AND2_X1 U13400 ( .A1(_02692__PTR78), .A2(_02445__PTR0), .ZN(_02693__PTR46) );
  AND2_X1 U13401 ( .A1(_02692__PTR79), .A2(_02445__PTR0), .ZN(_02693__PTR47) );
  AND2_X1 U13402 ( .A1(_02692__PTR48), .A2(_02445__PTR0), .ZN(_02693__PTR48) );
  AND2_X1 U13403 ( .A1(_02692__PTR49), .A2(_02445__PTR0), .ZN(_02693__PTR49) );
  AND2_X1 U13404 ( .A1(_02692__PTR50), .A2(_02445__PTR0), .ZN(_02693__PTR50) );
  AND2_X1 U13405 ( .A1(_02692__PTR51), .A2(_02445__PTR0), .ZN(_02693__PTR51) );
  AND2_X1 U13406 ( .A1(_02692__PTR52), .A2(_02445__PTR0), .ZN(_02693__PTR52) );
  AND2_X1 U13407 ( .A1(_02692__PTR53), .A2(_02445__PTR0), .ZN(_02693__PTR53) );
  AND2_X1 U13408 ( .A1(_02692__PTR54), .A2(_02445__PTR0), .ZN(_02693__PTR54) );
  AND2_X1 U13409 ( .A1(_02692__PTR55), .A2(_02445__PTR0), .ZN(_02693__PTR55) );
  AND2_X1 U13410 ( .A1(_02692__PTR56), .A2(_02445__PTR0), .ZN(_02693__PTR56) );
  AND2_X1 U13411 ( .A1(_02692__PTR57), .A2(_02445__PTR0), .ZN(_02693__PTR57) );
  AND2_X1 U13412 ( .A1(_02692__PTR58), .A2(_02445__PTR0), .ZN(_02693__PTR58) );
  AND2_X1 U13413 ( .A1(_02692__PTR59), .A2(_02445__PTR0), .ZN(_02693__PTR59) );
  AND2_X1 U13414 ( .A1(_02692__PTR60), .A2(_02445__PTR0), .ZN(_02693__PTR60) );
  AND2_X1 U13415 ( .A1(_02692__PTR61), .A2(_02445__PTR0), .ZN(_02693__PTR61) );
  AND2_X1 U13416 ( .A1(_02692__PTR62), .A2(_02445__PTR0), .ZN(_02693__PTR62) );
  AND2_X1 U13417 ( .A1(_02692__PTR95), .A2(_02445__PTR0), .ZN(_02693__PTR63) );
  AND2_X1 U13418 ( .A1(_02692__PTR64), .A2(_02445__PTR2), .ZN(_02693__PTR64) );
  AND2_X1 U13419 ( .A1(_02692__PTR65), .A2(_02445__PTR2), .ZN(_02693__PTR65) );
  AND2_X1 U13420 ( .A1(_02692__PTR66), .A2(_02445__PTR2), .ZN(_02693__PTR66) );
  AND2_X1 U13421 ( .A1(_02692__PTR67), .A2(_02445__PTR2), .ZN(_02693__PTR67) );
  AND2_X1 U13422 ( .A1(_02692__PTR68), .A2(_02445__PTR2), .ZN(_02693__PTR68) );
  AND2_X1 U13423 ( .A1(_02692__PTR69), .A2(_02445__PTR2), .ZN(_02693__PTR69) );
  AND2_X1 U13424 ( .A1(_02692__PTR70), .A2(_02445__PTR2), .ZN(_02693__PTR70) );
  AND2_X1 U13425 ( .A1(_02692__PTR71), .A2(_02445__PTR2), .ZN(_02693__PTR71) );
  AND2_X1 U13426 ( .A1(_02692__PTR72), .A2(_02445__PTR2), .ZN(_02693__PTR72) );
  AND2_X1 U13427 ( .A1(_02692__PTR73), .A2(_02445__PTR2), .ZN(_02693__PTR73) );
  AND2_X1 U13428 ( .A1(_02692__PTR74), .A2(_02445__PTR2), .ZN(_02693__PTR74) );
  AND2_X1 U13429 ( .A1(_02692__PTR75), .A2(_02445__PTR2), .ZN(_02693__PTR75) );
  AND2_X1 U13430 ( .A1(_02692__PTR76), .A2(_02445__PTR2), .ZN(_02693__PTR76) );
  AND2_X1 U13431 ( .A1(_02692__PTR77), .A2(_02445__PTR2), .ZN(_02693__PTR77) );
  AND2_X1 U13432 ( .A1(_02692__PTR78), .A2(_02445__PTR2), .ZN(_02693__PTR78) );
  AND2_X1 U13433 ( .A1(_02692__PTR79), .A2(_02445__PTR2), .ZN(_02693__PTR79) );
  AND2_X1 U13434 ( .A1(_02692__PTR80), .A2(_02445__PTR2), .ZN(_02693__PTR80) );
  AND2_X1 U13435 ( .A1(_02692__PTR81), .A2(_02445__PTR2), .ZN(_02693__PTR81) );
  AND2_X1 U13436 ( .A1(_02692__PTR82), .A2(_02445__PTR2), .ZN(_02693__PTR82) );
  AND2_X1 U13437 ( .A1(_02692__PTR83), .A2(_02445__PTR2), .ZN(_02693__PTR83) );
  AND2_X1 U13438 ( .A1(_02692__PTR84), .A2(_02445__PTR2), .ZN(_02693__PTR84) );
  AND2_X1 U13439 ( .A1(_02692__PTR85), .A2(_02445__PTR2), .ZN(_02693__PTR85) );
  AND2_X1 U13440 ( .A1(_02692__PTR86), .A2(_02445__PTR2), .ZN(_02693__PTR86) );
  AND2_X1 U13441 ( .A1(_02692__PTR87), .A2(_02445__PTR2), .ZN(_02693__PTR87) );
  AND2_X1 U13442 ( .A1(_02692__PTR88), .A2(_02445__PTR2), .ZN(_02693__PTR88) );
  AND2_X1 U13443 ( .A1(_02692__PTR89), .A2(_02445__PTR2), .ZN(_02693__PTR89) );
  AND2_X1 U13444 ( .A1(_02692__PTR90), .A2(_02445__PTR2), .ZN(_02693__PTR90) );
  AND2_X1 U13445 ( .A1(_02692__PTR91), .A2(_02445__PTR2), .ZN(_02693__PTR91) );
  AND2_X1 U13446 ( .A1(_02692__PTR92), .A2(_02445__PTR2), .ZN(_02693__PTR92) );
  AND2_X1 U13447 ( .A1(_02692__PTR93), .A2(_02445__PTR2), .ZN(_02693__PTR93) );
  AND2_X1 U13448 ( .A1(_02692__PTR94), .A2(_02445__PTR2), .ZN(_02693__PTR94) );
  AND2_X1 U13449 ( .A1(_02692__PTR95), .A2(_02445__PTR2), .ZN(_02693__PTR95) );
  AND2_X1 U13450 ( .A1(P3_P1_lWord_PTR0), .A2(_02687__PTR0), .ZN(_02690__PTR0) );
  AND2_X1 U13451 ( .A1(P3_P1_lWord_PTR1), .A2(_02687__PTR0), .ZN(_02690__PTR1) );
  AND2_X1 U13452 ( .A1(P3_P1_lWord_PTR2), .A2(_02687__PTR0), .ZN(_02690__PTR2) );
  AND2_X1 U13453 ( .A1(P3_P1_lWord_PTR3), .A2(_02687__PTR0), .ZN(_02690__PTR3) );
  AND2_X1 U13454 ( .A1(P3_P1_lWord_PTR4), .A2(_02687__PTR0), .ZN(_02690__PTR4) );
  AND2_X1 U13455 ( .A1(P3_P1_lWord_PTR5), .A2(_02687__PTR0), .ZN(_02690__PTR5) );
  AND2_X1 U13456 ( .A1(P3_P1_lWord_PTR6), .A2(_02687__PTR0), .ZN(_02690__PTR6) );
  AND2_X1 U13457 ( .A1(P3_P1_lWord_PTR7), .A2(_02687__PTR0), .ZN(_02690__PTR7) );
  AND2_X1 U13458 ( .A1(P3_P1_lWord_PTR8), .A2(_02687__PTR0), .ZN(_02690__PTR8) );
  AND2_X1 U13459 ( .A1(P3_P1_lWord_PTR9), .A2(_02687__PTR0), .ZN(_02690__PTR9) );
  AND2_X1 U13460 ( .A1(P3_P1_lWord_PTR10), .A2(_02687__PTR0), .ZN(_02690__PTR10) );
  AND2_X1 U13461 ( .A1(P3_P1_lWord_PTR11), .A2(_02687__PTR0), .ZN(_02690__PTR11) );
  AND2_X1 U13462 ( .A1(P3_P1_lWord_PTR12), .A2(_02687__PTR0), .ZN(_02690__PTR12) );
  AND2_X1 U13463 ( .A1(P3_P1_lWord_PTR13), .A2(_02687__PTR0), .ZN(_02690__PTR13) );
  AND2_X1 U13464 ( .A1(P3_P1_lWord_PTR14), .A2(_02687__PTR0), .ZN(_02690__PTR14) );
  AND2_X1 U13465 ( .A1(P3_P1_lWord_PTR15), .A2(_02687__PTR0), .ZN(_02690__PTR15) );
  AND2_X1 U13466 ( .A1(_02689__PTR16), .A2(_02445__PTR2), .ZN(_02690__PTR16) );
  AND2_X1 U13467 ( .A1(_02689__PTR17), .A2(_02445__PTR2), .ZN(_02690__PTR17) );
  AND2_X1 U13468 ( .A1(_02689__PTR18), .A2(_02445__PTR2), .ZN(_02690__PTR18) );
  AND2_X1 U13469 ( .A1(_02689__PTR19), .A2(_02445__PTR2), .ZN(_02690__PTR19) );
  AND2_X1 U13470 ( .A1(_02689__PTR20), .A2(_02445__PTR2), .ZN(_02690__PTR20) );
  AND2_X1 U13471 ( .A1(_02689__PTR21), .A2(_02445__PTR2), .ZN(_02690__PTR21) );
  AND2_X1 U13472 ( .A1(_02689__PTR22), .A2(_02445__PTR2), .ZN(_02690__PTR22) );
  AND2_X1 U13473 ( .A1(_02689__PTR23), .A2(_02445__PTR2), .ZN(_02690__PTR23) );
  AND2_X1 U13474 ( .A1(_02689__PTR24), .A2(_02445__PTR2), .ZN(_02690__PTR24) );
  AND2_X1 U13475 ( .A1(_02689__PTR25), .A2(_02445__PTR2), .ZN(_02690__PTR25) );
  AND2_X1 U13476 ( .A1(_02689__PTR26), .A2(_02445__PTR2), .ZN(_02690__PTR26) );
  AND2_X1 U13477 ( .A1(_02689__PTR27), .A2(_02445__PTR2), .ZN(_02690__PTR27) );
  AND2_X1 U13478 ( .A1(_02689__PTR28), .A2(_02445__PTR2), .ZN(_02690__PTR28) );
  AND2_X1 U13479 ( .A1(_02689__PTR29), .A2(_02445__PTR2), .ZN(_02690__PTR29) );
  AND2_X1 U13480 ( .A1(_02689__PTR30), .A2(_02445__PTR2), .ZN(_02690__PTR30) );
  AND2_X1 U13481 ( .A1(_02689__PTR31), .A2(_02445__PTR2), .ZN(_02690__PTR31) );
  AND2_X1 U13482 ( .A1(_02689__PTR32), .A2(_02668__PTR4), .ZN(_02690__PTR32) );
  AND2_X1 U13483 ( .A1(_02689__PTR33), .A2(_02668__PTR4), .ZN(_02690__PTR33) );
  AND2_X1 U13484 ( .A1(_02689__PTR34), .A2(_02668__PTR4), .ZN(_02690__PTR34) );
  AND2_X1 U13485 ( .A1(_02689__PTR35), .A2(_02668__PTR4), .ZN(_02690__PTR35) );
  AND2_X1 U13486 ( .A1(_02689__PTR36), .A2(_02668__PTR4), .ZN(_02690__PTR36) );
  AND2_X1 U13487 ( .A1(_02689__PTR37), .A2(_02668__PTR4), .ZN(_02690__PTR37) );
  AND2_X1 U13488 ( .A1(_02689__PTR38), .A2(_02668__PTR4), .ZN(_02690__PTR38) );
  AND2_X1 U13489 ( .A1(_02689__PTR39), .A2(_02668__PTR4), .ZN(_02690__PTR39) );
  AND2_X1 U13490 ( .A1(_02689__PTR40), .A2(_02668__PTR4), .ZN(_02690__PTR40) );
  AND2_X1 U13491 ( .A1(_02689__PTR41), .A2(_02668__PTR4), .ZN(_02690__PTR41) );
  AND2_X1 U13492 ( .A1(_02689__PTR42), .A2(_02668__PTR4), .ZN(_02690__PTR42) );
  AND2_X1 U13493 ( .A1(_02689__PTR43), .A2(_02668__PTR4), .ZN(_02690__PTR43) );
  AND2_X1 U13494 ( .A1(_02689__PTR44), .A2(_02668__PTR4), .ZN(_02690__PTR44) );
  AND2_X1 U13495 ( .A1(_02689__PTR45), .A2(_02668__PTR4), .ZN(_02690__PTR45) );
  AND2_X1 U13496 ( .A1(_02689__PTR46), .A2(_02668__PTR4), .ZN(_02690__PTR46) );
  AND2_X1 U13497 ( .A1(_02689__PTR47), .A2(_02668__PTR4), .ZN(_02690__PTR47) );
  AND2_X1 U13498 ( .A1(P3_P1_uWord_PTR0), .A2(_02687__PTR0), .ZN(_02686__PTR0) );
  AND2_X1 U13499 ( .A1(P3_P1_uWord_PTR1), .A2(_02687__PTR0), .ZN(_02686__PTR1) );
  AND2_X1 U13500 ( .A1(P3_P1_uWord_PTR2), .A2(_02687__PTR0), .ZN(_02686__PTR2) );
  AND2_X1 U13501 ( .A1(P3_P1_uWord_PTR3), .A2(_02687__PTR0), .ZN(_02686__PTR3) );
  AND2_X1 U13502 ( .A1(P3_P1_uWord_PTR4), .A2(_02687__PTR0), .ZN(_02686__PTR4) );
  AND2_X1 U13503 ( .A1(P3_P1_uWord_PTR5), .A2(_02687__PTR0), .ZN(_02686__PTR5) );
  AND2_X1 U13504 ( .A1(P3_P1_uWord_PTR6), .A2(_02687__PTR0), .ZN(_02686__PTR6) );
  AND2_X1 U13505 ( .A1(P3_P1_uWord_PTR7), .A2(_02687__PTR0), .ZN(_02686__PTR7) );
  AND2_X1 U13506 ( .A1(P3_P1_uWord_PTR8), .A2(_02687__PTR0), .ZN(_02686__PTR8) );
  AND2_X1 U13507 ( .A1(P3_P1_uWord_PTR9), .A2(_02687__PTR0), .ZN(_02686__PTR9) );
  AND2_X1 U13508 ( .A1(P3_P1_uWord_PTR10), .A2(_02687__PTR0), .ZN(_02686__PTR10) );
  AND2_X1 U13509 ( .A1(P3_P1_uWord_PTR11), .A2(_02687__PTR0), .ZN(_02686__PTR11) );
  AND2_X1 U13510 ( .A1(P3_P1_uWord_PTR12), .A2(_02687__PTR0), .ZN(_02686__PTR12) );
  AND2_X1 U13511 ( .A1(P3_P1_uWord_PTR13), .A2(_02687__PTR0), .ZN(_02686__PTR13) );
  AND2_X1 U13512 ( .A1(P3_P1_uWord_PTR14), .A2(_02687__PTR0), .ZN(_02686__PTR14) );
  AND2_X1 U13513 ( .A1(_02685__PTR15), .A2(_02445__PTR2), .ZN(_02686__PTR15) );
  AND2_X1 U13514 ( .A1(_02685__PTR16), .A2(_02445__PTR2), .ZN(_02686__PTR16) );
  AND2_X1 U13515 ( .A1(_02685__PTR17), .A2(_02445__PTR2), .ZN(_02686__PTR17) );
  AND2_X1 U13516 ( .A1(_02685__PTR18), .A2(_02445__PTR2), .ZN(_02686__PTR18) );
  AND2_X1 U13517 ( .A1(_02685__PTR19), .A2(_02445__PTR2), .ZN(_02686__PTR19) );
  AND2_X1 U13518 ( .A1(_02685__PTR20), .A2(_02445__PTR2), .ZN(_02686__PTR20) );
  AND2_X1 U13519 ( .A1(_02685__PTR21), .A2(_02445__PTR2), .ZN(_02686__PTR21) );
  AND2_X1 U13520 ( .A1(_02685__PTR22), .A2(_02445__PTR2), .ZN(_02686__PTR22) );
  AND2_X1 U13521 ( .A1(_02685__PTR23), .A2(_02445__PTR2), .ZN(_02686__PTR23) );
  AND2_X1 U13522 ( .A1(_02685__PTR24), .A2(_02445__PTR2), .ZN(_02686__PTR24) );
  AND2_X1 U13523 ( .A1(_02685__PTR25), .A2(_02445__PTR2), .ZN(_02686__PTR25) );
  AND2_X1 U13524 ( .A1(_02685__PTR26), .A2(_02445__PTR2), .ZN(_02686__PTR26) );
  AND2_X1 U13525 ( .A1(_02685__PTR27), .A2(_02445__PTR2), .ZN(_02686__PTR27) );
  AND2_X1 U13526 ( .A1(_02685__PTR28), .A2(_02445__PTR2), .ZN(_02686__PTR28) );
  AND2_X1 U13527 ( .A1(_02685__PTR29), .A2(_02445__PTR2), .ZN(_02686__PTR29) );
  AND2_X1 U13528 ( .A1(_02685__PTR30), .A2(_02668__PTR4), .ZN(_02686__PTR30) );
  AND2_X1 U13529 ( .A1(_02685__PTR31), .A2(_02668__PTR4), .ZN(_02686__PTR31) );
  AND2_X1 U13530 ( .A1(_02685__PTR32), .A2(_02668__PTR4), .ZN(_02686__PTR32) );
  AND2_X1 U13531 ( .A1(_02685__PTR33), .A2(_02668__PTR4), .ZN(_02686__PTR33) );
  AND2_X1 U13532 ( .A1(_02685__PTR34), .A2(_02668__PTR4), .ZN(_02686__PTR34) );
  AND2_X1 U13533 ( .A1(_02685__PTR35), .A2(_02668__PTR4), .ZN(_02686__PTR35) );
  AND2_X1 U13534 ( .A1(_02685__PTR36), .A2(_02668__PTR4), .ZN(_02686__PTR36) );
  AND2_X1 U13535 ( .A1(_02685__PTR37), .A2(_02668__PTR4), .ZN(_02686__PTR37) );
  AND2_X1 U13536 ( .A1(_02685__PTR38), .A2(_02668__PTR4), .ZN(_02686__PTR38) );
  AND2_X1 U13537 ( .A1(_02685__PTR39), .A2(_02668__PTR4), .ZN(_02686__PTR39) );
  AND2_X1 U13538 ( .A1(_02685__PTR40), .A2(_02668__PTR4), .ZN(_02686__PTR40) );
  AND2_X1 U13539 ( .A1(_02685__PTR41), .A2(_02668__PTR4), .ZN(_02686__PTR41) );
  AND2_X1 U13540 ( .A1(_02685__PTR42), .A2(_02668__PTR4), .ZN(_02686__PTR42) );
  AND2_X1 U13541 ( .A1(_02685__PTR43), .A2(_02668__PTR4), .ZN(_02686__PTR43) );
  AND2_X1 U13542 ( .A1(_02685__PTR44), .A2(_02668__PTR4), .ZN(_02686__PTR44) );
  AND2_X1 U13543 ( .A1(P3_EBX_PTR0), .A2(_02680__PTR0), .ZN(_02679__PTR0) );
  AND2_X1 U13544 ( .A1(P3_EBX_PTR1), .A2(_02680__PTR0), .ZN(_02679__PTR1) );
  AND2_X1 U13545 ( .A1(P3_EBX_PTR2), .A2(_02680__PTR0), .ZN(_02679__PTR2) );
  AND2_X1 U13546 ( .A1(P3_EBX_PTR3), .A2(_02680__PTR0), .ZN(_02679__PTR3) );
  AND2_X1 U13547 ( .A1(P3_EBX_PTR4), .A2(_02680__PTR0), .ZN(_02679__PTR4) );
  AND2_X1 U13548 ( .A1(P3_EBX_PTR5), .A2(_02680__PTR0), .ZN(_02679__PTR5) );
  AND2_X1 U13549 ( .A1(P3_EBX_PTR6), .A2(_02680__PTR0), .ZN(_02679__PTR6) );
  AND2_X1 U13550 ( .A1(P3_EBX_PTR7), .A2(_02680__PTR0), .ZN(_02679__PTR7) );
  AND2_X1 U13551 ( .A1(P3_EBX_PTR8), .A2(_02680__PTR0), .ZN(_02679__PTR8) );
  AND2_X1 U13552 ( .A1(P3_EBX_PTR9), .A2(_02680__PTR0), .ZN(_02679__PTR9) );
  AND2_X1 U13553 ( .A1(P3_EBX_PTR10), .A2(_02680__PTR0), .ZN(_02679__PTR10) );
  AND2_X1 U13554 ( .A1(P3_EBX_PTR11), .A2(_02680__PTR0), .ZN(_02679__PTR11) );
  AND2_X1 U13555 ( .A1(P3_EBX_PTR12), .A2(_02680__PTR0), .ZN(_02679__PTR12) );
  AND2_X1 U13556 ( .A1(P3_EBX_PTR13), .A2(_02680__PTR0), .ZN(_02679__PTR13) );
  AND2_X1 U13557 ( .A1(P3_EBX_PTR14), .A2(_02680__PTR0), .ZN(_02679__PTR14) );
  AND2_X1 U13558 ( .A1(P3_EBX_PTR15), .A2(_02680__PTR0), .ZN(_02679__PTR15) );
  AND2_X1 U13559 ( .A1(P3_EBX_PTR16), .A2(_02680__PTR0), .ZN(_02679__PTR16) );
  AND2_X1 U13560 ( .A1(P3_EBX_PTR17), .A2(_02680__PTR0), .ZN(_02679__PTR17) );
  AND2_X1 U13561 ( .A1(P3_EBX_PTR18), .A2(_02680__PTR0), .ZN(_02679__PTR18) );
  AND2_X1 U13562 ( .A1(P3_EBX_PTR19), .A2(_02680__PTR0), .ZN(_02679__PTR19) );
  AND2_X1 U13563 ( .A1(P3_EBX_PTR20), .A2(_02680__PTR0), .ZN(_02679__PTR20) );
  AND2_X1 U13564 ( .A1(P3_EBX_PTR21), .A2(_02680__PTR0), .ZN(_02679__PTR21) );
  AND2_X1 U13565 ( .A1(P3_EBX_PTR22), .A2(_02680__PTR0), .ZN(_02679__PTR22) );
  AND2_X1 U13566 ( .A1(P3_EBX_PTR23), .A2(_02680__PTR0), .ZN(_02679__PTR23) );
  AND2_X1 U13567 ( .A1(P3_EBX_PTR24), .A2(_02680__PTR0), .ZN(_02679__PTR24) );
  AND2_X1 U13568 ( .A1(P3_EBX_PTR25), .A2(_02680__PTR0), .ZN(_02679__PTR25) );
  AND2_X1 U13569 ( .A1(P3_EBX_PTR26), .A2(_02680__PTR0), .ZN(_02679__PTR26) );
  AND2_X1 U13570 ( .A1(P3_EBX_PTR27), .A2(_02680__PTR0), .ZN(_02679__PTR27) );
  AND2_X1 U13571 ( .A1(P3_EBX_PTR28), .A2(_02680__PTR0), .ZN(_02679__PTR28) );
  AND2_X1 U13572 ( .A1(P3_EBX_PTR29), .A2(_02680__PTR0), .ZN(_02679__PTR29) );
  AND2_X1 U13573 ( .A1(P3_EBX_PTR30), .A2(_02680__PTR0), .ZN(_02679__PTR30) );
  AND2_X1 U13574 ( .A1(P3_EBX_PTR31), .A2(_02680__PTR0), .ZN(_02679__PTR31) );
  AND2_X1 U13575 ( .A1(_02678__PTR32), .A2(_02680__PTR1), .ZN(_02679__PTR32) );
  AND2_X1 U13576 ( .A1(_02678__PTR33), .A2(_02680__PTR1), .ZN(_02679__PTR33) );
  AND2_X1 U13577 ( .A1(_02678__PTR34), .A2(_02680__PTR1), .ZN(_02679__PTR34) );
  AND2_X1 U13578 ( .A1(_02678__PTR35), .A2(_02680__PTR1), .ZN(_02679__PTR35) );
  AND2_X1 U13579 ( .A1(_02678__PTR36), .A2(_02680__PTR1), .ZN(_02679__PTR36) );
  AND2_X1 U13580 ( .A1(_02678__PTR37), .A2(_02680__PTR1), .ZN(_02679__PTR37) );
  AND2_X1 U13581 ( .A1(_02678__PTR38), .A2(_02680__PTR1), .ZN(_02679__PTR38) );
  AND2_X1 U13582 ( .A1(_02678__PTR39), .A2(_02680__PTR1), .ZN(_02679__PTR39) );
  AND2_X1 U13583 ( .A1(_02678__PTR40), .A2(_02680__PTR1), .ZN(_02679__PTR40) );
  AND2_X1 U13584 ( .A1(_02678__PTR41), .A2(_02680__PTR1), .ZN(_02679__PTR41) );
  AND2_X1 U13585 ( .A1(_02678__PTR42), .A2(_02680__PTR1), .ZN(_02679__PTR42) );
  AND2_X1 U13586 ( .A1(_02678__PTR43), .A2(_02680__PTR1), .ZN(_02679__PTR43) );
  AND2_X1 U13587 ( .A1(_02678__PTR44), .A2(_02680__PTR1), .ZN(_02679__PTR44) );
  AND2_X1 U13588 ( .A1(_02678__PTR45), .A2(_02680__PTR1), .ZN(_02679__PTR45) );
  AND2_X1 U13589 ( .A1(_02678__PTR46), .A2(_02680__PTR1), .ZN(_02679__PTR46) );
  AND2_X1 U13590 ( .A1(_02678__PTR47), .A2(_02680__PTR1), .ZN(_02679__PTR47) );
  AND2_X1 U13591 ( .A1(_02678__PTR48), .A2(_02680__PTR1), .ZN(_02679__PTR48) );
  AND2_X1 U13592 ( .A1(_02678__PTR49), .A2(_02680__PTR1), .ZN(_02679__PTR49) );
  AND2_X1 U13593 ( .A1(_02678__PTR50), .A2(_02680__PTR1), .ZN(_02679__PTR50) );
  AND2_X1 U13594 ( .A1(_02678__PTR51), .A2(_02680__PTR1), .ZN(_02679__PTR51) );
  AND2_X1 U13595 ( .A1(_02678__PTR52), .A2(_02680__PTR1), .ZN(_02679__PTR52) );
  AND2_X1 U13596 ( .A1(_02678__PTR53), .A2(_02680__PTR1), .ZN(_02679__PTR53) );
  AND2_X1 U13597 ( .A1(_02678__PTR54), .A2(_02680__PTR1), .ZN(_02679__PTR54) );
  AND2_X1 U13598 ( .A1(_02678__PTR55), .A2(_02680__PTR1), .ZN(_02679__PTR55) );
  AND2_X1 U13599 ( .A1(_02678__PTR56), .A2(_02680__PTR1), .ZN(_02679__PTR56) );
  AND2_X1 U13600 ( .A1(_02678__PTR57), .A2(_02680__PTR1), .ZN(_02679__PTR57) );
  AND2_X1 U13601 ( .A1(_02678__PTR58), .A2(_02680__PTR1), .ZN(_02679__PTR58) );
  AND2_X1 U13602 ( .A1(_02678__PTR59), .A2(_02680__PTR1), .ZN(_02679__PTR59) );
  AND2_X1 U13603 ( .A1(_02678__PTR60), .A2(_02680__PTR1), .ZN(_02679__PTR60) );
  AND2_X1 U13604 ( .A1(_02678__PTR61), .A2(_02680__PTR1), .ZN(_02679__PTR61) );
  AND2_X1 U13605 ( .A1(_02678__PTR62), .A2(_02680__PTR1), .ZN(_02679__PTR62) );
  AND2_X1 U13606 ( .A1(_02678__PTR63), .A2(_02680__PTR1), .ZN(_02679__PTR63) );
  AND2_X1 U13607 ( .A1(_02678__PTR64), .A2(_02680__PTR2), .ZN(_02679__PTR64) );
  AND2_X1 U13608 ( .A1(_02678__PTR65), .A2(_02680__PTR2), .ZN(_02679__PTR65) );
  AND2_X1 U13609 ( .A1(_02678__PTR66), .A2(_02680__PTR2), .ZN(_02679__PTR66) );
  AND2_X1 U13610 ( .A1(_02678__PTR67), .A2(_02680__PTR2), .ZN(_02679__PTR67) );
  AND2_X1 U13611 ( .A1(_02678__PTR68), .A2(_02680__PTR2), .ZN(_02679__PTR68) );
  AND2_X1 U13612 ( .A1(_02678__PTR69), .A2(_02680__PTR2), .ZN(_02679__PTR69) );
  AND2_X1 U13613 ( .A1(_02678__PTR70), .A2(_02680__PTR2), .ZN(_02679__PTR70) );
  AND2_X1 U13614 ( .A1(_02678__PTR71), .A2(_02680__PTR2), .ZN(_02679__PTR71) );
  AND2_X1 U13615 ( .A1(_02678__PTR72), .A2(_02680__PTR2), .ZN(_02679__PTR72) );
  AND2_X1 U13616 ( .A1(_02678__PTR73), .A2(_02680__PTR2), .ZN(_02679__PTR73) );
  AND2_X1 U13617 ( .A1(_02678__PTR74), .A2(_02680__PTR2), .ZN(_02679__PTR74) );
  AND2_X1 U13618 ( .A1(_02678__PTR75), .A2(_02680__PTR2), .ZN(_02679__PTR75) );
  AND2_X1 U13619 ( .A1(_02678__PTR76), .A2(_02680__PTR2), .ZN(_02679__PTR76) );
  AND2_X1 U13620 ( .A1(_02678__PTR77), .A2(_02680__PTR2), .ZN(_02679__PTR77) );
  AND2_X1 U13621 ( .A1(_02678__PTR78), .A2(_02680__PTR2), .ZN(_02679__PTR78) );
  AND2_X1 U13622 ( .A1(_02678__PTR79), .A2(_02680__PTR2), .ZN(_02679__PTR79) );
  AND2_X1 U13623 ( .A1(_02678__PTR80), .A2(_02680__PTR2), .ZN(_02679__PTR80) );
  AND2_X1 U13624 ( .A1(_02678__PTR81), .A2(_02680__PTR2), .ZN(_02679__PTR81) );
  AND2_X1 U13625 ( .A1(_02678__PTR82), .A2(_02680__PTR2), .ZN(_02679__PTR82) );
  AND2_X1 U13626 ( .A1(_02678__PTR83), .A2(_02680__PTR2), .ZN(_02679__PTR83) );
  AND2_X1 U13627 ( .A1(_02678__PTR84), .A2(_02680__PTR2), .ZN(_02679__PTR84) );
  AND2_X1 U13628 ( .A1(_02678__PTR85), .A2(_02680__PTR2), .ZN(_02679__PTR85) );
  AND2_X1 U13629 ( .A1(_02678__PTR86), .A2(_02680__PTR2), .ZN(_02679__PTR86) );
  AND2_X1 U13630 ( .A1(_02678__PTR87), .A2(_02680__PTR2), .ZN(_02679__PTR87) );
  AND2_X1 U13631 ( .A1(_02678__PTR88), .A2(_02680__PTR2), .ZN(_02679__PTR88) );
  AND2_X1 U13632 ( .A1(_02678__PTR89), .A2(_02680__PTR2), .ZN(_02679__PTR89) );
  AND2_X1 U13633 ( .A1(_02678__PTR90), .A2(_02680__PTR2), .ZN(_02679__PTR90) );
  AND2_X1 U13634 ( .A1(_02678__PTR91), .A2(_02680__PTR2), .ZN(_02679__PTR91) );
  AND2_X1 U13635 ( .A1(_02678__PTR92), .A2(_02680__PTR2), .ZN(_02679__PTR92) );
  AND2_X1 U13636 ( .A1(_02678__PTR93), .A2(_02680__PTR2), .ZN(_02679__PTR93) );
  AND2_X1 U13637 ( .A1(_02678__PTR94), .A2(_02680__PTR2), .ZN(_02679__PTR94) );
  AND2_X1 U13638 ( .A1(_02678__PTR95), .A2(_02680__PTR2), .ZN(_02679__PTR95) );
  AND2_X1 U13639 ( .A1(P3_EAX_PTR0), .A2(_02676__PTR0), .ZN(_02675__PTR0) );
  AND2_X1 U13640 ( .A1(P3_EAX_PTR1), .A2(_02676__PTR0), .ZN(_02675__PTR1) );
  AND2_X1 U13641 ( .A1(P3_EAX_PTR2), .A2(_02676__PTR0), .ZN(_02675__PTR2) );
  AND2_X1 U13642 ( .A1(P3_EAX_PTR3), .A2(_02676__PTR0), .ZN(_02675__PTR3) );
  AND2_X1 U13643 ( .A1(P3_EAX_PTR4), .A2(_02676__PTR0), .ZN(_02675__PTR4) );
  AND2_X1 U13644 ( .A1(P3_EAX_PTR5), .A2(_02676__PTR0), .ZN(_02675__PTR5) );
  AND2_X1 U13645 ( .A1(P3_EAX_PTR6), .A2(_02676__PTR0), .ZN(_02675__PTR6) );
  AND2_X1 U13646 ( .A1(P3_EAX_PTR7), .A2(_02676__PTR0), .ZN(_02675__PTR7) );
  AND2_X1 U13647 ( .A1(P3_EAX_PTR8), .A2(_02676__PTR0), .ZN(_02675__PTR8) );
  AND2_X1 U13648 ( .A1(P3_EAX_PTR9), .A2(_02676__PTR0), .ZN(_02675__PTR9) );
  AND2_X1 U13649 ( .A1(P3_EAX_PTR10), .A2(_02676__PTR0), .ZN(_02675__PTR10) );
  AND2_X1 U13650 ( .A1(P3_EAX_PTR11), .A2(_02676__PTR0), .ZN(_02675__PTR11) );
  AND2_X1 U13651 ( .A1(P3_EAX_PTR12), .A2(_02676__PTR0), .ZN(_02675__PTR12) );
  AND2_X1 U13652 ( .A1(P3_EAX_PTR13), .A2(_02676__PTR0), .ZN(_02675__PTR13) );
  AND2_X1 U13653 ( .A1(P3_EAX_PTR14), .A2(_02676__PTR0), .ZN(_02675__PTR14) );
  AND2_X1 U13654 ( .A1(P3_EAX_PTR15), .A2(_02676__PTR0), .ZN(_02675__PTR15) );
  AND2_X1 U13655 ( .A1(P3_EAX_PTR16), .A2(_02676__PTR0), .ZN(_02675__PTR16) );
  AND2_X1 U13656 ( .A1(P3_EAX_PTR17), .A2(_02676__PTR0), .ZN(_02675__PTR17) );
  AND2_X1 U13657 ( .A1(P3_EAX_PTR18), .A2(_02676__PTR0), .ZN(_02675__PTR18) );
  AND2_X1 U13658 ( .A1(P3_EAX_PTR19), .A2(_02676__PTR0), .ZN(_02675__PTR19) );
  AND2_X1 U13659 ( .A1(P3_EAX_PTR20), .A2(_02676__PTR0), .ZN(_02675__PTR20) );
  AND2_X1 U13660 ( .A1(P3_EAX_PTR21), .A2(_02676__PTR0), .ZN(_02675__PTR21) );
  AND2_X1 U13661 ( .A1(P3_EAX_PTR22), .A2(_02676__PTR0), .ZN(_02675__PTR22) );
  AND2_X1 U13662 ( .A1(P3_EAX_PTR23), .A2(_02676__PTR0), .ZN(_02675__PTR23) );
  AND2_X1 U13663 ( .A1(P3_EAX_PTR24), .A2(_02676__PTR0), .ZN(_02675__PTR24) );
  AND2_X1 U13664 ( .A1(P3_EAX_PTR25), .A2(_02676__PTR0), .ZN(_02675__PTR25) );
  AND2_X1 U13665 ( .A1(P3_EAX_PTR26), .A2(_02676__PTR0), .ZN(_02675__PTR26) );
  AND2_X1 U13666 ( .A1(P3_EAX_PTR27), .A2(_02676__PTR0), .ZN(_02675__PTR27) );
  AND2_X1 U13667 ( .A1(P3_EAX_PTR28), .A2(_02676__PTR0), .ZN(_02675__PTR28) );
  AND2_X1 U13668 ( .A1(P3_EAX_PTR29), .A2(_02676__PTR0), .ZN(_02675__PTR29) );
  AND2_X1 U13669 ( .A1(P3_EAX_PTR30), .A2(_02676__PTR0), .ZN(_02675__PTR30) );
  AND2_X1 U13670 ( .A1(P3_EAX_PTR31), .A2(_02676__PTR0), .ZN(_02675__PTR31) );
  AND2_X1 U13671 ( .A1(_02674__PTR32), .A2(_02676__PTR1), .ZN(_02675__PTR32) );
  AND2_X1 U13672 ( .A1(_02674__PTR33), .A2(_02676__PTR1), .ZN(_02675__PTR33) );
  AND2_X1 U13673 ( .A1(_02674__PTR34), .A2(_02676__PTR1), .ZN(_02675__PTR34) );
  AND2_X1 U13674 ( .A1(_02674__PTR35), .A2(_02676__PTR1), .ZN(_02675__PTR35) );
  AND2_X1 U13675 ( .A1(_02674__PTR36), .A2(_02676__PTR1), .ZN(_02675__PTR36) );
  AND2_X1 U13676 ( .A1(_02674__PTR37), .A2(_02676__PTR1), .ZN(_02675__PTR37) );
  AND2_X1 U13677 ( .A1(_02674__PTR38), .A2(_02676__PTR1), .ZN(_02675__PTR38) );
  AND2_X1 U13678 ( .A1(_02674__PTR39), .A2(_02676__PTR1), .ZN(_02675__PTR39) );
  AND2_X1 U13679 ( .A1(_02674__PTR40), .A2(_02676__PTR1), .ZN(_02675__PTR40) );
  AND2_X1 U13680 ( .A1(_02674__PTR41), .A2(_02676__PTR1), .ZN(_02675__PTR41) );
  AND2_X1 U13681 ( .A1(_02674__PTR42), .A2(_02676__PTR1), .ZN(_02675__PTR42) );
  AND2_X1 U13682 ( .A1(_02674__PTR43), .A2(_02676__PTR1), .ZN(_02675__PTR43) );
  AND2_X1 U13683 ( .A1(_02674__PTR44), .A2(_02676__PTR1), .ZN(_02675__PTR44) );
  AND2_X1 U13684 ( .A1(_02674__PTR45), .A2(_02676__PTR1), .ZN(_02675__PTR45) );
  AND2_X1 U13685 ( .A1(_02674__PTR46), .A2(_02676__PTR1), .ZN(_02675__PTR46) );
  AND2_X1 U13686 ( .A1(_02674__PTR47), .A2(_02676__PTR1), .ZN(_02675__PTR47) );
  AND2_X1 U13687 ( .A1(_02674__PTR48), .A2(_02676__PTR1), .ZN(_02675__PTR48) );
  AND2_X1 U13688 ( .A1(_02674__PTR49), .A2(_02676__PTR1), .ZN(_02675__PTR49) );
  AND2_X1 U13689 ( .A1(_02674__PTR50), .A2(_02676__PTR1), .ZN(_02675__PTR50) );
  AND2_X1 U13690 ( .A1(_02674__PTR51), .A2(_02676__PTR1), .ZN(_02675__PTR51) );
  AND2_X1 U13691 ( .A1(_02674__PTR52), .A2(_02676__PTR1), .ZN(_02675__PTR52) );
  AND2_X1 U13692 ( .A1(_02674__PTR53), .A2(_02676__PTR1), .ZN(_02675__PTR53) );
  AND2_X1 U13693 ( .A1(_02674__PTR54), .A2(_02676__PTR1), .ZN(_02675__PTR54) );
  AND2_X1 U13694 ( .A1(_02674__PTR55), .A2(_02676__PTR1), .ZN(_02675__PTR55) );
  AND2_X1 U13695 ( .A1(_02674__PTR56), .A2(_02676__PTR1), .ZN(_02675__PTR56) );
  AND2_X1 U13696 ( .A1(_02674__PTR57), .A2(_02676__PTR1), .ZN(_02675__PTR57) );
  AND2_X1 U13697 ( .A1(_02674__PTR58), .A2(_02676__PTR1), .ZN(_02675__PTR58) );
  AND2_X1 U13698 ( .A1(_02674__PTR59), .A2(_02676__PTR1), .ZN(_02675__PTR59) );
  AND2_X1 U13699 ( .A1(_02674__PTR60), .A2(_02676__PTR1), .ZN(_02675__PTR60) );
  AND2_X1 U13700 ( .A1(_02674__PTR61), .A2(_02676__PTR1), .ZN(_02675__PTR61) );
  AND2_X1 U13701 ( .A1(_02674__PTR62), .A2(_02676__PTR1), .ZN(_02675__PTR62) );
  AND2_X1 U13702 ( .A1(_02674__PTR63), .A2(_02676__PTR1), .ZN(_02675__PTR63) );
  AND2_X1 U13703 ( .A1(_02674__PTR96), .A2(_02668__PTR3), .ZN(_02675__PTR64) );
  AND2_X1 U13704 ( .A1(_02674__PTR97), .A2(_02668__PTR3), .ZN(_02675__PTR65) );
  AND2_X1 U13705 ( .A1(_02674__PTR98), .A2(_02668__PTR3), .ZN(_02675__PTR66) );
  AND2_X1 U13706 ( .A1(_02674__PTR99), .A2(_02668__PTR3), .ZN(_02675__PTR67) );
  AND2_X1 U13707 ( .A1(_02674__PTR100), .A2(_02668__PTR3), .ZN(_02675__PTR68) );
  AND2_X1 U13708 ( .A1(_02674__PTR101), .A2(_02668__PTR3), .ZN(_02675__PTR69) );
  AND2_X1 U13709 ( .A1(_02674__PTR102), .A2(_02668__PTR3), .ZN(_02675__PTR70) );
  AND2_X1 U13710 ( .A1(_02674__PTR103), .A2(_02668__PTR3), .ZN(_02675__PTR71) );
  AND2_X1 U13711 ( .A1(_02674__PTR104), .A2(_02668__PTR3), .ZN(_02675__PTR72) );
  AND2_X1 U13712 ( .A1(_02674__PTR105), .A2(_02668__PTR3), .ZN(_02675__PTR73) );
  AND2_X1 U13713 ( .A1(_02674__PTR106), .A2(_02668__PTR3), .ZN(_02675__PTR74) );
  AND2_X1 U13714 ( .A1(_02674__PTR107), .A2(_02668__PTR3), .ZN(_02675__PTR75) );
  AND2_X1 U13715 ( .A1(_02674__PTR108), .A2(_02668__PTR3), .ZN(_02675__PTR76) );
  AND2_X1 U13716 ( .A1(_02674__PTR109), .A2(_02668__PTR3), .ZN(_02675__PTR77) );
  AND2_X1 U13717 ( .A1(_02674__PTR110), .A2(_02668__PTR3), .ZN(_02675__PTR78) );
  AND2_X1 U13718 ( .A1(_02674__PTR111), .A2(_02668__PTR3), .ZN(_02675__PTR79) );
  AND2_X1 U13719 ( .A1(_02674__PTR80), .A2(_02668__PTR3), .ZN(_02675__PTR80) );
  AND2_X1 U13720 ( .A1(_02674__PTR81), .A2(_02668__PTR3), .ZN(_02675__PTR81) );
  AND2_X1 U13721 ( .A1(_02674__PTR82), .A2(_02668__PTR3), .ZN(_02675__PTR82) );
  AND2_X1 U13722 ( .A1(_02674__PTR83), .A2(_02668__PTR3), .ZN(_02675__PTR83) );
  AND2_X1 U13723 ( .A1(_02674__PTR84), .A2(_02668__PTR3), .ZN(_02675__PTR84) );
  AND2_X1 U13724 ( .A1(_02674__PTR85), .A2(_02668__PTR3), .ZN(_02675__PTR85) );
  AND2_X1 U13725 ( .A1(_02674__PTR86), .A2(_02668__PTR3), .ZN(_02675__PTR86) );
  AND2_X1 U13726 ( .A1(_02674__PTR87), .A2(_02668__PTR3), .ZN(_02675__PTR87) );
  AND2_X1 U13727 ( .A1(_02674__PTR88), .A2(_02668__PTR3), .ZN(_02675__PTR88) );
  AND2_X1 U13728 ( .A1(_02674__PTR89), .A2(_02668__PTR3), .ZN(_02675__PTR89) );
  AND2_X1 U13729 ( .A1(_02674__PTR90), .A2(_02668__PTR3), .ZN(_02675__PTR90) );
  AND2_X1 U13730 ( .A1(_02674__PTR91), .A2(_02668__PTR3), .ZN(_02675__PTR91) );
  AND2_X1 U13731 ( .A1(_02674__PTR92), .A2(_02668__PTR3), .ZN(_02675__PTR92) );
  AND2_X1 U13732 ( .A1(_02674__PTR93), .A2(_02668__PTR3), .ZN(_02675__PTR93) );
  AND2_X1 U13733 ( .A1(_02674__PTR94), .A2(_02668__PTR3), .ZN(_02675__PTR94) );
  AND2_X1 U13734 ( .A1(_02674__PTR95), .A2(_02668__PTR3), .ZN(_02675__PTR95) );
  AND2_X1 U13735 ( .A1(_02674__PTR96), .A2(_02668__PTR4), .ZN(_02675__PTR96) );
  AND2_X1 U13736 ( .A1(_02674__PTR97), .A2(_02668__PTR4), .ZN(_02675__PTR97) );
  AND2_X1 U13737 ( .A1(_02674__PTR98), .A2(_02668__PTR4), .ZN(_02675__PTR98) );
  AND2_X1 U13738 ( .A1(_02674__PTR99), .A2(_02668__PTR4), .ZN(_02675__PTR99) );
  AND2_X1 U13739 ( .A1(_02674__PTR100), .A2(_02668__PTR4), .ZN(_02675__PTR100) );
  AND2_X1 U13740 ( .A1(_02674__PTR101), .A2(_02668__PTR4), .ZN(_02675__PTR101) );
  AND2_X1 U13741 ( .A1(_02674__PTR102), .A2(_02668__PTR4), .ZN(_02675__PTR102) );
  AND2_X1 U13742 ( .A1(_02674__PTR103), .A2(_02668__PTR4), .ZN(_02675__PTR103) );
  AND2_X1 U13743 ( .A1(_02674__PTR104), .A2(_02668__PTR4), .ZN(_02675__PTR104) );
  AND2_X1 U13744 ( .A1(_02674__PTR105), .A2(_02668__PTR4), .ZN(_02675__PTR105) );
  AND2_X1 U13745 ( .A1(_02674__PTR106), .A2(_02668__PTR4), .ZN(_02675__PTR106) );
  AND2_X1 U13746 ( .A1(_02674__PTR107), .A2(_02668__PTR4), .ZN(_02675__PTR107) );
  AND2_X1 U13747 ( .A1(_02674__PTR108), .A2(_02668__PTR4), .ZN(_02675__PTR108) );
  AND2_X1 U13748 ( .A1(_02674__PTR109), .A2(_02668__PTR4), .ZN(_02675__PTR109) );
  AND2_X1 U13749 ( .A1(_02674__PTR110), .A2(_02668__PTR4), .ZN(_02675__PTR110) );
  AND2_X1 U13750 ( .A1(_02674__PTR111), .A2(_02668__PTR4), .ZN(_02675__PTR111) );
  AND2_X1 U13751 ( .A1(_02674__PTR112), .A2(_02668__PTR4), .ZN(_02675__PTR112) );
  AND2_X1 U13752 ( .A1(_02674__PTR113), .A2(_02668__PTR4), .ZN(_02675__PTR113) );
  AND2_X1 U13753 ( .A1(_02674__PTR114), .A2(_02668__PTR4), .ZN(_02675__PTR114) );
  AND2_X1 U13754 ( .A1(_02674__PTR115), .A2(_02668__PTR4), .ZN(_02675__PTR115) );
  AND2_X1 U13755 ( .A1(_02674__PTR116), .A2(_02668__PTR4), .ZN(_02675__PTR116) );
  AND2_X1 U13756 ( .A1(_02674__PTR117), .A2(_02668__PTR4), .ZN(_02675__PTR117) );
  AND2_X1 U13757 ( .A1(_02674__PTR118), .A2(_02668__PTR4), .ZN(_02675__PTR118) );
  AND2_X1 U13758 ( .A1(_02674__PTR119), .A2(_02668__PTR4), .ZN(_02675__PTR119) );
  AND2_X1 U13759 ( .A1(_02674__PTR120), .A2(_02668__PTR4), .ZN(_02675__PTR120) );
  AND2_X1 U13760 ( .A1(_02674__PTR121), .A2(_02668__PTR4), .ZN(_02675__PTR121) );
  AND2_X1 U13761 ( .A1(_02674__PTR122), .A2(_02668__PTR4), .ZN(_02675__PTR122) );
  AND2_X1 U13762 ( .A1(_02674__PTR123), .A2(_02668__PTR4), .ZN(_02675__PTR123) );
  AND2_X1 U13763 ( .A1(_02674__PTR124), .A2(_02668__PTR4), .ZN(_02675__PTR124) );
  AND2_X1 U13764 ( .A1(_02674__PTR125), .A2(_02668__PTR4), .ZN(_02675__PTR125) );
  AND2_X1 U13765 ( .A1(_02674__PTR126), .A2(_02668__PTR4), .ZN(_02675__PTR126) );
  AND2_X1 U13766 ( .A1(_02674__PTR127), .A2(_02668__PTR4), .ZN(_02675__PTR127) );
  AND2_X1 U13767 ( .A1(_02674__PTR128), .A2(_02676__PTR4), .ZN(_02675__PTR128) );
  AND2_X1 U13768 ( .A1(_02674__PTR129), .A2(_02676__PTR4), .ZN(_02675__PTR129) );
  AND2_X1 U13769 ( .A1(_02674__PTR130), .A2(_02676__PTR4), .ZN(_02675__PTR130) );
  AND2_X1 U13770 ( .A1(_02674__PTR131), .A2(_02676__PTR4), .ZN(_02675__PTR131) );
  AND2_X1 U13771 ( .A1(_02674__PTR132), .A2(_02676__PTR4), .ZN(_02675__PTR132) );
  AND2_X1 U13772 ( .A1(_02674__PTR133), .A2(_02676__PTR4), .ZN(_02675__PTR133) );
  AND2_X1 U13773 ( .A1(_02674__PTR134), .A2(_02676__PTR4), .ZN(_02675__PTR134) );
  AND2_X1 U13774 ( .A1(_02674__PTR135), .A2(_02676__PTR4), .ZN(_02675__PTR135) );
  AND2_X1 U13775 ( .A1(_02674__PTR136), .A2(_02676__PTR4), .ZN(_02675__PTR136) );
  AND2_X1 U13776 ( .A1(_02674__PTR137), .A2(_02676__PTR4), .ZN(_02675__PTR137) );
  AND2_X1 U13777 ( .A1(_02674__PTR138), .A2(_02676__PTR4), .ZN(_02675__PTR138) );
  AND2_X1 U13778 ( .A1(_02674__PTR139), .A2(_02676__PTR4), .ZN(_02675__PTR139) );
  AND2_X1 U13779 ( .A1(_02674__PTR140), .A2(_02676__PTR4), .ZN(_02675__PTR140) );
  AND2_X1 U13780 ( .A1(_02674__PTR141), .A2(_02676__PTR4), .ZN(_02675__PTR141) );
  AND2_X1 U13781 ( .A1(_02674__PTR142), .A2(_02676__PTR4), .ZN(_02675__PTR142) );
  AND2_X1 U13782 ( .A1(_02674__PTR143), .A2(_02676__PTR4), .ZN(_02675__PTR143) );
  AND2_X1 U13783 ( .A1(_02674__PTR144), .A2(_02676__PTR4), .ZN(_02675__PTR144) );
  AND2_X1 U13784 ( .A1(_02674__PTR145), .A2(_02676__PTR4), .ZN(_02675__PTR145) );
  AND2_X1 U13785 ( .A1(_02674__PTR146), .A2(_02676__PTR4), .ZN(_02675__PTR146) );
  AND2_X1 U13786 ( .A1(_02674__PTR147), .A2(_02676__PTR4), .ZN(_02675__PTR147) );
  AND2_X1 U13787 ( .A1(_02674__PTR148), .A2(_02676__PTR4), .ZN(_02675__PTR148) );
  AND2_X1 U13788 ( .A1(_02674__PTR149), .A2(_02676__PTR4), .ZN(_02675__PTR149) );
  AND2_X1 U13789 ( .A1(_02674__PTR150), .A2(_02676__PTR4), .ZN(_02675__PTR150) );
  AND2_X1 U13790 ( .A1(_02674__PTR151), .A2(_02676__PTR4), .ZN(_02675__PTR151) );
  AND2_X1 U13791 ( .A1(_02674__PTR152), .A2(_02676__PTR4), .ZN(_02675__PTR152) );
  AND2_X1 U13792 ( .A1(_02674__PTR153), .A2(_02676__PTR4), .ZN(_02675__PTR153) );
  AND2_X1 U13793 ( .A1(_02674__PTR154), .A2(_02676__PTR4), .ZN(_02675__PTR154) );
  AND2_X1 U13794 ( .A1(_02674__PTR155), .A2(_02676__PTR4), .ZN(_02675__PTR155) );
  AND2_X1 U13795 ( .A1(_02674__PTR156), .A2(_02676__PTR4), .ZN(_02675__PTR156) );
  AND2_X1 U13796 ( .A1(_02674__PTR157), .A2(_02676__PTR4), .ZN(_02675__PTR157) );
  AND2_X1 U13797 ( .A1(_02674__PTR158), .A2(_02676__PTR4), .ZN(_02675__PTR158) );
  AND2_X1 U13798 ( .A1(_02674__PTR159), .A2(_02676__PTR4), .ZN(_02675__PTR159) );
  AND2_X1 U13799 ( .A1(_02439__PTR0), .A2(_02437__PTR0), .ZN(_02440__PTR0) );
  AND2_X1 U13800 ( .A1(_02439__PTR1), .A2(_02437__PTR1), .ZN(_02440__PTR1) );
  AND2_X1 U13801 ( .A1(_02439__PTR2), .A2(_02441__PTR2), .ZN(_02440__PTR2) );
  AND2_X1 U13802 ( .A1(_02439__PTR3), .A2(_02437__PTR3), .ZN(_02440__PTR3) );
  AND2_X1 U13803 ( .A1(_02435__PTR0), .A2(_02437__PTR0), .ZN(_02436__PTR0) );
  AND2_X1 U13804 ( .A1(_02435__PTR1), .A2(_02437__PTR1), .ZN(_02436__PTR1) );
  AND2_X1 U13805 ( .A1(_02435__PTR2), .A2(_02437__PTR2), .ZN(_02436__PTR2) );
  AND2_X1 U13806 ( .A1(_02435__PTR3), .A2(_02437__PTR3), .ZN(_02436__PTR3) );
  AND2_X1 U13807 ( .A1(_02465__PTR3), .A2(_02664__PTR0), .ZN(_02667__PTR0) );
  AND2_X1 U13808 ( .A1(_02465__PTR4), .A2(_02664__PTR0), .ZN(_02667__PTR1) );
  AND2_X1 U13809 ( .A1(_02465__PTR5), .A2(_02664__PTR0), .ZN(_02667__PTR2) );
  AND2_X1 U13810 ( .A1(_02465__PTR6), .A2(_02664__PTR0), .ZN(_02667__PTR3) );
  AND2_X1 U13811 ( .A1(P3_P1_InstQueueRd_Addr_PTR0), .A2(_02664__PTR1), .ZN(_02667__PTR5) );
  AND2_X1 U13812 ( .A1(_02471__PTR4), .A2(_02664__PTR1), .ZN(_02667__PTR6) );
  AND2_X1 U13813 ( .A1(_02471__PTR5), .A2(_02664__PTR1), .ZN(_02667__PTR7) );
  AND2_X1 U13814 ( .A1(_02471__PTR6), .A2(_02664__PTR1), .ZN(_02667__PTR8) );
  AND2_X1 U13815 ( .A1(P3_P1_InstQueueRd_Addr_PTR0), .A2(_02437__PTR0), .ZN(_02667__PTR10) );
  AND2_X1 U13816 ( .A1(_02666__PTR11), .A2(_02437__PTR0), .ZN(_02667__PTR11) );
  AND2_X1 U13817 ( .A1(_02666__PTR12), .A2(_02437__PTR0), .ZN(_02667__PTR12) );
  AND2_X1 U13818 ( .A1(_02666__PTR13), .A2(_02437__PTR0), .ZN(_02667__PTR13) );
  AND2_X1 U13819 ( .A1(_02666__PTR14), .A2(_02437__PTR0), .ZN(_02667__PTR14) );
  AND2_X1 U13820 ( .A1(P3_P1_InstQueueRd_Addr_PTR0), .A2(_02668__PTR3), .ZN(_02667__PTR15) );
  AND2_X1 U13821 ( .A1(_02666__PTR21), .A2(_02668__PTR3), .ZN(_02667__PTR16) );
  AND2_X1 U13822 ( .A1(_02666__PTR22), .A2(_02668__PTR3), .ZN(_02667__PTR17) );
  AND2_X1 U13823 ( .A1(_02666__PTR23), .A2(_02668__PTR3), .ZN(_02667__PTR18) );
  AND2_X1 U13824 ( .A1(_02666__PTR19), .A2(_02668__PTR3), .ZN(_02667__PTR19) );
  AND2_X1 U13825 ( .A1(P3_P1_InstQueueRd_Addr_PTR0), .A2(_02668__PTR4), .ZN(_02667__PTR20) );
  AND2_X1 U13826 ( .A1(_02666__PTR21), .A2(_02668__PTR4), .ZN(_02667__PTR21) );
  AND2_X1 U13827 ( .A1(_02666__PTR22), .A2(_02668__PTR4), .ZN(_02667__PTR22) );
  AND2_X1 U13828 ( .A1(_02666__PTR23), .A2(_02668__PTR4), .ZN(_02667__PTR23) );
  AND2_X1 U13829 ( .A1(_02666__PTR24), .A2(_02668__PTR4), .ZN(_02667__PTR24) );
  AND2_X1 U13830 ( .A1(_02666__PTR25), .A2(_02664__PTR4), .ZN(_02667__PTR25) );
  AND2_X1 U13831 ( .A1(_02666__PTR26), .A2(_02664__PTR4), .ZN(_02667__PTR26) );
  AND2_X1 U13832 ( .A1(_02666__PTR27), .A2(_02664__PTR4), .ZN(_02667__PTR27) );
  AND2_X1 U13833 ( .A1(_02666__PTR28), .A2(_02664__PTR4), .ZN(_02667__PTR28) );
  AND2_X1 U13834 ( .A1(_02666__PTR29), .A2(_02664__PTR4), .ZN(_02667__PTR29) );
  AND2_X1 U13835 ( .A1(P3_P1_InstQueueRd_Addr_PTR0), .A2(_02668__PTR6), .ZN(_02667__PTR30) );
  AND2_X1 U13836 ( .A1(P3_P1_InstQueueRd_Addr_PTR1), .A2(_02668__PTR6), .ZN(_02667__PTR31) );
  AND2_X1 U13837 ( .A1(P3_P1_InstQueueRd_Addr_PTR2), .A2(_02668__PTR6), .ZN(_02667__PTR32) );
  AND2_X1 U13838 ( .A1(P3_P1_InstQueueRd_Addr_PTR3), .A2(_02668__PTR6), .ZN(_02667__PTR33) );
  AND2_X1 U13839 ( .A1(P3_P1_InstQueueRd_Addr_PTR4), .A2(_02668__PTR6), .ZN(_02667__PTR34) );
  AND2_X1 U13840 ( .A1(_02454__PTR0), .A2(_02456__PTR0), .ZN(_02455__PTR0) );
  AND2_X1 U13841 ( .A1(P3_CodeFetch), .A2(_02445__PTR3), .ZN(_02455__PTR1) );
  AND2_X1 U13842 ( .A1(_02443__PTR0), .A2(_02445__PTR0), .ZN(_02444__PTR0) );
  AND2_X1 U13843 ( .A1(_02443__PTR1), .A2(_02437__PTR1), .ZN(_02444__PTR1) );
  AND2_X1 U13844 ( .A1(_02443__PTR2), .A2(_02445__PTR2), .ZN(_02444__PTR2) );
  AND2_X1 U13845 ( .A1(P3_RequestPending), .A2(_02445__PTR3), .ZN(_02444__PTR3) );
  AND2_X1 U13846 ( .A1(_02450__PTR0), .A2(_02452__PTR0), .ZN(_02451__PTR0) );
  AND2_X1 U13847 ( .A1(_02450__PTR1), .A2(_02452__PTR1), .ZN(_02451__PTR1) );
  AND2_X1 U13848 ( .A1(P3_MemoryFetch), .A2(_02445__PTR3), .ZN(_02451__PTR2) );
  AND2_X1 U13849 ( .A1(_02447__PTR0), .A2(_02437__PTR0), .ZN(_02448__PTR0) );
  AND2_X1 U13850 ( .A1(_02447__PTR1), .A2(_02437__PTR1), .ZN(_02448__PTR1) );
  AND2_X1 U13851 ( .A1(P3_ReadRequest), .A2(_02445__PTR3), .ZN(_02448__PTR2) );
  AND2_X1 U13852 ( .A1(P3_rEIP_PTR0), .A2(_02445__PTR3), .ZN(_02683__PTR0) );
  AND2_X1 U13853 ( .A1(P3_rEIP_PTR1), .A2(_02445__PTR3), .ZN(_02683__PTR1) );
  AND2_X1 U13854 ( .A1(P3_rEIP_PTR2), .A2(_02445__PTR3), .ZN(_02683__PTR2) );
  AND2_X1 U13855 ( .A1(P3_rEIP_PTR3), .A2(_02445__PTR3), .ZN(_02683__PTR3) );
  AND2_X1 U13856 ( .A1(P3_rEIP_PTR4), .A2(_02445__PTR3), .ZN(_02683__PTR4) );
  AND2_X1 U13857 ( .A1(P3_rEIP_PTR5), .A2(_02445__PTR3), .ZN(_02683__PTR5) );
  AND2_X1 U13858 ( .A1(P3_rEIP_PTR6), .A2(_02445__PTR3), .ZN(_02683__PTR6) );
  AND2_X1 U13859 ( .A1(P3_rEIP_PTR7), .A2(_02445__PTR3), .ZN(_02683__PTR7) );
  AND2_X1 U13860 ( .A1(P3_rEIP_PTR8), .A2(_02445__PTR3), .ZN(_02683__PTR8) );
  AND2_X1 U13861 ( .A1(P3_rEIP_PTR9), .A2(_02445__PTR3), .ZN(_02683__PTR9) );
  AND2_X1 U13862 ( .A1(P3_rEIP_PTR10), .A2(_02445__PTR3), .ZN(_02683__PTR10) );
  AND2_X1 U13863 ( .A1(P3_rEIP_PTR11), .A2(_02445__PTR3), .ZN(_02683__PTR11) );
  AND2_X1 U13864 ( .A1(P3_rEIP_PTR12), .A2(_02445__PTR3), .ZN(_02683__PTR12) );
  AND2_X1 U13865 ( .A1(P3_rEIP_PTR13), .A2(_02445__PTR3), .ZN(_02683__PTR13) );
  AND2_X1 U13866 ( .A1(P3_rEIP_PTR14), .A2(_02445__PTR3), .ZN(_02683__PTR14) );
  AND2_X1 U13867 ( .A1(P3_rEIP_PTR15), .A2(_02445__PTR3), .ZN(_02683__PTR15) );
  AND2_X1 U13868 ( .A1(P3_rEIP_PTR16), .A2(_02445__PTR3), .ZN(_02683__PTR16) );
  AND2_X1 U13869 ( .A1(P3_rEIP_PTR17), .A2(_02445__PTR3), .ZN(_02683__PTR17) );
  AND2_X1 U13870 ( .A1(P3_rEIP_PTR18), .A2(_02445__PTR3), .ZN(_02683__PTR18) );
  AND2_X1 U13871 ( .A1(P3_rEIP_PTR19), .A2(_02445__PTR3), .ZN(_02683__PTR19) );
  AND2_X1 U13872 ( .A1(P3_rEIP_PTR20), .A2(_02445__PTR3), .ZN(_02683__PTR20) );
  AND2_X1 U13873 ( .A1(P3_rEIP_PTR21), .A2(_02445__PTR3), .ZN(_02683__PTR21) );
  AND2_X1 U13874 ( .A1(P3_rEIP_PTR22), .A2(_02445__PTR3), .ZN(_02683__PTR22) );
  AND2_X1 U13875 ( .A1(P3_rEIP_PTR23), .A2(_02445__PTR3), .ZN(_02683__PTR23) );
  AND2_X1 U13876 ( .A1(P3_rEIP_PTR24), .A2(_02445__PTR3), .ZN(_02683__PTR24) );
  AND2_X1 U13877 ( .A1(P3_rEIP_PTR25), .A2(_02445__PTR3), .ZN(_02683__PTR25) );
  AND2_X1 U13878 ( .A1(P3_rEIP_PTR26), .A2(_02445__PTR3), .ZN(_02683__PTR26) );
  AND2_X1 U13879 ( .A1(P3_rEIP_PTR27), .A2(_02445__PTR3), .ZN(_02683__PTR27) );
  AND2_X1 U13880 ( .A1(P3_rEIP_PTR28), .A2(_02445__PTR3), .ZN(_02683__PTR28) );
  AND2_X1 U13881 ( .A1(P3_rEIP_PTR29), .A2(_02445__PTR3), .ZN(_02683__PTR29) );
  AND2_X1 U13882 ( .A1(P3_rEIP_PTR30), .A2(_02445__PTR3), .ZN(_02683__PTR30) );
  AND2_X1 U13883 ( .A1(P3_rEIP_PTR31), .A2(_02445__PTR3), .ZN(_02683__PTR31) );
  AND2_X1 U13884 ( .A1(_02682__PTR32), .A2(_02452__PTR0), .ZN(_02683__PTR32) );
  AND2_X1 U13885 ( .A1(_02682__PTR33), .A2(_02452__PTR0), .ZN(_02683__PTR33) );
  AND2_X1 U13886 ( .A1(_02682__PTR34), .A2(_02452__PTR0), .ZN(_02683__PTR34) );
  AND2_X1 U13887 ( .A1(_02682__PTR35), .A2(_02452__PTR0), .ZN(_02683__PTR35) );
  AND2_X1 U13888 ( .A1(_02682__PTR36), .A2(_02452__PTR0), .ZN(_02683__PTR36) );
  AND2_X1 U13889 ( .A1(_02682__PTR37), .A2(_02452__PTR0), .ZN(_02683__PTR37) );
  AND2_X1 U13890 ( .A1(_02682__PTR38), .A2(_02452__PTR0), .ZN(_02683__PTR38) );
  AND2_X1 U13891 ( .A1(_02682__PTR39), .A2(_02452__PTR0), .ZN(_02683__PTR39) );
  AND2_X1 U13892 ( .A1(_02682__PTR40), .A2(_02452__PTR0), .ZN(_02683__PTR40) );
  AND2_X1 U13893 ( .A1(_02682__PTR41), .A2(_02452__PTR0), .ZN(_02683__PTR41) );
  AND2_X1 U13894 ( .A1(_02682__PTR42), .A2(_02452__PTR0), .ZN(_02683__PTR42) );
  AND2_X1 U13895 ( .A1(_02682__PTR43), .A2(_02452__PTR0), .ZN(_02683__PTR43) );
  AND2_X1 U13896 ( .A1(_02682__PTR44), .A2(_02452__PTR0), .ZN(_02683__PTR44) );
  AND2_X1 U13897 ( .A1(_02682__PTR45), .A2(_02452__PTR0), .ZN(_02683__PTR45) );
  AND2_X1 U13898 ( .A1(_02682__PTR46), .A2(_02452__PTR0), .ZN(_02683__PTR46) );
  AND2_X1 U13899 ( .A1(_02682__PTR47), .A2(_02452__PTR0), .ZN(_02683__PTR47) );
  AND2_X1 U13900 ( .A1(_02682__PTR48), .A2(_02452__PTR0), .ZN(_02683__PTR48) );
  AND2_X1 U13901 ( .A1(_02682__PTR49), .A2(_02452__PTR0), .ZN(_02683__PTR49) );
  AND2_X1 U13902 ( .A1(_02682__PTR50), .A2(_02452__PTR0), .ZN(_02683__PTR50) );
  AND2_X1 U13903 ( .A1(_02682__PTR51), .A2(_02452__PTR0), .ZN(_02683__PTR51) );
  AND2_X1 U13904 ( .A1(_02682__PTR52), .A2(_02452__PTR0), .ZN(_02683__PTR52) );
  AND2_X1 U13905 ( .A1(_02682__PTR53), .A2(_02452__PTR0), .ZN(_02683__PTR53) );
  AND2_X1 U13906 ( .A1(_02682__PTR54), .A2(_02452__PTR0), .ZN(_02683__PTR54) );
  AND2_X1 U13907 ( .A1(_02682__PTR55), .A2(_02452__PTR0), .ZN(_02683__PTR55) );
  AND2_X1 U13908 ( .A1(_02682__PTR56), .A2(_02452__PTR0), .ZN(_02683__PTR56) );
  AND2_X1 U13909 ( .A1(_02682__PTR57), .A2(_02452__PTR0), .ZN(_02683__PTR57) );
  AND2_X1 U13910 ( .A1(_02682__PTR58), .A2(_02452__PTR0), .ZN(_02683__PTR58) );
  AND2_X1 U13911 ( .A1(_02682__PTR59), .A2(_02452__PTR0), .ZN(_02683__PTR59) );
  AND2_X1 U13912 ( .A1(_02682__PTR60), .A2(_02452__PTR0), .ZN(_02683__PTR60) );
  AND2_X1 U13913 ( .A1(_02682__PTR61), .A2(_02452__PTR0), .ZN(_02683__PTR61) );
  AND2_X1 U13914 ( .A1(_02682__PTR62), .A2(_02452__PTR0), .ZN(_02683__PTR62) );
  AND2_X1 U13915 ( .A1(_02682__PTR63), .A2(_02452__PTR0), .ZN(_02683__PTR63) );
  AND2_X1 U13916 ( .A1(_02682__PTR64), .A2(_02445__PTR2), .ZN(_02683__PTR64) );
  AND2_X1 U13917 ( .A1(_02682__PTR65), .A2(_02445__PTR2), .ZN(_02683__PTR65) );
  AND2_X1 U13918 ( .A1(_02682__PTR66), .A2(_02445__PTR2), .ZN(_02683__PTR66) );
  AND2_X1 U13919 ( .A1(_02682__PTR67), .A2(_02445__PTR2), .ZN(_02683__PTR67) );
  AND2_X1 U13920 ( .A1(_02682__PTR68), .A2(_02445__PTR2), .ZN(_02683__PTR68) );
  AND2_X1 U13921 ( .A1(_02682__PTR69), .A2(_02445__PTR2), .ZN(_02683__PTR69) );
  AND2_X1 U13922 ( .A1(_02682__PTR70), .A2(_02445__PTR2), .ZN(_02683__PTR70) );
  AND2_X1 U13923 ( .A1(_02682__PTR71), .A2(_02445__PTR2), .ZN(_02683__PTR71) );
  AND2_X1 U13924 ( .A1(_02682__PTR72), .A2(_02445__PTR2), .ZN(_02683__PTR72) );
  AND2_X1 U13925 ( .A1(_02682__PTR73), .A2(_02445__PTR2), .ZN(_02683__PTR73) );
  AND2_X1 U13926 ( .A1(_02682__PTR74), .A2(_02445__PTR2), .ZN(_02683__PTR74) );
  AND2_X1 U13927 ( .A1(_02682__PTR75), .A2(_02445__PTR2), .ZN(_02683__PTR75) );
  AND2_X1 U13928 ( .A1(_02682__PTR76), .A2(_02445__PTR2), .ZN(_02683__PTR76) );
  AND2_X1 U13929 ( .A1(_02682__PTR77), .A2(_02445__PTR2), .ZN(_02683__PTR77) );
  AND2_X1 U13930 ( .A1(_02682__PTR78), .A2(_02445__PTR2), .ZN(_02683__PTR78) );
  AND2_X1 U13931 ( .A1(_02682__PTR79), .A2(_02445__PTR2), .ZN(_02683__PTR79) );
  AND2_X1 U13932 ( .A1(_02682__PTR80), .A2(_02445__PTR2), .ZN(_02683__PTR80) );
  AND2_X1 U13933 ( .A1(_02682__PTR81), .A2(_02445__PTR2), .ZN(_02683__PTR81) );
  AND2_X1 U13934 ( .A1(_02682__PTR82), .A2(_02445__PTR2), .ZN(_02683__PTR82) );
  AND2_X1 U13935 ( .A1(_02682__PTR83), .A2(_02445__PTR2), .ZN(_02683__PTR83) );
  AND2_X1 U13936 ( .A1(_02682__PTR84), .A2(_02445__PTR2), .ZN(_02683__PTR84) );
  AND2_X1 U13937 ( .A1(_02682__PTR85), .A2(_02445__PTR2), .ZN(_02683__PTR85) );
  AND2_X1 U13938 ( .A1(_02682__PTR86), .A2(_02445__PTR2), .ZN(_02683__PTR86) );
  AND2_X1 U13939 ( .A1(_02682__PTR87), .A2(_02445__PTR2), .ZN(_02683__PTR87) );
  AND2_X1 U13940 ( .A1(_02682__PTR88), .A2(_02445__PTR2), .ZN(_02683__PTR88) );
  AND2_X1 U13941 ( .A1(_02682__PTR89), .A2(_02445__PTR2), .ZN(_02683__PTR89) );
  AND2_X1 U13942 ( .A1(_02682__PTR90), .A2(_02445__PTR2), .ZN(_02683__PTR90) );
  AND2_X1 U13943 ( .A1(_02682__PTR91), .A2(_02445__PTR2), .ZN(_02683__PTR91) );
  AND2_X1 U13944 ( .A1(_02682__PTR92), .A2(_02445__PTR2), .ZN(_02683__PTR92) );
  AND2_X1 U13945 ( .A1(_02682__PTR93), .A2(_02445__PTR2), .ZN(_02683__PTR93) );
  AND2_X1 U13946 ( .A1(_02682__PTR94), .A2(_02445__PTR2), .ZN(_02683__PTR94) );
  AND2_X1 U13947 ( .A1(_02682__PTR95), .A2(_02445__PTR2), .ZN(_02683__PTR95) );
  AND2_X1 U13948 ( .A1(_02682__PTR96), .A2(_02668__PTR4), .ZN(_02683__PTR96) );
  AND2_X1 U13949 ( .A1(_02682__PTR97), .A2(_02668__PTR4), .ZN(_02683__PTR97) );
  AND2_X1 U13950 ( .A1(_02682__PTR98), .A2(_02668__PTR4), .ZN(_02683__PTR98) );
  AND2_X1 U13951 ( .A1(_02682__PTR99), .A2(_02668__PTR4), .ZN(_02683__PTR99) );
  AND2_X1 U13952 ( .A1(_02682__PTR100), .A2(_02668__PTR4), .ZN(_02683__PTR100) );
  AND2_X1 U13953 ( .A1(_02682__PTR101), .A2(_02668__PTR4), .ZN(_02683__PTR101) );
  AND2_X1 U13954 ( .A1(_02682__PTR102), .A2(_02668__PTR4), .ZN(_02683__PTR102) );
  AND2_X1 U13955 ( .A1(_02682__PTR103), .A2(_02668__PTR4), .ZN(_02683__PTR103) );
  AND2_X1 U13956 ( .A1(_02682__PTR104), .A2(_02668__PTR4), .ZN(_02683__PTR104) );
  AND2_X1 U13957 ( .A1(_02682__PTR105), .A2(_02668__PTR4), .ZN(_02683__PTR105) );
  AND2_X1 U13958 ( .A1(_02682__PTR106), .A2(_02668__PTR4), .ZN(_02683__PTR106) );
  AND2_X1 U13959 ( .A1(_02682__PTR107), .A2(_02668__PTR4), .ZN(_02683__PTR107) );
  AND2_X1 U13960 ( .A1(_02682__PTR108), .A2(_02668__PTR4), .ZN(_02683__PTR108) );
  AND2_X1 U13961 ( .A1(_02682__PTR109), .A2(_02668__PTR4), .ZN(_02683__PTR109) );
  AND2_X1 U13962 ( .A1(_02682__PTR110), .A2(_02668__PTR4), .ZN(_02683__PTR110) );
  AND2_X1 U13963 ( .A1(_02682__PTR111), .A2(_02668__PTR4), .ZN(_02683__PTR111) );
  AND2_X1 U13964 ( .A1(_02682__PTR112), .A2(_02668__PTR4), .ZN(_02683__PTR112) );
  AND2_X1 U13965 ( .A1(_02682__PTR113), .A2(_02668__PTR4), .ZN(_02683__PTR113) );
  AND2_X1 U13966 ( .A1(_02682__PTR114), .A2(_02668__PTR4), .ZN(_02683__PTR114) );
  AND2_X1 U13967 ( .A1(_02682__PTR115), .A2(_02668__PTR4), .ZN(_02683__PTR115) );
  AND2_X1 U13968 ( .A1(_02682__PTR116), .A2(_02668__PTR4), .ZN(_02683__PTR116) );
  AND2_X1 U13969 ( .A1(_02682__PTR117), .A2(_02668__PTR4), .ZN(_02683__PTR117) );
  AND2_X1 U13970 ( .A1(_02682__PTR118), .A2(_02668__PTR4), .ZN(_02683__PTR118) );
  AND2_X1 U13971 ( .A1(_02682__PTR119), .A2(_02668__PTR4), .ZN(_02683__PTR119) );
  AND2_X1 U13972 ( .A1(_02682__PTR120), .A2(_02668__PTR4), .ZN(_02683__PTR120) );
  AND2_X1 U13973 ( .A1(_02682__PTR121), .A2(_02668__PTR4), .ZN(_02683__PTR121) );
  AND2_X1 U13974 ( .A1(_02682__PTR122), .A2(_02668__PTR4), .ZN(_02683__PTR122) );
  AND2_X1 U13975 ( .A1(_02682__PTR123), .A2(_02668__PTR4), .ZN(_02683__PTR123) );
  AND2_X1 U13976 ( .A1(_02682__PTR124), .A2(_02668__PTR4), .ZN(_02683__PTR124) );
  AND2_X1 U13977 ( .A1(_02682__PTR125), .A2(_02668__PTR4), .ZN(_02683__PTR125) );
  AND2_X1 U13978 ( .A1(_02682__PTR126), .A2(_02668__PTR4), .ZN(_02683__PTR126) );
  AND2_X1 U13979 ( .A1(_02682__PTR127), .A2(_02668__PTR4), .ZN(_02683__PTR127) );
  AND2_X1 U13980 ( .A1(_02662__PTR0), .A2(_02664__PTR0), .ZN(_02663__PTR0) );
  AND2_X1 U13981 ( .A1(_02662__PTR1), .A2(_02664__PTR0), .ZN(_02663__PTR1) );
  AND2_X1 U13982 ( .A1(_02662__PTR2), .A2(_02664__PTR0), .ZN(_02663__PTR2) );
  AND2_X1 U13983 ( .A1(_02662__PTR3), .A2(_02664__PTR0), .ZN(_02663__PTR3) );
  AND2_X1 U13984 ( .A1(_02662__PTR4), .A2(_02664__PTR0), .ZN(_02663__PTR4) );
  AND2_X1 U13985 ( .A1(_02662__PTR5), .A2(_02664__PTR0), .ZN(_02663__PTR5) );
  AND2_X1 U13986 ( .A1(_02662__PTR6), .A2(_02664__PTR0), .ZN(_02663__PTR6) );
  AND2_X1 U13987 ( .A1(_02662__PTR7), .A2(_02664__PTR0), .ZN(_02663__PTR7) );
  AND2_X1 U13988 ( .A1(_02662__PTR8), .A2(_02664__PTR0), .ZN(_02663__PTR8) );
  AND2_X1 U13989 ( .A1(_02662__PTR9), .A2(_02664__PTR0), .ZN(_02663__PTR9) );
  AND2_X1 U13990 ( .A1(_02662__PTR10), .A2(_02664__PTR0), .ZN(_02663__PTR10) );
  AND2_X1 U13991 ( .A1(_02662__PTR11), .A2(_02664__PTR0), .ZN(_02663__PTR11) );
  AND2_X1 U13992 ( .A1(_02662__PTR12), .A2(_02664__PTR0), .ZN(_02663__PTR12) );
  AND2_X1 U13993 ( .A1(_02662__PTR13), .A2(_02664__PTR0), .ZN(_02663__PTR13) );
  AND2_X1 U13994 ( .A1(_02662__PTR14), .A2(_02664__PTR0), .ZN(_02663__PTR14) );
  AND2_X1 U13995 ( .A1(_02662__PTR15), .A2(_02664__PTR0), .ZN(_02663__PTR15) );
  AND2_X1 U13996 ( .A1(_02662__PTR16), .A2(_02664__PTR0), .ZN(_02663__PTR16) );
  AND2_X1 U13997 ( .A1(_02662__PTR17), .A2(_02664__PTR0), .ZN(_02663__PTR17) );
  AND2_X1 U13998 ( .A1(_02662__PTR18), .A2(_02664__PTR0), .ZN(_02663__PTR18) );
  AND2_X1 U13999 ( .A1(_02662__PTR19), .A2(_02664__PTR0), .ZN(_02663__PTR19) );
  AND2_X1 U14000 ( .A1(_02662__PTR20), .A2(_02664__PTR0), .ZN(_02663__PTR20) );
  AND2_X1 U14001 ( .A1(_02662__PTR21), .A2(_02664__PTR0), .ZN(_02663__PTR21) );
  AND2_X1 U14002 ( .A1(_02662__PTR22), .A2(_02664__PTR0), .ZN(_02663__PTR22) );
  AND2_X1 U14003 ( .A1(_02662__PTR23), .A2(_02664__PTR0), .ZN(_02663__PTR23) );
  AND2_X1 U14004 ( .A1(_02662__PTR24), .A2(_02664__PTR0), .ZN(_02663__PTR24) );
  AND2_X1 U14005 ( .A1(_02662__PTR25), .A2(_02664__PTR0), .ZN(_02663__PTR25) );
  AND2_X1 U14006 ( .A1(_02662__PTR26), .A2(_02664__PTR0), .ZN(_02663__PTR26) );
  AND2_X1 U14007 ( .A1(_02662__PTR27), .A2(_02664__PTR0), .ZN(_02663__PTR27) );
  AND2_X1 U14008 ( .A1(_02662__PTR28), .A2(_02664__PTR0), .ZN(_02663__PTR28) );
  AND2_X1 U14009 ( .A1(_02662__PTR29), .A2(_02664__PTR0), .ZN(_02663__PTR29) );
  AND2_X1 U14010 ( .A1(_02662__PTR30), .A2(_02664__PTR0), .ZN(_02663__PTR30) );
  AND2_X1 U14011 ( .A1(_02662__PTR31), .A2(_02664__PTR0), .ZN(_02663__PTR31) );
  AND2_X1 U14012 ( .A1(P3_P1_InstAddrPointer_PTR0), .A2(_02664__PTR1), .ZN(_02663__PTR32) );
  AND2_X1 U14013 ( .A1(_02662__PTR33), .A2(_02664__PTR1), .ZN(_02663__PTR33) );
  AND2_X1 U14014 ( .A1(_02662__PTR34), .A2(_02664__PTR1), .ZN(_02663__PTR34) );
  AND2_X1 U14015 ( .A1(_02662__PTR35), .A2(_02664__PTR1), .ZN(_02663__PTR35) );
  AND2_X1 U14016 ( .A1(_02662__PTR36), .A2(_02664__PTR1), .ZN(_02663__PTR36) );
  AND2_X1 U14017 ( .A1(_02662__PTR37), .A2(_02664__PTR1), .ZN(_02663__PTR37) );
  AND2_X1 U14018 ( .A1(_02662__PTR38), .A2(_02664__PTR1), .ZN(_02663__PTR38) );
  AND2_X1 U14019 ( .A1(_02662__PTR39), .A2(_02664__PTR1), .ZN(_02663__PTR39) );
  AND2_X1 U14020 ( .A1(_02662__PTR40), .A2(_02664__PTR1), .ZN(_02663__PTR40) );
  AND2_X1 U14021 ( .A1(_02662__PTR41), .A2(_02664__PTR1), .ZN(_02663__PTR41) );
  AND2_X1 U14022 ( .A1(_02662__PTR42), .A2(_02664__PTR1), .ZN(_02663__PTR42) );
  AND2_X1 U14023 ( .A1(_02662__PTR43), .A2(_02664__PTR1), .ZN(_02663__PTR43) );
  AND2_X1 U14024 ( .A1(_02662__PTR44), .A2(_02664__PTR1), .ZN(_02663__PTR44) );
  AND2_X1 U14025 ( .A1(_02662__PTR45), .A2(_02664__PTR1), .ZN(_02663__PTR45) );
  AND2_X1 U14026 ( .A1(_02662__PTR46), .A2(_02664__PTR1), .ZN(_02663__PTR46) );
  AND2_X1 U14027 ( .A1(_02662__PTR47), .A2(_02664__PTR1), .ZN(_02663__PTR47) );
  AND2_X1 U14028 ( .A1(_02662__PTR48), .A2(_02664__PTR1), .ZN(_02663__PTR48) );
  AND2_X1 U14029 ( .A1(_02662__PTR49), .A2(_02664__PTR1), .ZN(_02663__PTR49) );
  AND2_X1 U14030 ( .A1(_02662__PTR50), .A2(_02664__PTR1), .ZN(_02663__PTR50) );
  AND2_X1 U14031 ( .A1(_02662__PTR51), .A2(_02664__PTR1), .ZN(_02663__PTR51) );
  AND2_X1 U14032 ( .A1(_02662__PTR52), .A2(_02664__PTR1), .ZN(_02663__PTR52) );
  AND2_X1 U14033 ( .A1(_02662__PTR53), .A2(_02664__PTR1), .ZN(_02663__PTR53) );
  AND2_X1 U14034 ( .A1(_02662__PTR54), .A2(_02664__PTR1), .ZN(_02663__PTR54) );
  AND2_X1 U14035 ( .A1(_02662__PTR55), .A2(_02664__PTR1), .ZN(_02663__PTR55) );
  AND2_X1 U14036 ( .A1(_02662__PTR56), .A2(_02664__PTR1), .ZN(_02663__PTR56) );
  AND2_X1 U14037 ( .A1(_02662__PTR57), .A2(_02664__PTR1), .ZN(_02663__PTR57) );
  AND2_X1 U14038 ( .A1(_02662__PTR58), .A2(_02664__PTR1), .ZN(_02663__PTR58) );
  AND2_X1 U14039 ( .A1(_02662__PTR59), .A2(_02664__PTR1), .ZN(_02663__PTR59) );
  AND2_X1 U14040 ( .A1(_02662__PTR60), .A2(_02664__PTR1), .ZN(_02663__PTR60) );
  AND2_X1 U14041 ( .A1(_02662__PTR61), .A2(_02664__PTR1), .ZN(_02663__PTR61) );
  AND2_X1 U14042 ( .A1(_02662__PTR62), .A2(_02664__PTR1), .ZN(_02663__PTR62) );
  AND2_X1 U14043 ( .A1(_02662__PTR63), .A2(_02664__PTR1), .ZN(_02663__PTR63) );
  AND2_X1 U14044 ( .A1(P3_P1_InstAddrPointer_PTR0), .A2(_02437__PTR0), .ZN(_02663__PTR64) );
  AND2_X1 U14045 ( .A1(_02662__PTR65), .A2(_02437__PTR0), .ZN(_02663__PTR65) );
  AND2_X1 U14046 ( .A1(_02662__PTR66), .A2(_02437__PTR0), .ZN(_02663__PTR66) );
  AND2_X1 U14047 ( .A1(_02662__PTR67), .A2(_02437__PTR0), .ZN(_02663__PTR67) );
  AND2_X1 U14048 ( .A1(_02662__PTR68), .A2(_02437__PTR0), .ZN(_02663__PTR68) );
  AND2_X1 U14049 ( .A1(_02662__PTR69), .A2(_02437__PTR0), .ZN(_02663__PTR69) );
  AND2_X1 U14050 ( .A1(_02662__PTR70), .A2(_02437__PTR0), .ZN(_02663__PTR70) );
  AND2_X1 U14051 ( .A1(_02662__PTR71), .A2(_02437__PTR0), .ZN(_02663__PTR71) );
  AND2_X1 U14052 ( .A1(_02662__PTR72), .A2(_02437__PTR0), .ZN(_02663__PTR72) );
  AND2_X1 U14053 ( .A1(_02662__PTR73), .A2(_02437__PTR0), .ZN(_02663__PTR73) );
  AND2_X1 U14054 ( .A1(_02662__PTR74), .A2(_02437__PTR0), .ZN(_02663__PTR74) );
  AND2_X1 U14055 ( .A1(_02662__PTR75), .A2(_02437__PTR0), .ZN(_02663__PTR75) );
  AND2_X1 U14056 ( .A1(_02662__PTR76), .A2(_02437__PTR0), .ZN(_02663__PTR76) );
  AND2_X1 U14057 ( .A1(_02662__PTR77), .A2(_02437__PTR0), .ZN(_02663__PTR77) );
  AND2_X1 U14058 ( .A1(_02662__PTR78), .A2(_02437__PTR0), .ZN(_02663__PTR78) );
  AND2_X1 U14059 ( .A1(_02662__PTR79), .A2(_02437__PTR0), .ZN(_02663__PTR79) );
  AND2_X1 U14060 ( .A1(_02662__PTR80), .A2(_02437__PTR0), .ZN(_02663__PTR80) );
  AND2_X1 U14061 ( .A1(_02662__PTR81), .A2(_02437__PTR0), .ZN(_02663__PTR81) );
  AND2_X1 U14062 ( .A1(_02662__PTR82), .A2(_02437__PTR0), .ZN(_02663__PTR82) );
  AND2_X1 U14063 ( .A1(_02662__PTR83), .A2(_02437__PTR0), .ZN(_02663__PTR83) );
  AND2_X1 U14064 ( .A1(_02662__PTR84), .A2(_02437__PTR0), .ZN(_02663__PTR84) );
  AND2_X1 U14065 ( .A1(_02662__PTR85), .A2(_02437__PTR0), .ZN(_02663__PTR85) );
  AND2_X1 U14066 ( .A1(_02662__PTR86), .A2(_02437__PTR0), .ZN(_02663__PTR86) );
  AND2_X1 U14067 ( .A1(_02662__PTR87), .A2(_02437__PTR0), .ZN(_02663__PTR87) );
  AND2_X1 U14068 ( .A1(_02662__PTR88), .A2(_02437__PTR0), .ZN(_02663__PTR88) );
  AND2_X1 U14069 ( .A1(_02662__PTR89), .A2(_02437__PTR0), .ZN(_02663__PTR89) );
  AND2_X1 U14070 ( .A1(_02662__PTR90), .A2(_02437__PTR0), .ZN(_02663__PTR90) );
  AND2_X1 U14071 ( .A1(_02662__PTR91), .A2(_02437__PTR0), .ZN(_02663__PTR91) );
  AND2_X1 U14072 ( .A1(_02662__PTR92), .A2(_02437__PTR0), .ZN(_02663__PTR92) );
  AND2_X1 U14073 ( .A1(_02662__PTR93), .A2(_02437__PTR0), .ZN(_02663__PTR93) );
  AND2_X1 U14074 ( .A1(_02662__PTR94), .A2(_02437__PTR0), .ZN(_02663__PTR94) );
  AND2_X1 U14075 ( .A1(_02662__PTR95), .A2(_02437__PTR0), .ZN(_02663__PTR95) );
  AND2_X1 U14076 ( .A1(P3_P1_InstAddrPointer_PTR0), .A2(_02437__PTR1), .ZN(_02663__PTR96) );
  AND2_X1 U14077 ( .A1(_02662__PTR97), .A2(_02437__PTR1), .ZN(_02663__PTR97) );
  AND2_X1 U14078 ( .A1(_02662__PTR98), .A2(_02437__PTR1), .ZN(_02663__PTR98) );
  AND2_X1 U14079 ( .A1(_02662__PTR99), .A2(_02437__PTR1), .ZN(_02663__PTR99) );
  AND2_X1 U14080 ( .A1(_02662__PTR100), .A2(_02437__PTR1), .ZN(_02663__PTR100) );
  AND2_X1 U14081 ( .A1(_02662__PTR101), .A2(_02437__PTR1), .ZN(_02663__PTR101) );
  AND2_X1 U14082 ( .A1(_02662__PTR102), .A2(_02437__PTR1), .ZN(_02663__PTR102) );
  AND2_X1 U14083 ( .A1(_02662__PTR103), .A2(_02437__PTR1), .ZN(_02663__PTR103) );
  AND2_X1 U14084 ( .A1(_02662__PTR104), .A2(_02437__PTR1), .ZN(_02663__PTR104) );
  AND2_X1 U14085 ( .A1(_02662__PTR105), .A2(_02437__PTR1), .ZN(_02663__PTR105) );
  AND2_X1 U14086 ( .A1(_02662__PTR106), .A2(_02437__PTR1), .ZN(_02663__PTR106) );
  AND2_X1 U14087 ( .A1(_02662__PTR107), .A2(_02437__PTR1), .ZN(_02663__PTR107) );
  AND2_X1 U14088 ( .A1(_02662__PTR108), .A2(_02437__PTR1), .ZN(_02663__PTR108) );
  AND2_X1 U14089 ( .A1(_02662__PTR109), .A2(_02437__PTR1), .ZN(_02663__PTR109) );
  AND2_X1 U14090 ( .A1(_02662__PTR110), .A2(_02437__PTR1), .ZN(_02663__PTR110) );
  AND2_X1 U14091 ( .A1(_02662__PTR111), .A2(_02437__PTR1), .ZN(_02663__PTR111) );
  AND2_X1 U14092 ( .A1(_02662__PTR112), .A2(_02437__PTR1), .ZN(_02663__PTR112) );
  AND2_X1 U14093 ( .A1(_02662__PTR113), .A2(_02437__PTR1), .ZN(_02663__PTR113) );
  AND2_X1 U14094 ( .A1(_02662__PTR114), .A2(_02437__PTR1), .ZN(_02663__PTR114) );
  AND2_X1 U14095 ( .A1(_02662__PTR115), .A2(_02437__PTR1), .ZN(_02663__PTR115) );
  AND2_X1 U14096 ( .A1(_02662__PTR116), .A2(_02437__PTR1), .ZN(_02663__PTR116) );
  AND2_X1 U14097 ( .A1(_02662__PTR117), .A2(_02437__PTR1), .ZN(_02663__PTR117) );
  AND2_X1 U14098 ( .A1(_02662__PTR118), .A2(_02437__PTR1), .ZN(_02663__PTR118) );
  AND2_X1 U14099 ( .A1(_02662__PTR119), .A2(_02437__PTR1), .ZN(_02663__PTR119) );
  AND2_X1 U14100 ( .A1(_02662__PTR120), .A2(_02437__PTR1), .ZN(_02663__PTR120) );
  AND2_X1 U14101 ( .A1(_02662__PTR121), .A2(_02437__PTR1), .ZN(_02663__PTR121) );
  AND2_X1 U14102 ( .A1(_02662__PTR122), .A2(_02437__PTR1), .ZN(_02663__PTR122) );
  AND2_X1 U14103 ( .A1(_02662__PTR123), .A2(_02437__PTR1), .ZN(_02663__PTR123) );
  AND2_X1 U14104 ( .A1(_02662__PTR124), .A2(_02437__PTR1), .ZN(_02663__PTR124) );
  AND2_X1 U14105 ( .A1(_02662__PTR125), .A2(_02437__PTR1), .ZN(_02663__PTR125) );
  AND2_X1 U14106 ( .A1(_02662__PTR126), .A2(_02437__PTR1), .ZN(_02663__PTR126) );
  AND2_X1 U14107 ( .A1(_02662__PTR127), .A2(_02437__PTR1), .ZN(_02663__PTR127) );
  AND2_X1 U14108 ( .A1(_02662__PTR128), .A2(_02664__PTR4), .ZN(_02663__PTR128) );
  AND2_X1 U14109 ( .A1(_02662__PTR129), .A2(_02664__PTR4), .ZN(_02663__PTR129) );
  AND2_X1 U14110 ( .A1(_02662__PTR130), .A2(_02664__PTR4), .ZN(_02663__PTR130) );
  AND2_X1 U14111 ( .A1(_02662__PTR131), .A2(_02664__PTR4), .ZN(_02663__PTR131) );
  AND2_X1 U14112 ( .A1(_02662__PTR132), .A2(_02664__PTR4), .ZN(_02663__PTR132) );
  AND2_X1 U14113 ( .A1(_02662__PTR133), .A2(_02664__PTR4), .ZN(_02663__PTR133) );
  AND2_X1 U14114 ( .A1(_02662__PTR134), .A2(_02664__PTR4), .ZN(_02663__PTR134) );
  AND2_X1 U14115 ( .A1(_02662__PTR135), .A2(_02664__PTR4), .ZN(_02663__PTR135) );
  AND2_X1 U14116 ( .A1(_02662__PTR136), .A2(_02664__PTR4), .ZN(_02663__PTR136) );
  AND2_X1 U14117 ( .A1(_02662__PTR137), .A2(_02664__PTR4), .ZN(_02663__PTR137) );
  AND2_X1 U14118 ( .A1(_02662__PTR138), .A2(_02664__PTR4), .ZN(_02663__PTR138) );
  AND2_X1 U14119 ( .A1(_02662__PTR139), .A2(_02664__PTR4), .ZN(_02663__PTR139) );
  AND2_X1 U14120 ( .A1(_02662__PTR140), .A2(_02664__PTR4), .ZN(_02663__PTR140) );
  AND2_X1 U14121 ( .A1(_02662__PTR141), .A2(_02664__PTR4), .ZN(_02663__PTR141) );
  AND2_X1 U14122 ( .A1(_02662__PTR142), .A2(_02664__PTR4), .ZN(_02663__PTR142) );
  AND2_X1 U14123 ( .A1(_02662__PTR143), .A2(_02664__PTR4), .ZN(_02663__PTR143) );
  AND2_X1 U14124 ( .A1(_02662__PTR144), .A2(_02664__PTR4), .ZN(_02663__PTR144) );
  AND2_X1 U14125 ( .A1(_02662__PTR145), .A2(_02664__PTR4), .ZN(_02663__PTR145) );
  AND2_X1 U14126 ( .A1(_02662__PTR146), .A2(_02664__PTR4), .ZN(_02663__PTR146) );
  AND2_X1 U14127 ( .A1(_02662__PTR147), .A2(_02664__PTR4), .ZN(_02663__PTR147) );
  AND2_X1 U14128 ( .A1(_02662__PTR148), .A2(_02664__PTR4), .ZN(_02663__PTR148) );
  AND2_X1 U14129 ( .A1(_02662__PTR149), .A2(_02664__PTR4), .ZN(_02663__PTR149) );
  AND2_X1 U14130 ( .A1(_02662__PTR150), .A2(_02664__PTR4), .ZN(_02663__PTR150) );
  AND2_X1 U14131 ( .A1(_02662__PTR151), .A2(_02664__PTR4), .ZN(_02663__PTR151) );
  AND2_X1 U14132 ( .A1(_02662__PTR152), .A2(_02664__PTR4), .ZN(_02663__PTR152) );
  AND2_X1 U14133 ( .A1(_02662__PTR153), .A2(_02664__PTR4), .ZN(_02663__PTR153) );
  AND2_X1 U14134 ( .A1(_02662__PTR154), .A2(_02664__PTR4), .ZN(_02663__PTR154) );
  AND2_X1 U14135 ( .A1(_02662__PTR155), .A2(_02664__PTR4), .ZN(_02663__PTR155) );
  AND2_X1 U14136 ( .A1(_02662__PTR156), .A2(_02664__PTR4), .ZN(_02663__PTR156) );
  AND2_X1 U14137 ( .A1(_02662__PTR157), .A2(_02664__PTR4), .ZN(_02663__PTR157) );
  AND2_X1 U14138 ( .A1(_02662__PTR158), .A2(_02664__PTR4), .ZN(_02663__PTR158) );
  AND2_X1 U14139 ( .A1(_02662__PTR159), .A2(_02664__PTR4), .ZN(_02663__PTR159) );
  AND2_X1 U14140 ( .A1(_02662__PTR160), .A2(_02437__PTR2), .ZN(_02663__PTR160) );
  AND2_X1 U14141 ( .A1(_02662__PTR161), .A2(_02437__PTR2), .ZN(_02663__PTR161) );
  AND2_X1 U14142 ( .A1(_02662__PTR162), .A2(_02437__PTR2), .ZN(_02663__PTR162) );
  AND2_X1 U14143 ( .A1(_02662__PTR163), .A2(_02437__PTR2), .ZN(_02663__PTR163) );
  AND2_X1 U14144 ( .A1(_02662__PTR164), .A2(_02437__PTR2), .ZN(_02663__PTR164) );
  AND2_X1 U14145 ( .A1(_02662__PTR165), .A2(_02437__PTR2), .ZN(_02663__PTR165) );
  AND2_X1 U14146 ( .A1(_02662__PTR166), .A2(_02437__PTR2), .ZN(_02663__PTR166) );
  AND2_X1 U14147 ( .A1(_02662__PTR167), .A2(_02437__PTR2), .ZN(_02663__PTR167) );
  AND2_X1 U14148 ( .A1(_02662__PTR168), .A2(_02437__PTR2), .ZN(_02663__PTR168) );
  AND2_X1 U14149 ( .A1(_02662__PTR169), .A2(_02437__PTR2), .ZN(_02663__PTR169) );
  AND2_X1 U14150 ( .A1(_02662__PTR170), .A2(_02437__PTR2), .ZN(_02663__PTR170) );
  AND2_X1 U14151 ( .A1(_02662__PTR171), .A2(_02437__PTR2), .ZN(_02663__PTR171) );
  AND2_X1 U14152 ( .A1(_02662__PTR172), .A2(_02437__PTR2), .ZN(_02663__PTR172) );
  AND2_X1 U14153 ( .A1(_02662__PTR173), .A2(_02437__PTR2), .ZN(_02663__PTR173) );
  AND2_X1 U14154 ( .A1(_02662__PTR174), .A2(_02437__PTR2), .ZN(_02663__PTR174) );
  AND2_X1 U14155 ( .A1(_02662__PTR175), .A2(_02437__PTR2), .ZN(_02663__PTR175) );
  AND2_X1 U14156 ( .A1(_02662__PTR176), .A2(_02437__PTR2), .ZN(_02663__PTR176) );
  AND2_X1 U14157 ( .A1(_02662__PTR177), .A2(_02437__PTR2), .ZN(_02663__PTR177) );
  AND2_X1 U14158 ( .A1(_02662__PTR178), .A2(_02437__PTR2), .ZN(_02663__PTR178) );
  AND2_X1 U14159 ( .A1(_02662__PTR179), .A2(_02437__PTR2), .ZN(_02663__PTR179) );
  AND2_X1 U14160 ( .A1(_02662__PTR180), .A2(_02437__PTR2), .ZN(_02663__PTR180) );
  AND2_X1 U14161 ( .A1(_02662__PTR181), .A2(_02437__PTR2), .ZN(_02663__PTR181) );
  AND2_X1 U14162 ( .A1(_02662__PTR182), .A2(_02437__PTR2), .ZN(_02663__PTR182) );
  AND2_X1 U14163 ( .A1(_02662__PTR183), .A2(_02437__PTR2), .ZN(_02663__PTR183) );
  AND2_X1 U14164 ( .A1(_02662__PTR184), .A2(_02437__PTR2), .ZN(_02663__PTR184) );
  AND2_X1 U14165 ( .A1(_02662__PTR185), .A2(_02437__PTR2), .ZN(_02663__PTR185) );
  AND2_X1 U14166 ( .A1(_02662__PTR186), .A2(_02437__PTR2), .ZN(_02663__PTR186) );
  AND2_X1 U14167 ( .A1(_02662__PTR187), .A2(_02437__PTR2), .ZN(_02663__PTR187) );
  AND2_X1 U14168 ( .A1(_02662__PTR188), .A2(_02437__PTR2), .ZN(_02663__PTR188) );
  AND2_X1 U14169 ( .A1(_02662__PTR189), .A2(_02437__PTR2), .ZN(_02663__PTR189) );
  AND2_X1 U14170 ( .A1(_02662__PTR190), .A2(_02437__PTR2), .ZN(_02663__PTR190) );
  AND2_X1 U14171 ( .A1(_02662__PTR191), .A2(_02437__PTR2), .ZN(_02663__PTR191) );
  AND2_X1 U14172 ( .A1(_02662__PTR192), .A2(_02437__PTR3), .ZN(_02663__PTR192) );
  AND2_X1 U14173 ( .A1(_02662__PTR193), .A2(_02437__PTR3), .ZN(_02663__PTR193) );
  AND2_X1 U14174 ( .A1(_02662__PTR194), .A2(_02437__PTR3), .ZN(_02663__PTR194) );
  AND2_X1 U14175 ( .A1(_02662__PTR195), .A2(_02437__PTR3), .ZN(_02663__PTR195) );
  AND2_X1 U14176 ( .A1(_02662__PTR196), .A2(_02437__PTR3), .ZN(_02663__PTR196) );
  AND2_X1 U14177 ( .A1(_02662__PTR197), .A2(_02437__PTR3), .ZN(_02663__PTR197) );
  AND2_X1 U14178 ( .A1(_02662__PTR198), .A2(_02437__PTR3), .ZN(_02663__PTR198) );
  AND2_X1 U14179 ( .A1(_02662__PTR199), .A2(_02437__PTR3), .ZN(_02663__PTR199) );
  AND2_X1 U14180 ( .A1(_02662__PTR200), .A2(_02437__PTR3), .ZN(_02663__PTR200) );
  AND2_X1 U14181 ( .A1(_02662__PTR201), .A2(_02437__PTR3), .ZN(_02663__PTR201) );
  AND2_X1 U14182 ( .A1(_02662__PTR202), .A2(_02437__PTR3), .ZN(_02663__PTR202) );
  AND2_X1 U14183 ( .A1(_02662__PTR203), .A2(_02437__PTR3), .ZN(_02663__PTR203) );
  AND2_X1 U14184 ( .A1(_02662__PTR204), .A2(_02437__PTR3), .ZN(_02663__PTR204) );
  AND2_X1 U14185 ( .A1(_02662__PTR205), .A2(_02437__PTR3), .ZN(_02663__PTR205) );
  AND2_X1 U14186 ( .A1(_02662__PTR206), .A2(_02437__PTR3), .ZN(_02663__PTR206) );
  AND2_X1 U14187 ( .A1(_02662__PTR207), .A2(_02437__PTR3), .ZN(_02663__PTR207) );
  AND2_X1 U14188 ( .A1(_02662__PTR208), .A2(_02437__PTR3), .ZN(_02663__PTR208) );
  AND2_X1 U14189 ( .A1(_02662__PTR209), .A2(_02437__PTR3), .ZN(_02663__PTR209) );
  AND2_X1 U14190 ( .A1(_02662__PTR210), .A2(_02437__PTR3), .ZN(_02663__PTR210) );
  AND2_X1 U14191 ( .A1(_02662__PTR211), .A2(_02437__PTR3), .ZN(_02663__PTR211) );
  AND2_X1 U14192 ( .A1(_02662__PTR212), .A2(_02437__PTR3), .ZN(_02663__PTR212) );
  AND2_X1 U14193 ( .A1(_02662__PTR213), .A2(_02437__PTR3), .ZN(_02663__PTR213) );
  AND2_X1 U14194 ( .A1(_02662__PTR214), .A2(_02437__PTR3), .ZN(_02663__PTR214) );
  AND2_X1 U14195 ( .A1(_02662__PTR215), .A2(_02437__PTR3), .ZN(_02663__PTR215) );
  AND2_X1 U14196 ( .A1(_02662__PTR216), .A2(_02437__PTR3), .ZN(_02663__PTR216) );
  AND2_X1 U14197 ( .A1(_02662__PTR217), .A2(_02437__PTR3), .ZN(_02663__PTR217) );
  AND2_X1 U14198 ( .A1(_02662__PTR218), .A2(_02437__PTR3), .ZN(_02663__PTR218) );
  AND2_X1 U14199 ( .A1(_02662__PTR219), .A2(_02437__PTR3), .ZN(_02663__PTR219) );
  AND2_X1 U14200 ( .A1(_02662__PTR220), .A2(_02437__PTR3), .ZN(_02663__PTR220) );
  AND2_X1 U14201 ( .A1(_02662__PTR221), .A2(_02437__PTR3), .ZN(_02663__PTR221) );
  AND2_X1 U14202 ( .A1(_02662__PTR222), .A2(_02437__PTR3), .ZN(_02663__PTR222) );
  AND2_X1 U14203 ( .A1(_02662__PTR223), .A2(_02437__PTR3), .ZN(_02663__PTR223) );
  AND2_X1 U14204 ( .A1(P3_P1_PhyAddrPointer_PTR0), .A2(_02672__PTR0), .ZN(_02671__PTR0) );
  AND2_X1 U14205 ( .A1(P3_P1_PhyAddrPointer_PTR1), .A2(_02672__PTR0), .ZN(_02671__PTR1) );
  AND2_X1 U14206 ( .A1(P3_P1_PhyAddrPointer_PTR2), .A2(_02672__PTR0), .ZN(_02671__PTR2) );
  AND2_X1 U14207 ( .A1(P3_P1_PhyAddrPointer_PTR3), .A2(_02672__PTR0), .ZN(_02671__PTR3) );
  AND2_X1 U14208 ( .A1(P3_P1_PhyAddrPointer_PTR4), .A2(_02672__PTR0), .ZN(_02671__PTR4) );
  AND2_X1 U14209 ( .A1(P3_P1_PhyAddrPointer_PTR5), .A2(_02672__PTR0), .ZN(_02671__PTR5) );
  AND2_X1 U14210 ( .A1(P3_P1_PhyAddrPointer_PTR6), .A2(_02672__PTR0), .ZN(_02671__PTR6) );
  AND2_X1 U14211 ( .A1(P3_P1_PhyAddrPointer_PTR7), .A2(_02672__PTR0), .ZN(_02671__PTR7) );
  AND2_X1 U14212 ( .A1(P3_P1_PhyAddrPointer_PTR8), .A2(_02672__PTR0), .ZN(_02671__PTR8) );
  AND2_X1 U14213 ( .A1(P3_P1_PhyAddrPointer_PTR9), .A2(_02672__PTR0), .ZN(_02671__PTR9) );
  AND2_X1 U14214 ( .A1(P3_P1_PhyAddrPointer_PTR10), .A2(_02672__PTR0), .ZN(_02671__PTR10) );
  AND2_X1 U14215 ( .A1(P3_P1_PhyAddrPointer_PTR11), .A2(_02672__PTR0), .ZN(_02671__PTR11) );
  AND2_X1 U14216 ( .A1(P3_P1_PhyAddrPointer_PTR12), .A2(_02672__PTR0), .ZN(_02671__PTR12) );
  AND2_X1 U14217 ( .A1(P3_P1_PhyAddrPointer_PTR13), .A2(_02672__PTR0), .ZN(_02671__PTR13) );
  AND2_X1 U14218 ( .A1(P3_P1_PhyAddrPointer_PTR14), .A2(_02672__PTR0), .ZN(_02671__PTR14) );
  AND2_X1 U14219 ( .A1(P3_P1_PhyAddrPointer_PTR15), .A2(_02672__PTR0), .ZN(_02671__PTR15) );
  AND2_X1 U14220 ( .A1(P3_P1_PhyAddrPointer_PTR16), .A2(_02672__PTR0), .ZN(_02671__PTR16) );
  AND2_X1 U14221 ( .A1(P3_P1_PhyAddrPointer_PTR17), .A2(_02672__PTR0), .ZN(_02671__PTR17) );
  AND2_X1 U14222 ( .A1(P3_P1_PhyAddrPointer_PTR18), .A2(_02672__PTR0), .ZN(_02671__PTR18) );
  AND2_X1 U14223 ( .A1(P3_P1_PhyAddrPointer_PTR19), .A2(_02672__PTR0), .ZN(_02671__PTR19) );
  AND2_X1 U14224 ( .A1(P3_P1_PhyAddrPointer_PTR20), .A2(_02672__PTR0), .ZN(_02671__PTR20) );
  AND2_X1 U14225 ( .A1(P3_P1_PhyAddrPointer_PTR21), .A2(_02672__PTR0), .ZN(_02671__PTR21) );
  AND2_X1 U14226 ( .A1(P3_P1_PhyAddrPointer_PTR22), .A2(_02672__PTR0), .ZN(_02671__PTR22) );
  AND2_X1 U14227 ( .A1(P3_P1_PhyAddrPointer_PTR23), .A2(_02672__PTR0), .ZN(_02671__PTR23) );
  AND2_X1 U14228 ( .A1(P3_P1_PhyAddrPointer_PTR24), .A2(_02672__PTR0), .ZN(_02671__PTR24) );
  AND2_X1 U14229 ( .A1(P3_P1_PhyAddrPointer_PTR25), .A2(_02672__PTR0), .ZN(_02671__PTR25) );
  AND2_X1 U14230 ( .A1(P3_P1_PhyAddrPointer_PTR26), .A2(_02672__PTR0), .ZN(_02671__PTR26) );
  AND2_X1 U14231 ( .A1(P3_P1_PhyAddrPointer_PTR27), .A2(_02672__PTR0), .ZN(_02671__PTR27) );
  AND2_X1 U14232 ( .A1(P3_P1_PhyAddrPointer_PTR28), .A2(_02672__PTR0), .ZN(_02671__PTR28) );
  AND2_X1 U14233 ( .A1(P3_P1_PhyAddrPointer_PTR29), .A2(_02672__PTR0), .ZN(_02671__PTR29) );
  AND2_X1 U14234 ( .A1(P3_P1_PhyAddrPointer_PTR30), .A2(_02672__PTR0), .ZN(_02671__PTR30) );
  AND2_X1 U14235 ( .A1(P3_P1_PhyAddrPointer_PTR31), .A2(_02672__PTR0), .ZN(_02671__PTR31) );
  AND2_X1 U14236 ( .A1(_02670__PTR32), .A2(_02437__PTR2), .ZN(_02671__PTR32) );
  AND2_X1 U14237 ( .A1(_02670__PTR33), .A2(_02437__PTR2), .ZN(_02671__PTR33) );
  AND2_X1 U14238 ( .A1(_02670__PTR34), .A2(_02437__PTR2), .ZN(_02671__PTR34) );
  AND2_X1 U14239 ( .A1(_02670__PTR35), .A2(_02437__PTR2), .ZN(_02671__PTR35) );
  AND2_X1 U14240 ( .A1(_02670__PTR36), .A2(_02437__PTR2), .ZN(_02671__PTR36) );
  AND2_X1 U14241 ( .A1(_02670__PTR37), .A2(_02437__PTR2), .ZN(_02671__PTR37) );
  AND2_X1 U14242 ( .A1(_02670__PTR38), .A2(_02437__PTR2), .ZN(_02671__PTR38) );
  AND2_X1 U14243 ( .A1(_02670__PTR39), .A2(_02437__PTR2), .ZN(_02671__PTR39) );
  AND2_X1 U14244 ( .A1(_02670__PTR40), .A2(_02437__PTR2), .ZN(_02671__PTR40) );
  AND2_X1 U14245 ( .A1(_02670__PTR41), .A2(_02437__PTR2), .ZN(_02671__PTR41) );
  AND2_X1 U14246 ( .A1(_02670__PTR42), .A2(_02437__PTR2), .ZN(_02671__PTR42) );
  AND2_X1 U14247 ( .A1(_02670__PTR43), .A2(_02437__PTR2), .ZN(_02671__PTR43) );
  AND2_X1 U14248 ( .A1(_02670__PTR44), .A2(_02437__PTR2), .ZN(_02671__PTR44) );
  AND2_X1 U14249 ( .A1(_02670__PTR45), .A2(_02437__PTR2), .ZN(_02671__PTR45) );
  AND2_X1 U14250 ( .A1(_02670__PTR46), .A2(_02437__PTR2), .ZN(_02671__PTR46) );
  AND2_X1 U14251 ( .A1(_02670__PTR47), .A2(_02437__PTR2), .ZN(_02671__PTR47) );
  AND2_X1 U14252 ( .A1(_02670__PTR48), .A2(_02437__PTR2), .ZN(_02671__PTR48) );
  AND2_X1 U14253 ( .A1(_02670__PTR49), .A2(_02437__PTR2), .ZN(_02671__PTR49) );
  AND2_X1 U14254 ( .A1(_02670__PTR50), .A2(_02437__PTR2), .ZN(_02671__PTR50) );
  AND2_X1 U14255 ( .A1(_02670__PTR51), .A2(_02437__PTR2), .ZN(_02671__PTR51) );
  AND2_X1 U14256 ( .A1(_02670__PTR52), .A2(_02437__PTR2), .ZN(_02671__PTR52) );
  AND2_X1 U14257 ( .A1(_02670__PTR53), .A2(_02437__PTR2), .ZN(_02671__PTR53) );
  AND2_X1 U14258 ( .A1(_02670__PTR54), .A2(_02437__PTR2), .ZN(_02671__PTR54) );
  AND2_X1 U14259 ( .A1(_02670__PTR55), .A2(_02437__PTR2), .ZN(_02671__PTR55) );
  AND2_X1 U14260 ( .A1(_02670__PTR56), .A2(_02437__PTR2), .ZN(_02671__PTR56) );
  AND2_X1 U14261 ( .A1(_02670__PTR57), .A2(_02437__PTR2), .ZN(_02671__PTR57) );
  AND2_X1 U14262 ( .A1(_02670__PTR58), .A2(_02437__PTR2), .ZN(_02671__PTR58) );
  AND2_X1 U14263 ( .A1(_02670__PTR59), .A2(_02437__PTR2), .ZN(_02671__PTR59) );
  AND2_X1 U14264 ( .A1(_02670__PTR60), .A2(_02437__PTR2), .ZN(_02671__PTR60) );
  AND2_X1 U14265 ( .A1(_02670__PTR61), .A2(_02437__PTR2), .ZN(_02671__PTR61) );
  AND2_X1 U14266 ( .A1(_02670__PTR62), .A2(_02437__PTR2), .ZN(_02671__PTR62) );
  AND2_X1 U14267 ( .A1(_02670__PTR63), .A2(_02437__PTR2), .ZN(_02671__PTR63) );
  AND2_X1 U14268 ( .A1(_02670__PTR64), .A2(_02437__PTR3), .ZN(_02671__PTR64) );
  AND2_X1 U14269 ( .A1(_02670__PTR65), .A2(_02437__PTR3), .ZN(_02671__PTR65) );
  AND2_X1 U14270 ( .A1(_02670__PTR66), .A2(_02437__PTR3), .ZN(_02671__PTR66) );
  AND2_X1 U14271 ( .A1(_02670__PTR67), .A2(_02437__PTR3), .ZN(_02671__PTR67) );
  AND2_X1 U14272 ( .A1(_02670__PTR68), .A2(_02437__PTR3), .ZN(_02671__PTR68) );
  AND2_X1 U14273 ( .A1(_02670__PTR69), .A2(_02437__PTR3), .ZN(_02671__PTR69) );
  AND2_X1 U14274 ( .A1(_02670__PTR70), .A2(_02437__PTR3), .ZN(_02671__PTR70) );
  AND2_X1 U14275 ( .A1(_02670__PTR71), .A2(_02437__PTR3), .ZN(_02671__PTR71) );
  AND2_X1 U14276 ( .A1(_02670__PTR72), .A2(_02437__PTR3), .ZN(_02671__PTR72) );
  AND2_X1 U14277 ( .A1(_02670__PTR73), .A2(_02437__PTR3), .ZN(_02671__PTR73) );
  AND2_X1 U14278 ( .A1(_02670__PTR74), .A2(_02437__PTR3), .ZN(_02671__PTR74) );
  AND2_X1 U14279 ( .A1(_02670__PTR75), .A2(_02437__PTR3), .ZN(_02671__PTR75) );
  AND2_X1 U14280 ( .A1(_02670__PTR76), .A2(_02437__PTR3), .ZN(_02671__PTR76) );
  AND2_X1 U14281 ( .A1(_02670__PTR77), .A2(_02437__PTR3), .ZN(_02671__PTR77) );
  AND2_X1 U14282 ( .A1(_02670__PTR78), .A2(_02437__PTR3), .ZN(_02671__PTR78) );
  AND2_X1 U14283 ( .A1(_02670__PTR79), .A2(_02437__PTR3), .ZN(_02671__PTR79) );
  AND2_X1 U14284 ( .A1(_02670__PTR80), .A2(_02437__PTR3), .ZN(_02671__PTR80) );
  AND2_X1 U14285 ( .A1(_02670__PTR81), .A2(_02437__PTR3), .ZN(_02671__PTR81) );
  AND2_X1 U14286 ( .A1(_02670__PTR82), .A2(_02437__PTR3), .ZN(_02671__PTR82) );
  AND2_X1 U14287 ( .A1(_02670__PTR83), .A2(_02437__PTR3), .ZN(_02671__PTR83) );
  AND2_X1 U14288 ( .A1(_02670__PTR84), .A2(_02437__PTR3), .ZN(_02671__PTR84) );
  AND2_X1 U14289 ( .A1(_02670__PTR85), .A2(_02437__PTR3), .ZN(_02671__PTR85) );
  AND2_X1 U14290 ( .A1(_02670__PTR86), .A2(_02437__PTR3), .ZN(_02671__PTR86) );
  AND2_X1 U14291 ( .A1(_02670__PTR87), .A2(_02437__PTR3), .ZN(_02671__PTR87) );
  AND2_X1 U14292 ( .A1(_02670__PTR88), .A2(_02437__PTR3), .ZN(_02671__PTR88) );
  AND2_X1 U14293 ( .A1(_02670__PTR89), .A2(_02437__PTR3), .ZN(_02671__PTR89) );
  AND2_X1 U14294 ( .A1(_02670__PTR90), .A2(_02437__PTR3), .ZN(_02671__PTR90) );
  AND2_X1 U14295 ( .A1(_02670__PTR91), .A2(_02437__PTR3), .ZN(_02671__PTR91) );
  AND2_X1 U14296 ( .A1(_02670__PTR92), .A2(_02437__PTR3), .ZN(_02671__PTR92) );
  AND2_X1 U14297 ( .A1(_02670__PTR93), .A2(_02437__PTR3), .ZN(_02671__PTR93) );
  AND2_X1 U14298 ( .A1(_02670__PTR94), .A2(_02437__PTR3), .ZN(_02671__PTR94) );
  AND2_X1 U14299 ( .A1(_02670__PTR95), .A2(_02437__PTR3), .ZN(_02671__PTR95) );
  AND2_X1 U14300 ( .A1(P3_P1_State2_PTR0), .A2(_02698__PTR0), .ZN(_02697__PTR0) );
  AND2_X1 U14301 ( .A1(P3_P1_State2_PTR1), .A2(_02698__PTR0), .ZN(_02697__PTR1) );
  AND2_X1 U14302 ( .A1(P3_P1_State2_PTR2), .A2(_02698__PTR0), .ZN(_02697__PTR2) );
  AND2_X1 U14303 ( .A1(P3_P1_State2_PTR3), .A2(_02698__PTR0), .ZN(_02697__PTR3) );
  AND2_X1 U14304 ( .A1(_02696__PTR4), .A2(_02445__PTR2), .ZN(_02697__PTR4) );
  AND2_X1 U14305 ( .A1(_02696__PTR5), .A2(_02445__PTR2), .ZN(_02697__PTR5) );
  AND2_X1 U14306 ( .A1(_02696__PTR6), .A2(_02445__PTR2), .ZN(_02697__PTR6) );
  AND2_X1 U14307 ( .A1(_02696__PTR7), .A2(_02445__PTR2), .ZN(_02697__PTR7) );
  XOR2_X1 U14308 ( .A(P1_P1_InstQueueRd_Addr_PTR3), .B(_02750__PTR2), .Z(_01884__PTR6) );
  XOR2_X1 U14309 ( .A(_02943__PTR4), .B(_02944__PTR3), .Z(_02746__PTR4) );
  XOR2_X1 U14310 ( .A(_02829__PTR1), .B(P1_P1_InstAddrPointer_PTR0), .Z(_02831__PTR1) );
  XOR2_X1 U14311 ( .A(_02084__PTR33), .B(_02084__PTR0), .Z(_02949__PTR1) );
  XOR2_X1 U14312 ( .A(_02941__PTR4), .B(_02942__PTR3), .Z(_02739__PTR4) );
  XOR2_X1 U14313 ( .A(_01932__PTR40), .B(_01836__PTR0), .Z(_02737__PTR0) );
  XOR2_X1 U14314 ( .A(_01932__PTR41), .B(_02735__PTR1), .Z(_02737__PTR1) );
  XOR2_X1 U14315 ( .A(_01932__PTR42), .B(_02735__PTR2), .Z(_02737__PTR2) );
  XOR2_X1 U14316 ( .A(_01932__PTR43), .B(_02735__PTR3), .Z(_02737__PTR3) );
  XOR2_X1 U14317 ( .A(_01932__PTR44), .B(_02735__PTR4), .Z(_02737__PTR4) );
  AND2_X1 U14318 ( .A1(_01932__PTR40), .A2(_01836__PTR0), .ZN(_02738__PTR0) );
  AND2_X1 U14319 ( .A1(_01932__PTR41), .A2(_02735__PTR1), .ZN(_02738__PTR1) );
  AND2_X1 U14320 ( .A1(_01932__PTR42), .A2(_02735__PTR2), .ZN(_02738__PTR2) );
  AND2_X1 U14321 ( .A1(_01932__PTR43), .A2(_02735__PTR3), .ZN(_02738__PTR3) );
  AND2_X1 U14322 ( .A1(_01932__PTR44), .A2(_02735__PTR4), .ZN(_02738__PTR4) );
  XOR2_X1 U14323 ( .A(P1_EBX_PTR1), .B(P1_EBX_PTR0), .Z(_02100__PTR33) );
  XOR2_X1 U14324 ( .A(P1_EBX_PTR2), .B(_02828__PTR1), .Z(_02100__PTR34) );
  XOR2_X1 U14325 ( .A(P1_EBX_PTR3), .B(_02828__PTR2), .Z(_02100__PTR35) );
  XOR2_X1 U14326 ( .A(P1_EBX_PTR4), .B(_02828__PTR3), .Z(_02100__PTR36) );
  XOR2_X1 U14327 ( .A(P1_EBX_PTR5), .B(_02828__PTR4), .Z(_02100__PTR37) );
  XOR2_X1 U14328 ( .A(P1_EBX_PTR6), .B(_02828__PTR5), .Z(_02100__PTR38) );
  XOR2_X1 U14329 ( .A(P1_EBX_PTR7), .B(_02828__PTR6), .Z(_02100__PTR39) );
  XOR2_X1 U14330 ( .A(P1_EBX_PTR8), .B(_02828__PTR7), .Z(_02100__PTR40) );
  XOR2_X1 U14331 ( .A(P1_EBX_PTR9), .B(_02828__PTR8), .Z(_02100__PTR41) );
  XOR2_X1 U14332 ( .A(P1_EBX_PTR10), .B(_02828__PTR9), .Z(_02100__PTR42) );
  XOR2_X1 U14333 ( .A(P1_EBX_PTR11), .B(_02828__PTR10), .Z(_02100__PTR43) );
  XOR2_X1 U14334 ( .A(P1_EBX_PTR12), .B(_02828__PTR11), .Z(_02100__PTR44) );
  XOR2_X1 U14335 ( .A(P1_EBX_PTR13), .B(_02828__PTR12), .Z(_02100__PTR45) );
  XOR2_X1 U14336 ( .A(P1_EBX_PTR14), .B(_02828__PTR13), .Z(_02100__PTR46) );
  XOR2_X1 U14337 ( .A(P1_EBX_PTR15), .B(_02828__PTR14), .Z(_02100__PTR47) );
  XOR2_X1 U14338 ( .A(P1_EBX_PTR16), .B(_02828__PTR15), .Z(_02100__PTR48) );
  XOR2_X1 U14339 ( .A(P1_EBX_PTR17), .B(_02828__PTR16), .Z(_02100__PTR49) );
  XOR2_X1 U14340 ( .A(P1_EBX_PTR18), .B(_02828__PTR17), .Z(_02100__PTR50) );
  XOR2_X1 U14341 ( .A(P1_EBX_PTR19), .B(_02828__PTR18), .Z(_02100__PTR51) );
  XOR2_X1 U14342 ( .A(P1_EBX_PTR20), .B(_02828__PTR19), .Z(_02100__PTR52) );
  XOR2_X1 U14343 ( .A(P1_EBX_PTR21), .B(_02828__PTR20), .Z(_02100__PTR53) );
  XOR2_X1 U14344 ( .A(P1_EBX_PTR22), .B(_02828__PTR21), .Z(_02100__PTR54) );
  XOR2_X1 U14345 ( .A(P1_EBX_PTR23), .B(_02828__PTR22), .Z(_02100__PTR55) );
  XOR2_X1 U14346 ( .A(P1_EBX_PTR24), .B(_02828__PTR23), .Z(_02100__PTR56) );
  XOR2_X1 U14347 ( .A(P1_EBX_PTR25), .B(_02828__PTR24), .Z(_02100__PTR57) );
  XOR2_X1 U14348 ( .A(P1_EBX_PTR26), .B(_02828__PTR25), .Z(_02100__PTR58) );
  XOR2_X1 U14349 ( .A(P1_EBX_PTR27), .B(_02828__PTR26), .Z(_02100__PTR59) );
  XOR2_X1 U14350 ( .A(P1_EBX_PTR28), .B(_02828__PTR27), .Z(_02100__PTR60) );
  XOR2_X1 U14351 ( .A(P1_EBX_PTR29), .B(_02828__PTR28), .Z(_02100__PTR61) );
  XOR2_X1 U14352 ( .A(P1_EBX_PTR30), .B(_02828__PTR29), .Z(_02100__PTR62) );
  XOR2_X1 U14353 ( .A(P1_EBX_PTR31), .B(_02828__PTR30), .Z(_02100__PTR63) );
  XOR2_X1 U14354 ( .A(P1_EAX_PTR1), .B(P1_EAX_PTR0), .Z(_02096__PTR33) );
  XOR2_X1 U14355 ( .A(P1_EAX_PTR2), .B(_02827__PTR1), .Z(_02096__PTR34) );
  XOR2_X1 U14356 ( .A(P1_EAX_PTR3), .B(_02827__PTR2), .Z(_02096__PTR35) );
  XOR2_X1 U14357 ( .A(P1_EAX_PTR4), .B(_02827__PTR3), .Z(_02096__PTR36) );
  XOR2_X1 U14358 ( .A(P1_EAX_PTR5), .B(_02827__PTR4), .Z(_02096__PTR37) );
  XOR2_X1 U14359 ( .A(P1_EAX_PTR6), .B(_02827__PTR5), .Z(_02096__PTR38) );
  XOR2_X1 U14360 ( .A(P1_EAX_PTR7), .B(_02827__PTR6), .Z(_02096__PTR39) );
  XOR2_X1 U14361 ( .A(P1_EAX_PTR8), .B(_02827__PTR7), .Z(_02096__PTR40) );
  XOR2_X1 U14362 ( .A(P1_EAX_PTR9), .B(_02827__PTR8), .Z(_02096__PTR41) );
  XOR2_X1 U14363 ( .A(P1_EAX_PTR10), .B(_02827__PTR9), .Z(_02096__PTR42) );
  XOR2_X1 U14364 ( .A(P1_EAX_PTR11), .B(_02827__PTR10), .Z(_02096__PTR43) );
  XOR2_X1 U14365 ( .A(P1_EAX_PTR12), .B(_02827__PTR11), .Z(_02096__PTR44) );
  XOR2_X1 U14366 ( .A(P1_EAX_PTR13), .B(_02827__PTR12), .Z(_02096__PTR45) );
  XOR2_X1 U14367 ( .A(P1_EAX_PTR14), .B(_02827__PTR13), .Z(_02096__PTR46) );
  XOR2_X1 U14368 ( .A(P1_EAX_PTR15), .B(_02827__PTR14), .Z(_02096__PTR47) );
  XOR2_X1 U14369 ( .A(P1_EAX_PTR16), .B(_02827__PTR15), .Z(_02096__PTR48) );
  XOR2_X1 U14370 ( .A(P1_EAX_PTR17), .B(_02827__PTR16), .Z(_02096__PTR49) );
  XOR2_X1 U14371 ( .A(P1_EAX_PTR18), .B(_02827__PTR17), .Z(_02096__PTR50) );
  XOR2_X1 U14372 ( .A(P1_EAX_PTR19), .B(_02827__PTR18), .Z(_02096__PTR51) );
  XOR2_X1 U14373 ( .A(P1_EAX_PTR20), .B(_02827__PTR19), .Z(_02096__PTR52) );
  XOR2_X1 U14374 ( .A(P1_EAX_PTR21), .B(_02827__PTR20), .Z(_02096__PTR53) );
  XOR2_X1 U14375 ( .A(P1_EAX_PTR22), .B(_02827__PTR21), .Z(_02096__PTR54) );
  XOR2_X1 U14376 ( .A(P1_EAX_PTR23), .B(_02827__PTR22), .Z(_02096__PTR55) );
  XOR2_X1 U14377 ( .A(P1_EAX_PTR24), .B(_02827__PTR23), .Z(_02096__PTR56) );
  XOR2_X1 U14378 ( .A(P1_EAX_PTR25), .B(_02827__PTR24), .Z(_02096__PTR57) );
  XOR2_X1 U14379 ( .A(P1_EAX_PTR26), .B(_02827__PTR25), .Z(_02096__PTR58) );
  XOR2_X1 U14380 ( .A(P1_EAX_PTR27), .B(_02827__PTR26), .Z(_02096__PTR59) );
  XOR2_X1 U14381 ( .A(P1_EAX_PTR28), .B(_02827__PTR27), .Z(_02096__PTR60) );
  XOR2_X1 U14382 ( .A(P1_EAX_PTR29), .B(_02827__PTR28), .Z(_02096__PTR61) );
  XOR2_X1 U14383 ( .A(P1_EAX_PTR30), .B(_02827__PTR29), .Z(_02096__PTR62) );
  XOR2_X1 U14384 ( .A(P1_EAX_PTR31), .B(_02827__PTR30), .Z(_02096__PTR63) );
  XOR2_X1 U14385 ( .A(P1_EAX_PTR17), .B(_02824__PTR0), .Z(_02826__PTR1) );
  XOR2_X1 U14386 ( .A(P1_EAX_PTR18), .B(_02824__PTR1), .Z(_02826__PTR2) );
  XOR2_X1 U14387 ( .A(P1_EAX_PTR19), .B(_02824__PTR2), .Z(_02826__PTR3) );
  XOR2_X1 U14388 ( .A(P1_EAX_PTR20), .B(_02824__PTR3), .Z(_02826__PTR4) );
  XOR2_X1 U14389 ( .A(P1_EAX_PTR21), .B(_02824__PTR4), .Z(_02826__PTR5) );
  XOR2_X1 U14390 ( .A(P1_EAX_PTR22), .B(_02824__PTR5), .Z(_02826__PTR6) );
  XOR2_X1 U14391 ( .A(P1_EAX_PTR23), .B(_02824__PTR6), .Z(_02826__PTR7) );
  XOR2_X1 U14392 ( .A(P1_EAX_PTR24), .B(_02824__PTR7), .Z(_02826__PTR8) );
  XOR2_X1 U14393 ( .A(P1_EAX_PTR25), .B(_02824__PTR8), .Z(_02826__PTR9) );
  XOR2_X1 U14394 ( .A(P1_EAX_PTR26), .B(_02824__PTR9), .Z(_02826__PTR10) );
  XOR2_X1 U14395 ( .A(P1_EAX_PTR27), .B(_02824__PTR10), .Z(_02826__PTR11) );
  XOR2_X1 U14396 ( .A(P1_EAX_PTR28), .B(_02824__PTR11), .Z(_02826__PTR12) );
  XOR2_X1 U14397 ( .A(P1_EAX_PTR29), .B(_02824__PTR12), .Z(_02826__PTR13) );
  XOR2_X1 U14398 ( .A(P1_EAX_PTR30), .B(_02824__PTR13), .Z(_02826__PTR14) );
  XOR2_X1 U14399 ( .A(_02823_), .B(P1_EAX_PTR16), .Z(_02825__PTR0) );
  AND2_X1 U14400 ( .A1(_02823_), .A2(P1_EAX_PTR16), .ZN(_02824__PTR0) );
  XOR2_X1 U14401 ( .A(P1_rEIP_PTR2), .B(P1_rEIP_PTR1), .Z(_02822__PTR1) );
  XOR2_X1 U14402 ( .A(P1_rEIP_PTR3), .B(_02821__PTR1), .Z(_02822__PTR2) );
  XOR2_X1 U14403 ( .A(P1_rEIP_PTR4), .B(_02821__PTR2), .Z(_02822__PTR3) );
  XOR2_X1 U14404 ( .A(P1_rEIP_PTR5), .B(_02821__PTR3), .Z(_02822__PTR4) );
  XOR2_X1 U14405 ( .A(P1_rEIP_PTR6), .B(_02821__PTR4), .Z(_02822__PTR5) );
  XOR2_X1 U14406 ( .A(P1_rEIP_PTR7), .B(_02821__PTR5), .Z(_02822__PTR6) );
  XOR2_X1 U14407 ( .A(P1_rEIP_PTR8), .B(_02821__PTR6), .Z(_02822__PTR7) );
  XOR2_X1 U14408 ( .A(P1_rEIP_PTR9), .B(_02821__PTR7), .Z(_02822__PTR8) );
  XOR2_X1 U14409 ( .A(P1_rEIP_PTR10), .B(_02821__PTR8), .Z(_02822__PTR9) );
  XOR2_X1 U14410 ( .A(P1_rEIP_PTR11), .B(_02821__PTR9), .Z(_02822__PTR10) );
  XOR2_X1 U14411 ( .A(P1_rEIP_PTR12), .B(_02821__PTR10), .Z(_02822__PTR11) );
  XOR2_X1 U14412 ( .A(P1_rEIP_PTR13), .B(_02821__PTR11), .Z(_02822__PTR12) );
  XOR2_X1 U14413 ( .A(P1_rEIP_PTR14), .B(_02821__PTR12), .Z(_02822__PTR13) );
  XOR2_X1 U14414 ( .A(P1_rEIP_PTR15), .B(_02821__PTR13), .Z(_02822__PTR14) );
  XOR2_X1 U14415 ( .A(P1_rEIP_PTR16), .B(_02821__PTR14), .Z(_02822__PTR15) );
  XOR2_X1 U14416 ( .A(P1_rEIP_PTR17), .B(_02821__PTR15), .Z(_02822__PTR16) );
  XOR2_X1 U14417 ( .A(P1_rEIP_PTR18), .B(_02821__PTR16), .Z(_02822__PTR17) );
  XOR2_X1 U14418 ( .A(P1_rEIP_PTR19), .B(_02821__PTR17), .Z(_02822__PTR18) );
  XOR2_X1 U14419 ( .A(P1_rEIP_PTR20), .B(_02821__PTR18), .Z(_02822__PTR19) );
  XOR2_X1 U14420 ( .A(P1_rEIP_PTR21), .B(_02821__PTR19), .Z(_02822__PTR20) );
  XOR2_X1 U14421 ( .A(P1_rEIP_PTR22), .B(_02821__PTR20), .Z(_02822__PTR21) );
  XOR2_X1 U14422 ( .A(P1_rEIP_PTR23), .B(_02821__PTR21), .Z(_02822__PTR22) );
  XOR2_X1 U14423 ( .A(P1_rEIP_PTR24), .B(_02821__PTR22), .Z(_02822__PTR23) );
  XOR2_X1 U14424 ( .A(P1_rEIP_PTR25), .B(_02821__PTR23), .Z(_02822__PTR24) );
  XOR2_X1 U14425 ( .A(P1_rEIP_PTR26), .B(_02821__PTR24), .Z(_02822__PTR25) );
  XOR2_X1 U14426 ( .A(P1_rEIP_PTR27), .B(_02821__PTR25), .Z(_02822__PTR26) );
  XOR2_X1 U14427 ( .A(P1_rEIP_PTR28), .B(_02821__PTR26), .Z(_02822__PTR27) );
  XOR2_X1 U14428 ( .A(P1_rEIP_PTR29), .B(_02821__PTR27), .Z(_02822__PTR28) );
  XOR2_X1 U14429 ( .A(P1_rEIP_PTR30), .B(_02821__PTR28), .Z(_02822__PTR29) );
  XOR2_X1 U14430 ( .A(P1_rEIP_PTR31), .B(_02821__PTR29), .Z(_02822__PTR30) );
  XOR2_X1 U14431 ( .A(_02734__PTR1), .B(_02100__PTR32), .Z(_02948__PTR1) );
  XOR2_X1 U14432 ( .A(_02734__PTR2), .B(_02947__PTR1), .Z(_02948__PTR2) );
  XOR2_X1 U14433 ( .A(_02734__PTR3), .B(_02947__PTR2), .Z(_02948__PTR3) );
  XOR2_X1 U14434 ( .A(_02734__PTR4), .B(_02947__PTR3), .Z(_02948__PTR4) );
  XOR2_X1 U14435 ( .A(_02734__PTR5), .B(_02947__PTR4), .Z(_02948__PTR5) );
  XOR2_X1 U14436 ( .A(_02734__PTR6), .B(_02947__PTR5), .Z(_02948__PTR6) );
  XOR2_X1 U14437 ( .A(_02734__PTR7), .B(_02947__PTR6), .Z(_02948__PTR7) );
  XOR2_X1 U14438 ( .A(_02734__PTR8), .B(_02947__PTR7), .Z(_02948__PTR8) );
  XOR2_X1 U14439 ( .A(_02734__PTR9), .B(_02947__PTR8), .Z(_02948__PTR9) );
  XOR2_X1 U14440 ( .A(_02734__PTR10), .B(_02947__PTR9), .Z(_02948__PTR10) );
  XOR2_X1 U14441 ( .A(_02734__PTR11), .B(_02947__PTR10), .Z(_02948__PTR11) );
  XOR2_X1 U14442 ( .A(_02734__PTR12), .B(_02947__PTR11), .Z(_02948__PTR12) );
  XOR2_X1 U14443 ( .A(_02734__PTR13), .B(_02947__PTR12), .Z(_02948__PTR13) );
  XOR2_X1 U14444 ( .A(_02734__PTR14), .B(_02947__PTR13), .Z(_02948__PTR14) );
  XOR2_X1 U14445 ( .A(_02734__PTR15), .B(_02947__PTR14), .Z(_02948__PTR15) );
  XOR2_X1 U14446 ( .A(_02734__PTR16), .B(_02947__PTR15), .Z(_02948__PTR16) );
  XOR2_X1 U14447 ( .A(_02734__PTR17), .B(_02947__PTR16), .Z(_02948__PTR17) );
  XOR2_X1 U14448 ( .A(_02734__PTR18), .B(_02947__PTR17), .Z(_02948__PTR18) );
  XOR2_X1 U14449 ( .A(_02734__PTR19), .B(_02947__PTR18), .Z(_02948__PTR19) );
  XOR2_X1 U14450 ( .A(_02734__PTR20), .B(_02947__PTR19), .Z(_02948__PTR20) );
  XOR2_X1 U14451 ( .A(_02734__PTR21), .B(_02947__PTR20), .Z(_02948__PTR21) );
  XOR2_X1 U14452 ( .A(_02734__PTR22), .B(_02947__PTR21), .Z(_02948__PTR22) );
  XOR2_X1 U14453 ( .A(_02734__PTR23), .B(_02947__PTR22), .Z(_02948__PTR23) );
  XOR2_X1 U14454 ( .A(_02734__PTR24), .B(_02947__PTR23), .Z(_02948__PTR24) );
  XOR2_X1 U14455 ( .A(_02734__PTR25), .B(_02947__PTR24), .Z(_02948__PTR25) );
  XOR2_X1 U14456 ( .A(_02734__PTR26), .B(_02947__PTR25), .Z(_02948__PTR26) );
  XOR2_X1 U14457 ( .A(_02734__PTR27), .B(_02947__PTR26), .Z(_02948__PTR27) );
  XOR2_X1 U14458 ( .A(_02734__PTR28), .B(_02947__PTR27), .Z(_02948__PTR28) );
  XOR2_X1 U14459 ( .A(_02734__PTR29), .B(_02947__PTR28), .Z(_02948__PTR29) );
  XOR2_X1 U14460 ( .A(_02734__PTR30), .B(_02947__PTR29), .Z(_02948__PTR30) );
  XOR2_X1 U14461 ( .A(_02732__PTR31), .B(_02947__PTR30), .Z(_02948__PTR31) );
  XOR2_X1 U14462 ( .A(_02932__PTR1), .B(_02931__PTR0), .Z(_02717__PTR1) );
  XOR2_X1 U14463 ( .A(_02932__PTR2), .B(_02931__PTR1), .Z(_02717__PTR2) );
  XOR2_X1 U14464 ( .A(_02932__PTR3), .B(_02931__PTR2), .Z(_02717__PTR3) );
  XOR2_X1 U14465 ( .A(_02932__PTR4), .B(_02931__PTR3), .Z(_02717__PTR4) );
  XOR2_X1 U14466 ( .A(P1_P1_InstQueueWr_Addr_PTR0), .B(_01884__PTR3), .Z(_02718__PTR0) );
  XOR2_X1 U14467 ( .A(P1_P1_InstQueueWr_Addr_PTR1), .B(_01890__PTR4), .Z(_02932__PTR1) );
  XOR2_X1 U14468 ( .A(P1_P1_InstQueueWr_Addr_PTR2), .B(_01886__PTR5), .Z(_02932__PTR2) );
  XOR2_X1 U14469 ( .A(P1_P1_InstQueueWr_Addr_PTR3), .B(_02930__PTR3), .Z(_02932__PTR3) );
  XOR2_X1 U14470 ( .A(P1_P1_InstQueueWr_Addr_PTR4), .B(_02751__PTR4), .Z(_02932__PTR4) );
  AND2_X1 U14471 ( .A1(P1_P1_InstQueueWr_Addr_PTR0), .A2(_01884__PTR3), .ZN(_02933__PTR0) );
  AND2_X1 U14472 ( .A1(P1_P1_InstQueueWr_Addr_PTR1), .A2(_01890__PTR4), .ZN(_02933__PTR1) );
  AND2_X1 U14473 ( .A1(P1_P1_InstQueueWr_Addr_PTR2), .A2(_01886__PTR5), .ZN(_02933__PTR2) );
  AND2_X1 U14474 ( .A1(P1_P1_InstQueueWr_Addr_PTR3), .A2(_02930__PTR3), .ZN(_02933__PTR3) );
  AND2_X1 U14475 ( .A1(P1_P1_InstQueueWr_Addr_PTR4), .A2(_02751__PTR4), .ZN(_02933__PTR4) );
  XOR2_X1 U14476 ( .A(_01886__PTR5), .B(_02750__PTR1), .Z(_02820__PTR2) );
  XOR2_X1 U14477 ( .A(P1_P1_InstQueueRd_Addr_PTR3), .B(_02819__PTR2), .Z(_02820__PTR3) );
  XOR2_X1 U14478 ( .A(P1_P1_InstQueueRd_Addr_PTR2), .B(P1_P1_InstQueueRd_Addr_PTR1), .Z(_01890__PTR5) );
  XOR2_X1 U14479 ( .A(P1_P1_InstQueueRd_Addr_PTR3), .B(_02817__PTR1), .Z(_01890__PTR6) );
  XOR2_X1 U14480 ( .A(P1_P1_InstQueueRd_Addr_PTR4), .B(_02817__PTR2), .Z(_02818__PTR3) );
  XOR2_X1 U14481 ( .A(_01887__PTR1), .B(_02814__PTR0), .Z(_02816__PTR1) );
  XOR2_X1 U14482 ( .A(_01887__PTR2), .B(_02814__PTR1), .Z(_02816__PTR2) );
  XOR2_X1 U14483 ( .A(_01887__PTR3), .B(_02814__PTR2), .Z(_02816__PTR3) );
  XOR2_X1 U14484 ( .A(_01887__PTR4), .B(_02814__PTR3), .Z(_02816__PTR4) );
  XOR2_X1 U14485 ( .A(_01887__PTR5), .B(_02814__PTR4), .Z(_02816__PTR5) );
  XOR2_X1 U14486 ( .A(_01887__PTR6), .B(_02814__PTR5), .Z(_02816__PTR6) );
  XOR2_X1 U14487 ( .A(_01887__PTR7), .B(_02814__PTR6), .Z(_02816__PTR7) );
  XOR2_X1 U14488 ( .A(_01887__PTR0), .B(_01889__PTR7), .Z(_02815__PTR0) );
  AND2_X1 U14489 ( .A1(_01887__PTR0), .A2(_01889__PTR7), .ZN(_02814__PTR0) );
  XOR2_X1 U14490 ( .A(_01890__PTR4), .B(P1_P1_InstQueueRd_Addr_PTR0), .Z(_01888__PTR4) );
  XOR2_X1 U14491 ( .A(P1_P1_InstQueueRd_Addr_PTR2), .B(_02813__PTR1), .Z(_01888__PTR5) );
  XOR2_X1 U14492 ( .A(P1_P1_InstQueueRd_Addr_PTR3), .B(_02813__PTR2), .Z(_01888__PTR6) );
  XOR2_X1 U14493 ( .A(P1_P1_InstQueueRd_Addr_PTR3), .B(P1_P1_InstQueueRd_Addr_PTR2), .Z(_01886__PTR6) );
  XOR2_X1 U14494 ( .A(_02745__PTR2), .B(_02798__PTR1), .Z(_02807__PTR2) );
  XOR2_X1 U14495 ( .A(P1_P1_InstAddrPointer_PTR3), .B(_02806__PTR2), .Z(_02807__PTR3) );
  XOR2_X1 U14496 ( .A(P1_P1_InstAddrPointer_PTR4), .B(_02806__PTR3), .Z(_02807__PTR4) );
  XOR2_X1 U14497 ( .A(P1_P1_InstAddrPointer_PTR5), .B(_02806__PTR4), .Z(_02807__PTR5) );
  XOR2_X1 U14498 ( .A(P1_P1_InstAddrPointer_PTR6), .B(_02806__PTR5), .Z(_02807__PTR6) );
  XOR2_X1 U14499 ( .A(P1_P1_InstAddrPointer_PTR7), .B(_02806__PTR6), .Z(_02807__PTR7) );
  XOR2_X1 U14500 ( .A(P1_P1_InstAddrPointer_PTR8), .B(_02806__PTR7), .Z(_02807__PTR8) );
  XOR2_X1 U14501 ( .A(P1_P1_InstAddrPointer_PTR9), .B(_02806__PTR8), .Z(_02807__PTR9) );
  XOR2_X1 U14502 ( .A(P1_P1_InstAddrPointer_PTR10), .B(_02806__PTR9), .Z(_02807__PTR10) );
  XOR2_X1 U14503 ( .A(P1_P1_InstAddrPointer_PTR11), .B(_02806__PTR10), .Z(_02807__PTR11) );
  XOR2_X1 U14504 ( .A(P1_P1_InstAddrPointer_PTR12), .B(_02806__PTR11), .Z(_02807__PTR12) );
  XOR2_X1 U14505 ( .A(P1_P1_InstAddrPointer_PTR13), .B(_02806__PTR12), .Z(_02807__PTR13) );
  XOR2_X1 U14506 ( .A(P1_P1_InstAddrPointer_PTR14), .B(_02806__PTR13), .Z(_02807__PTR14) );
  XOR2_X1 U14507 ( .A(P1_P1_InstAddrPointer_PTR15), .B(_02806__PTR14), .Z(_02807__PTR15) );
  XOR2_X1 U14508 ( .A(P1_P1_InstAddrPointer_PTR16), .B(_02806__PTR15), .Z(_02807__PTR16) );
  XOR2_X1 U14509 ( .A(P1_P1_InstAddrPointer_PTR17), .B(_02806__PTR16), .Z(_02807__PTR17) );
  XOR2_X1 U14510 ( .A(P1_P1_InstAddrPointer_PTR18), .B(_02806__PTR17), .Z(_02807__PTR18) );
  XOR2_X1 U14511 ( .A(P1_P1_InstAddrPointer_PTR19), .B(_02806__PTR18), .Z(_02807__PTR19) );
  XOR2_X1 U14512 ( .A(P1_P1_InstAddrPointer_PTR20), .B(_02806__PTR19), .Z(_02807__PTR20) );
  XOR2_X1 U14513 ( .A(P1_P1_InstAddrPointer_PTR21), .B(_02806__PTR20), .Z(_02807__PTR21) );
  XOR2_X1 U14514 ( .A(P1_P1_InstAddrPointer_PTR22), .B(_02806__PTR21), .Z(_02807__PTR22) );
  XOR2_X1 U14515 ( .A(P1_P1_InstAddrPointer_PTR23), .B(_02806__PTR22), .Z(_02807__PTR23) );
  XOR2_X1 U14516 ( .A(P1_P1_InstAddrPointer_PTR24), .B(_02806__PTR23), .Z(_02807__PTR24) );
  XOR2_X1 U14517 ( .A(P1_P1_InstAddrPointer_PTR25), .B(_02806__PTR24), .Z(_02807__PTR25) );
  XOR2_X1 U14518 ( .A(P1_P1_InstAddrPointer_PTR26), .B(_02806__PTR25), .Z(_02807__PTR26) );
  XOR2_X1 U14519 ( .A(P1_P1_InstAddrPointer_PTR27), .B(_02806__PTR26), .Z(_02807__PTR27) );
  XOR2_X1 U14520 ( .A(P1_P1_InstAddrPointer_PTR28), .B(_02806__PTR27), .Z(_02807__PTR28) );
  XOR2_X1 U14521 ( .A(P1_P1_InstAddrPointer_PTR29), .B(_02806__PTR28), .Z(_02807__PTR29) );
  XOR2_X1 U14522 ( .A(P1_P1_InstAddrPointer_PTR30), .B(_02806__PTR29), .Z(_02807__PTR30) );
  XOR2_X1 U14523 ( .A(P1_P1_InstAddrPointer_PTR31), .B(_02806__PTR30), .Z(_02807__PTR31) );
  XOR2_X1 U14524 ( .A(_02809__PTR1), .B(_02808__PTR0), .Z(_02810__PTR1) );
  XOR2_X1 U14525 ( .A(_02809__PTR2), .B(_02808__PTR1), .Z(_02810__PTR2) );
  XOR2_X1 U14526 ( .A(_02809__PTR3), .B(_02808__PTR2), .Z(_02810__PTR3) );
  XOR2_X1 U14527 ( .A(_02809__PTR4), .B(_02808__PTR3), .Z(_02810__PTR4) );
  XOR2_X1 U14528 ( .A(_02809__PTR5), .B(_02808__PTR4), .Z(_02810__PTR5) );
  XOR2_X1 U14529 ( .A(_02809__PTR6), .B(_02808__PTR5), .Z(_02810__PTR6) );
  XOR2_X1 U14530 ( .A(_02809__PTR7), .B(_02808__PTR6), .Z(_02810__PTR7) );
  XOR2_X1 U14531 ( .A(_02807__PTR8), .B(_02808__PTR7), .Z(_02810__PTR8) );
  XOR2_X1 U14532 ( .A(_02807__PTR9), .B(_02808__PTR8), .Z(_02810__PTR9) );
  XOR2_X1 U14533 ( .A(_02807__PTR10), .B(_02808__PTR9), .Z(_02810__PTR10) );
  XOR2_X1 U14534 ( .A(_02807__PTR11), .B(_02808__PTR10), .Z(_02810__PTR11) );
  XOR2_X1 U14535 ( .A(_02807__PTR12), .B(_02808__PTR11), .Z(_02810__PTR12) );
  XOR2_X1 U14536 ( .A(_02807__PTR13), .B(_02808__PTR12), .Z(_02810__PTR13) );
  XOR2_X1 U14537 ( .A(_02807__PTR14), .B(_02808__PTR13), .Z(_02810__PTR14) );
  XOR2_X1 U14538 ( .A(_02807__PTR15), .B(_02808__PTR14), .Z(_02810__PTR15) );
  XOR2_X1 U14539 ( .A(_02807__PTR16), .B(_02808__PTR15), .Z(_02810__PTR16) );
  XOR2_X1 U14540 ( .A(_02807__PTR17), .B(_02808__PTR16), .Z(_02810__PTR17) );
  XOR2_X1 U14541 ( .A(_02807__PTR18), .B(_02808__PTR17), .Z(_02810__PTR18) );
  XOR2_X1 U14542 ( .A(_02807__PTR19), .B(_02808__PTR18), .Z(_02810__PTR19) );
  XOR2_X1 U14543 ( .A(_02807__PTR20), .B(_02808__PTR19), .Z(_02810__PTR20) );
  XOR2_X1 U14544 ( .A(_02807__PTR21), .B(_02808__PTR20), .Z(_02810__PTR21) );
  XOR2_X1 U14545 ( .A(_02807__PTR22), .B(_02808__PTR21), .Z(_02810__PTR22) );
  XOR2_X1 U14546 ( .A(_02807__PTR23), .B(_02808__PTR22), .Z(_02810__PTR23) );
  XOR2_X1 U14547 ( .A(_02807__PTR24), .B(_02808__PTR23), .Z(_02810__PTR24) );
  XOR2_X1 U14548 ( .A(_02807__PTR25), .B(_02808__PTR24), .Z(_02810__PTR25) );
  XOR2_X1 U14549 ( .A(_02807__PTR26), .B(_02808__PTR25), .Z(_02810__PTR26) );
  XOR2_X1 U14550 ( .A(_02807__PTR27), .B(_02808__PTR26), .Z(_02810__PTR27) );
  XOR2_X1 U14551 ( .A(_02807__PTR28), .B(_02808__PTR27), .Z(_02810__PTR28) );
  XOR2_X1 U14552 ( .A(_02807__PTR29), .B(_02808__PTR28), .Z(_02810__PTR29) );
  XOR2_X1 U14553 ( .A(_02807__PTR30), .B(_02808__PTR29), .Z(_02810__PTR30) );
  XOR2_X1 U14554 ( .A(_02807__PTR31), .B(_02808__PTR30), .Z(_02810__PTR31) );
  XOR2_X1 U14555 ( .A(_02084__PTR0), .B(_01885__PTR0), .Z(_02809__PTR0) );
  XOR2_X1 U14556 ( .A(_02084__PTR1), .B(_01885__PTR1), .Z(_02809__PTR1) );
  XOR2_X1 U14557 ( .A(_02807__PTR2), .B(_01885__PTR2), .Z(_02809__PTR2) );
  XOR2_X1 U14558 ( .A(_02807__PTR3), .B(_01885__PTR3), .Z(_02809__PTR3) );
  XOR2_X1 U14559 ( .A(_02807__PTR4), .B(_01885__PTR4), .Z(_02809__PTR4) );
  XOR2_X1 U14560 ( .A(_02807__PTR5), .B(_01885__PTR5), .Z(_02809__PTR5) );
  XOR2_X1 U14561 ( .A(_02807__PTR6), .B(_01885__PTR6), .Z(_02809__PTR6) );
  XOR2_X1 U14562 ( .A(_02807__PTR7), .B(_01885__PTR7), .Z(_02809__PTR7) );
  AND2_X1 U14563 ( .A1(_02084__PTR0), .A2(_01885__PTR0), .ZN(_02808__PTR0) );
  AND2_X1 U14564 ( .A1(_02084__PTR1), .A2(_01885__PTR1), .ZN(_02811__PTR1) );
  AND2_X1 U14565 ( .A1(_02807__PTR2), .A2(_01885__PTR2), .ZN(_02811__PTR2) );
  AND2_X1 U14566 ( .A1(_02807__PTR3), .A2(_01885__PTR3), .ZN(_02811__PTR3) );
  AND2_X1 U14567 ( .A1(_02807__PTR4), .A2(_01885__PTR4), .ZN(_02811__PTR4) );
  AND2_X1 U14568 ( .A1(_02807__PTR5), .A2(_01885__PTR5), .ZN(_02811__PTR5) );
  AND2_X1 U14569 ( .A1(_02807__PTR6), .A2(_01885__PTR6), .ZN(_02811__PTR6) );
  AND2_X1 U14570 ( .A1(_02807__PTR7), .A2(_01885__PTR7), .ZN(_02811__PTR7) );
  XOR2_X1 U14571 ( .A(P1_P1_InstAddrPointer_PTR2), .B(P1_P1_InstAddrPointer_PTR1), .Z(_02084__PTR34) );
  XOR2_X1 U14572 ( .A(P1_P1_InstAddrPointer_PTR3), .B(_02801__PTR1), .Z(_02084__PTR35) );
  XOR2_X1 U14573 ( .A(P1_P1_InstAddrPointer_PTR4), .B(_02801__PTR2), .Z(_02084__PTR36) );
  XOR2_X1 U14574 ( .A(P1_P1_InstAddrPointer_PTR5), .B(_02801__PTR3), .Z(_02084__PTR37) );
  XOR2_X1 U14575 ( .A(P1_P1_InstAddrPointer_PTR6), .B(_02801__PTR4), .Z(_02084__PTR38) );
  XOR2_X1 U14576 ( .A(P1_P1_InstAddrPointer_PTR7), .B(_02801__PTR5), .Z(_02084__PTR39) );
  XOR2_X1 U14577 ( .A(P1_P1_InstAddrPointer_PTR8), .B(_02801__PTR6), .Z(_02084__PTR40) );
  XOR2_X1 U14578 ( .A(P1_P1_InstAddrPointer_PTR9), .B(_02801__PTR7), .Z(_02084__PTR41) );
  XOR2_X1 U14579 ( .A(P1_P1_InstAddrPointer_PTR10), .B(_02801__PTR8), .Z(_02084__PTR42) );
  XOR2_X1 U14580 ( .A(P1_P1_InstAddrPointer_PTR11), .B(_02801__PTR9), .Z(_02084__PTR43) );
  XOR2_X1 U14581 ( .A(P1_P1_InstAddrPointer_PTR12), .B(_02801__PTR10), .Z(_02084__PTR44) );
  XOR2_X1 U14582 ( .A(P1_P1_InstAddrPointer_PTR13), .B(_02801__PTR11), .Z(_02084__PTR45) );
  XOR2_X1 U14583 ( .A(P1_P1_InstAddrPointer_PTR14), .B(_02801__PTR12), .Z(_02084__PTR46) );
  XOR2_X1 U14584 ( .A(P1_P1_InstAddrPointer_PTR15), .B(_02801__PTR13), .Z(_02084__PTR47) );
  XOR2_X1 U14585 ( .A(P1_P1_InstAddrPointer_PTR16), .B(_02801__PTR14), .Z(_02084__PTR48) );
  XOR2_X1 U14586 ( .A(P1_P1_InstAddrPointer_PTR17), .B(_02801__PTR15), .Z(_02084__PTR49) );
  XOR2_X1 U14587 ( .A(P1_P1_InstAddrPointer_PTR18), .B(_02801__PTR16), .Z(_02084__PTR50) );
  XOR2_X1 U14588 ( .A(P1_P1_InstAddrPointer_PTR19), .B(_02801__PTR17), .Z(_02084__PTR51) );
  XOR2_X1 U14589 ( .A(P1_P1_InstAddrPointer_PTR20), .B(_02801__PTR18), .Z(_02084__PTR52) );
  XOR2_X1 U14590 ( .A(P1_P1_InstAddrPointer_PTR21), .B(_02801__PTR19), .Z(_02084__PTR53) );
  XOR2_X1 U14591 ( .A(P1_P1_InstAddrPointer_PTR22), .B(_02801__PTR20), .Z(_02084__PTR54) );
  XOR2_X1 U14592 ( .A(P1_P1_InstAddrPointer_PTR23), .B(_02801__PTR21), .Z(_02084__PTR55) );
  XOR2_X1 U14593 ( .A(P1_P1_InstAddrPointer_PTR24), .B(_02801__PTR22), .Z(_02084__PTR56) );
  XOR2_X1 U14594 ( .A(P1_P1_InstAddrPointer_PTR25), .B(_02801__PTR23), .Z(_02084__PTR57) );
  XOR2_X1 U14595 ( .A(P1_P1_InstAddrPointer_PTR26), .B(_02801__PTR24), .Z(_02084__PTR58) );
  XOR2_X1 U14596 ( .A(P1_P1_InstAddrPointer_PTR27), .B(_02801__PTR25), .Z(_02084__PTR59) );
  XOR2_X1 U14597 ( .A(P1_P1_InstAddrPointer_PTR28), .B(_02801__PTR26), .Z(_02084__PTR60) );
  XOR2_X1 U14598 ( .A(P1_P1_InstAddrPointer_PTR29), .B(_02801__PTR27), .Z(_02084__PTR61) );
  XOR2_X1 U14599 ( .A(P1_P1_InstAddrPointer_PTR30), .B(_02801__PTR28), .Z(_02084__PTR62) );
  XOR2_X1 U14600 ( .A(P1_P1_InstAddrPointer_PTR31), .B(_02801__PTR29), .Z(_02084__PTR63) );
  XOR2_X1 U14601 ( .A(_02803__PTR1), .B(_02802__PTR0), .Z(_02804__PTR1) );
  XOR2_X1 U14602 ( .A(_02803__PTR2), .B(_02802__PTR1), .Z(_02804__PTR2) );
  XOR2_X1 U14603 ( .A(_02803__PTR3), .B(_02802__PTR2), .Z(_02804__PTR3) );
  XOR2_X1 U14604 ( .A(_02803__PTR4), .B(_02802__PTR3), .Z(_02804__PTR4) );
  XOR2_X1 U14605 ( .A(_02803__PTR5), .B(_02802__PTR4), .Z(_02804__PTR5) );
  XOR2_X1 U14606 ( .A(_02803__PTR6), .B(_02802__PTR5), .Z(_02804__PTR6) );
  XOR2_X1 U14607 ( .A(_02803__PTR7), .B(_02802__PTR6), .Z(_02804__PTR7) );
  XOR2_X1 U14608 ( .A(_02084__PTR40), .B(_02802__PTR7), .Z(_02804__PTR8) );
  XOR2_X1 U14609 ( .A(_02084__PTR41), .B(_02802__PTR8), .Z(_02804__PTR9) );
  XOR2_X1 U14610 ( .A(_02084__PTR42), .B(_02802__PTR9), .Z(_02804__PTR10) );
  XOR2_X1 U14611 ( .A(_02084__PTR43), .B(_02802__PTR10), .Z(_02804__PTR11) );
  XOR2_X1 U14612 ( .A(_02084__PTR44), .B(_02802__PTR11), .Z(_02804__PTR12) );
  XOR2_X1 U14613 ( .A(_02084__PTR45), .B(_02802__PTR12), .Z(_02804__PTR13) );
  XOR2_X1 U14614 ( .A(_02084__PTR46), .B(_02802__PTR13), .Z(_02804__PTR14) );
  XOR2_X1 U14615 ( .A(_02084__PTR47), .B(_02802__PTR14), .Z(_02804__PTR15) );
  XOR2_X1 U14616 ( .A(_02084__PTR48), .B(_02802__PTR15), .Z(_02804__PTR16) );
  XOR2_X1 U14617 ( .A(_02084__PTR49), .B(_02802__PTR16), .Z(_02804__PTR17) );
  XOR2_X1 U14618 ( .A(_02084__PTR50), .B(_02802__PTR17), .Z(_02804__PTR18) );
  XOR2_X1 U14619 ( .A(_02084__PTR51), .B(_02802__PTR18), .Z(_02804__PTR19) );
  XOR2_X1 U14620 ( .A(_02084__PTR52), .B(_02802__PTR19), .Z(_02804__PTR20) );
  XOR2_X1 U14621 ( .A(_02084__PTR53), .B(_02802__PTR20), .Z(_02804__PTR21) );
  XOR2_X1 U14622 ( .A(_02084__PTR54), .B(_02802__PTR21), .Z(_02804__PTR22) );
  XOR2_X1 U14623 ( .A(_02084__PTR55), .B(_02802__PTR22), .Z(_02804__PTR23) );
  XOR2_X1 U14624 ( .A(_02084__PTR56), .B(_02802__PTR23), .Z(_02804__PTR24) );
  XOR2_X1 U14625 ( .A(_02084__PTR57), .B(_02802__PTR24), .Z(_02804__PTR25) );
  XOR2_X1 U14626 ( .A(_02084__PTR58), .B(_02802__PTR25), .Z(_02804__PTR26) );
  XOR2_X1 U14627 ( .A(_02084__PTR59), .B(_02802__PTR26), .Z(_02804__PTR27) );
  XOR2_X1 U14628 ( .A(_02084__PTR60), .B(_02802__PTR27), .Z(_02804__PTR28) );
  XOR2_X1 U14629 ( .A(_02084__PTR61), .B(_02802__PTR28), .Z(_02804__PTR29) );
  XOR2_X1 U14630 ( .A(_02084__PTR62), .B(_02802__PTR29), .Z(_02804__PTR30) );
  XOR2_X1 U14631 ( .A(_02084__PTR63), .B(_02802__PTR30), .Z(_02804__PTR31) );
  XOR2_X1 U14632 ( .A(P1_P1_InstAddrPointer_PTR0), .B(_01885__PTR0), .Z(_02803__PTR0) );
  XOR2_X1 U14633 ( .A(_02084__PTR33), .B(_01885__PTR1), .Z(_02803__PTR1) );
  XOR2_X1 U14634 ( .A(_02084__PTR34), .B(_01885__PTR2), .Z(_02803__PTR2) );
  XOR2_X1 U14635 ( .A(_02084__PTR35), .B(_01885__PTR3), .Z(_02803__PTR3) );
  XOR2_X1 U14636 ( .A(_02084__PTR36), .B(_01885__PTR4), .Z(_02803__PTR4) );
  XOR2_X1 U14637 ( .A(_02084__PTR37), .B(_01885__PTR5), .Z(_02803__PTR5) );
  XOR2_X1 U14638 ( .A(_02084__PTR38), .B(_01885__PTR6), .Z(_02803__PTR6) );
  XOR2_X1 U14639 ( .A(_02084__PTR39), .B(_01885__PTR7), .Z(_02803__PTR7) );
  AND2_X1 U14640 ( .A1(P1_P1_InstAddrPointer_PTR0), .A2(_01885__PTR0), .ZN(_02802__PTR0) );
  AND2_X1 U14641 ( .A1(_02084__PTR33), .A2(_01885__PTR1), .ZN(_02805__PTR1) );
  AND2_X1 U14642 ( .A1(_02084__PTR34), .A2(_01885__PTR2), .ZN(_02805__PTR2) );
  AND2_X1 U14643 ( .A1(_02084__PTR35), .A2(_01885__PTR3), .ZN(_02805__PTR3) );
  AND2_X1 U14644 ( .A1(_02084__PTR36), .A2(_01885__PTR4), .ZN(_02805__PTR4) );
  AND2_X1 U14645 ( .A1(_02084__PTR37), .A2(_01885__PTR5), .ZN(_02805__PTR5) );
  AND2_X1 U14646 ( .A1(_02084__PTR38), .A2(_01885__PTR6), .ZN(_02805__PTR6) );
  AND2_X1 U14647 ( .A1(_02084__PTR39), .A2(_01885__PTR7), .ZN(_02805__PTR7) );
  XOR2_X1 U14648 ( .A(_01885__PTR7), .B(_02724__PTR6), .Z(_02935__PTR7) );
  XOR2_X1 U14649 ( .A(P1_P1_InstAddrPointer_PTR1), .B(P1_P1_InstAddrPointer_PTR0), .Z(_02084__PTR1) );
  XOR2_X1 U14650 ( .A(P1_P1_InstAddrPointer_PTR2), .B(_02798__PTR1), .Z(_02084__PTR2) );
  XOR2_X1 U14651 ( .A(P1_P1_InstAddrPointer_PTR3), .B(_02798__PTR2), .Z(_02084__PTR3) );
  XOR2_X1 U14652 ( .A(P1_P1_InstAddrPointer_PTR4), .B(_02798__PTR3), .Z(_02084__PTR4) );
  XOR2_X1 U14653 ( .A(P1_P1_InstAddrPointer_PTR5), .B(_02798__PTR4), .Z(_02084__PTR5) );
  XOR2_X1 U14654 ( .A(P1_P1_InstAddrPointer_PTR6), .B(_02798__PTR5), .Z(_02084__PTR6) );
  XOR2_X1 U14655 ( .A(P1_P1_InstAddrPointer_PTR7), .B(_02798__PTR6), .Z(_02084__PTR7) );
  XOR2_X1 U14656 ( .A(P1_P1_InstAddrPointer_PTR8), .B(_02798__PTR7), .Z(_02084__PTR8) );
  XOR2_X1 U14657 ( .A(P1_P1_InstAddrPointer_PTR9), .B(_02798__PTR8), .Z(_02084__PTR9) );
  XOR2_X1 U14658 ( .A(P1_P1_InstAddrPointer_PTR10), .B(_02798__PTR9), .Z(_02084__PTR10) );
  XOR2_X1 U14659 ( .A(P1_P1_InstAddrPointer_PTR11), .B(_02798__PTR10), .Z(_02084__PTR11) );
  XOR2_X1 U14660 ( .A(P1_P1_InstAddrPointer_PTR12), .B(_02798__PTR11), .Z(_02084__PTR12) );
  XOR2_X1 U14661 ( .A(P1_P1_InstAddrPointer_PTR13), .B(_02798__PTR12), .Z(_02084__PTR13) );
  XOR2_X1 U14662 ( .A(P1_P1_InstAddrPointer_PTR14), .B(_02798__PTR13), .Z(_02084__PTR14) );
  XOR2_X1 U14663 ( .A(P1_P1_InstAddrPointer_PTR15), .B(_02798__PTR14), .Z(_02084__PTR15) );
  XOR2_X1 U14664 ( .A(P1_P1_InstAddrPointer_PTR16), .B(_02798__PTR15), .Z(_02084__PTR16) );
  XOR2_X1 U14665 ( .A(P1_P1_InstAddrPointer_PTR17), .B(_02798__PTR16), .Z(_02084__PTR17) );
  XOR2_X1 U14666 ( .A(P1_P1_InstAddrPointer_PTR18), .B(_02798__PTR17), .Z(_02084__PTR18) );
  XOR2_X1 U14667 ( .A(P1_P1_InstAddrPointer_PTR19), .B(_02798__PTR18), .Z(_02084__PTR19) );
  XOR2_X1 U14668 ( .A(P1_P1_InstAddrPointer_PTR20), .B(_02798__PTR19), .Z(_02084__PTR20) );
  XOR2_X1 U14669 ( .A(P1_P1_InstAddrPointer_PTR21), .B(_02798__PTR20), .Z(_02084__PTR21) );
  XOR2_X1 U14670 ( .A(P1_P1_InstAddrPointer_PTR22), .B(_02798__PTR21), .Z(_02084__PTR22) );
  XOR2_X1 U14671 ( .A(P1_P1_InstAddrPointer_PTR23), .B(_02798__PTR22), .Z(_02084__PTR23) );
  XOR2_X1 U14672 ( .A(P1_P1_InstAddrPointer_PTR24), .B(_02798__PTR23), .Z(_02084__PTR24) );
  XOR2_X1 U14673 ( .A(P1_P1_InstAddrPointer_PTR25), .B(_02798__PTR24), .Z(_02084__PTR25) );
  XOR2_X1 U14674 ( .A(P1_P1_InstAddrPointer_PTR26), .B(_02798__PTR25), .Z(_02084__PTR26) );
  XOR2_X1 U14675 ( .A(P1_P1_InstAddrPointer_PTR27), .B(_02798__PTR26), .Z(_02084__PTR27) );
  XOR2_X1 U14676 ( .A(P1_P1_InstAddrPointer_PTR28), .B(_02798__PTR27), .Z(_02084__PTR28) );
  XOR2_X1 U14677 ( .A(P1_P1_InstAddrPointer_PTR29), .B(_02798__PTR28), .Z(_02084__PTR29) );
  XOR2_X1 U14678 ( .A(P1_P1_InstAddrPointer_PTR30), .B(_02798__PTR29), .Z(_02084__PTR30) );
  XOR2_X1 U14679 ( .A(P1_P1_InstAddrPointer_PTR31), .B(_02798__PTR30), .Z(_02084__PTR31) );
  XOR2_X1 U14680 ( .A(_02809__PTR1), .B(_02937__PTR0), .Z(_02939__PTR1) );
  XOR2_X1 U14681 ( .A(_02938__PTR2), .B(_02937__PTR1), .Z(_02939__PTR2) );
  XOR2_X1 U14682 ( .A(_02938__PTR3), .B(_02937__PTR2), .Z(_02939__PTR3) );
  XOR2_X1 U14683 ( .A(_02938__PTR4), .B(_02937__PTR3), .Z(_02939__PTR4) );
  XOR2_X1 U14684 ( .A(_02938__PTR5), .B(_02937__PTR4), .Z(_02939__PTR5) );
  XOR2_X1 U14685 ( .A(_02938__PTR6), .B(_02937__PTR5), .Z(_02939__PTR6) );
  XOR2_X1 U14686 ( .A(_02938__PTR7), .B(_02937__PTR6), .Z(_02939__PTR7) );
  XOR2_X1 U14687 ( .A(_02938__PTR8), .B(_02937__PTR7), .Z(_02939__PTR8) );
  XOR2_X1 U14688 ( .A(_02938__PTR9), .B(_02937__PTR8), .Z(_02939__PTR9) );
  XOR2_X1 U14689 ( .A(_02938__PTR10), .B(_02937__PTR9), .Z(_02939__PTR10) );
  XOR2_X1 U14690 ( .A(_02938__PTR11), .B(_02937__PTR10), .Z(_02939__PTR11) );
  XOR2_X1 U14691 ( .A(_02938__PTR12), .B(_02937__PTR11), .Z(_02939__PTR12) );
  XOR2_X1 U14692 ( .A(_02938__PTR13), .B(_02937__PTR12), .Z(_02939__PTR13) );
  XOR2_X1 U14693 ( .A(_02938__PTR14), .B(_02937__PTR13), .Z(_02939__PTR14) );
  XOR2_X1 U14694 ( .A(_02938__PTR15), .B(_02937__PTR14), .Z(_02939__PTR15) );
  XOR2_X1 U14695 ( .A(_02938__PTR16), .B(_02937__PTR15), .Z(_02939__PTR16) );
  XOR2_X1 U14696 ( .A(_02938__PTR17), .B(_02937__PTR16), .Z(_02939__PTR17) );
  XOR2_X1 U14697 ( .A(_02938__PTR18), .B(_02937__PTR17), .Z(_02939__PTR18) );
  XOR2_X1 U14698 ( .A(_02938__PTR19), .B(_02937__PTR18), .Z(_02939__PTR19) );
  XOR2_X1 U14699 ( .A(_02938__PTR20), .B(_02937__PTR19), .Z(_02939__PTR20) );
  XOR2_X1 U14700 ( .A(_02938__PTR21), .B(_02937__PTR20), .Z(_02939__PTR21) );
  XOR2_X1 U14701 ( .A(_02938__PTR22), .B(_02937__PTR21), .Z(_02939__PTR22) );
  XOR2_X1 U14702 ( .A(_02938__PTR23), .B(_02937__PTR22), .Z(_02939__PTR23) );
  XOR2_X1 U14703 ( .A(_02938__PTR24), .B(_02937__PTR23), .Z(_02939__PTR24) );
  XOR2_X1 U14704 ( .A(_02938__PTR25), .B(_02937__PTR24), .Z(_02939__PTR25) );
  XOR2_X1 U14705 ( .A(_02938__PTR26), .B(_02937__PTR25), .Z(_02939__PTR26) );
  XOR2_X1 U14706 ( .A(_02938__PTR27), .B(_02937__PTR26), .Z(_02939__PTR27) );
  XOR2_X1 U14707 ( .A(_02938__PTR28), .B(_02937__PTR27), .Z(_02939__PTR28) );
  XOR2_X1 U14708 ( .A(_02938__PTR29), .B(_02937__PTR28), .Z(_02939__PTR29) );
  XOR2_X1 U14709 ( .A(_02938__PTR30), .B(_02937__PTR29), .Z(_02939__PTR30) );
  XOR2_X1 U14710 ( .A(_02938__PTR32), .B(_02937__PTR30), .Z(_02939__PTR31) );
  XOR2_X1 U14711 ( .A(_02084__PTR2), .B(_01885__PTR2), .Z(_02938__PTR2) );
  XOR2_X1 U14712 ( .A(_02084__PTR3), .B(_01885__PTR3), .Z(_02938__PTR3) );
  XOR2_X1 U14713 ( .A(_02084__PTR4), .B(_02936__PTR4), .Z(_02938__PTR4) );
  XOR2_X1 U14714 ( .A(_02084__PTR5), .B(_02936__PTR5), .Z(_02938__PTR5) );
  XOR2_X1 U14715 ( .A(_02084__PTR6), .B(_02936__PTR6), .Z(_02938__PTR6) );
  XOR2_X1 U14716 ( .A(_02084__PTR7), .B(_02936__PTR7), .Z(_02938__PTR7) );
  XOR2_X1 U14717 ( .A(_02084__PTR8), .B(_02934__PTR8), .Z(_02938__PTR8) );
  XOR2_X1 U14718 ( .A(_02084__PTR9), .B(_02934__PTR8), .Z(_02938__PTR9) );
  XOR2_X1 U14719 ( .A(_02084__PTR10), .B(_02934__PTR8), .Z(_02938__PTR10) );
  XOR2_X1 U14720 ( .A(_02084__PTR11), .B(_02934__PTR8), .Z(_02938__PTR11) );
  XOR2_X1 U14721 ( .A(_02084__PTR12), .B(_02934__PTR8), .Z(_02938__PTR12) );
  XOR2_X1 U14722 ( .A(_02084__PTR13), .B(_02934__PTR8), .Z(_02938__PTR13) );
  XOR2_X1 U14723 ( .A(_02084__PTR14), .B(_02934__PTR8), .Z(_02938__PTR14) );
  XOR2_X1 U14724 ( .A(_02084__PTR15), .B(_02934__PTR8), .Z(_02938__PTR15) );
  XOR2_X1 U14725 ( .A(_02084__PTR16), .B(_02934__PTR8), .Z(_02938__PTR16) );
  XOR2_X1 U14726 ( .A(_02084__PTR17), .B(_02934__PTR8), .Z(_02938__PTR17) );
  XOR2_X1 U14727 ( .A(_02084__PTR18), .B(_02934__PTR8), .Z(_02938__PTR18) );
  XOR2_X1 U14728 ( .A(_02084__PTR19), .B(_02934__PTR8), .Z(_02938__PTR19) );
  XOR2_X1 U14729 ( .A(_02084__PTR20), .B(_02934__PTR8), .Z(_02938__PTR20) );
  XOR2_X1 U14730 ( .A(_02084__PTR21), .B(_02934__PTR8), .Z(_02938__PTR21) );
  XOR2_X1 U14731 ( .A(_02084__PTR22), .B(_02934__PTR8), .Z(_02938__PTR22) );
  XOR2_X1 U14732 ( .A(_02084__PTR23), .B(_02934__PTR8), .Z(_02938__PTR23) );
  XOR2_X1 U14733 ( .A(_02084__PTR24), .B(_02934__PTR8), .Z(_02938__PTR24) );
  XOR2_X1 U14734 ( .A(_02084__PTR25), .B(_02934__PTR8), .Z(_02938__PTR25) );
  XOR2_X1 U14735 ( .A(_02084__PTR26), .B(_02934__PTR8), .Z(_02938__PTR26) );
  XOR2_X1 U14736 ( .A(_02084__PTR27), .B(_02934__PTR8), .Z(_02938__PTR27) );
  XOR2_X1 U14737 ( .A(_02084__PTR28), .B(_02934__PTR8), .Z(_02938__PTR28) );
  XOR2_X1 U14738 ( .A(_02084__PTR29), .B(_02934__PTR8), .Z(_02938__PTR29) );
  XOR2_X1 U14739 ( .A(_02084__PTR30), .B(_02934__PTR8), .Z(_02938__PTR30) );
  XOR2_X1 U14740 ( .A(_02084__PTR31), .B(_02934__PTR8), .Z(_02938__PTR32) );
  AND2_X1 U14741 ( .A1(_02084__PTR2), .A2(_01885__PTR2), .ZN(_02940__PTR2) );
  AND2_X1 U14742 ( .A1(_02084__PTR3), .A2(_01885__PTR3), .ZN(_02940__PTR3) );
  AND2_X1 U14743 ( .A1(_02084__PTR4), .A2(_02936__PTR4), .ZN(_02940__PTR4) );
  AND2_X1 U14744 ( .A1(_02084__PTR5), .A2(_02936__PTR5), .ZN(_02940__PTR5) );
  AND2_X1 U14745 ( .A1(_02084__PTR6), .A2(_02936__PTR6), .ZN(_02940__PTR6) );
  AND2_X1 U14746 ( .A1(_02084__PTR7), .A2(_02936__PTR7), .ZN(_02940__PTR7) );
  AND2_X1 U14747 ( .A1(_02084__PTR8), .A2(_02934__PTR8), .ZN(_02940__PTR8) );
  AND2_X1 U14748 ( .A1(_02084__PTR9), .A2(_02934__PTR8), .ZN(_02940__PTR9) );
  AND2_X1 U14749 ( .A1(_02084__PTR10), .A2(_02934__PTR8), .ZN(_02940__PTR10) );
  AND2_X1 U14750 ( .A1(_02084__PTR11), .A2(_02934__PTR8), .ZN(_02940__PTR11) );
  AND2_X1 U14751 ( .A1(_02084__PTR12), .A2(_02934__PTR8), .ZN(_02940__PTR12) );
  AND2_X1 U14752 ( .A1(_02084__PTR13), .A2(_02934__PTR8), .ZN(_02940__PTR13) );
  AND2_X1 U14753 ( .A1(_02084__PTR14), .A2(_02934__PTR8), .ZN(_02940__PTR14) );
  AND2_X1 U14754 ( .A1(_02084__PTR15), .A2(_02934__PTR8), .ZN(_02940__PTR15) );
  AND2_X1 U14755 ( .A1(_02084__PTR16), .A2(_02934__PTR8), .ZN(_02940__PTR16) );
  AND2_X1 U14756 ( .A1(_02084__PTR17), .A2(_02934__PTR8), .ZN(_02940__PTR17) );
  AND2_X1 U14757 ( .A1(_02084__PTR18), .A2(_02934__PTR8), .ZN(_02940__PTR18) );
  AND2_X1 U14758 ( .A1(_02084__PTR19), .A2(_02934__PTR8), .ZN(_02940__PTR19) );
  AND2_X1 U14759 ( .A1(_02084__PTR20), .A2(_02934__PTR8), .ZN(_02940__PTR20) );
  AND2_X1 U14760 ( .A1(_02084__PTR21), .A2(_02934__PTR8), .ZN(_02940__PTR21) );
  AND2_X1 U14761 ( .A1(_02084__PTR22), .A2(_02934__PTR8), .ZN(_02940__PTR22) );
  AND2_X1 U14762 ( .A1(_02084__PTR23), .A2(_02934__PTR8), .ZN(_02940__PTR23) );
  AND2_X1 U14763 ( .A1(_02084__PTR24), .A2(_02934__PTR8), .ZN(_02940__PTR24) );
  AND2_X1 U14764 ( .A1(_02084__PTR25), .A2(_02934__PTR8), .ZN(_02940__PTR25) );
  AND2_X1 U14765 ( .A1(_02084__PTR26), .A2(_02934__PTR8), .ZN(_02940__PTR26) );
  AND2_X1 U14766 ( .A1(_02084__PTR27), .A2(_02934__PTR8), .ZN(_02940__PTR27) );
  AND2_X1 U14767 ( .A1(_02084__PTR28), .A2(_02934__PTR8), .ZN(_02940__PTR28) );
  AND2_X1 U14768 ( .A1(_02084__PTR29), .A2(_02934__PTR8), .ZN(_02940__PTR29) );
  AND2_X1 U14769 ( .A1(_02084__PTR30), .A2(_02934__PTR8), .ZN(_02940__PTR30) );
  XOR2_X1 U14770 ( .A(_01885__PTR4), .B(_02724__PTR3), .Z(_02725__PTR4) );
  XOR2_X1 U14771 ( .A(_01885__PTR5), .B(_02724__PTR4), .Z(_02725__PTR5) );
  XOR2_X1 U14772 ( .A(_01885__PTR6), .B(_02724__PTR5), .Z(_02725__PTR6) );
  XOR2_X1 U14773 ( .A(P1_P1_InstQueueRd_Addr_PTR1), .B(P1_P1_InstQueueRd_Addr_PTR0), .Z(_01884__PTR4) );
  XOR2_X1 U14774 ( .A(P1_P1_InstQueueRd_Addr_PTR2), .B(_02750__PTR1), .Z(_01884__PTR5) );
  XOR2_X1 U14775 ( .A(P1_P1_InstQueueRd_Addr_PTR4), .B(_02750__PTR3), .Z(_02800__PTR4) );
  XOR2_X1 U14776 ( .A(P1_P1_PhyAddrPointer_PTR2), .B(P1_P1_PhyAddrPointer_PTR1), .Z(_01892__PTR130) );
  XOR2_X1 U14777 ( .A(P1_P1_PhyAddrPointer_PTR3), .B(_02797__PTR1), .Z(_01892__PTR131) );
  XOR2_X1 U14778 ( .A(P1_P1_PhyAddrPointer_PTR4), .B(_02797__PTR2), .Z(_01892__PTR132) );
  XOR2_X1 U14779 ( .A(P1_P1_PhyAddrPointer_PTR5), .B(_02797__PTR3), .Z(_01892__PTR133) );
  XOR2_X1 U14780 ( .A(P1_P1_PhyAddrPointer_PTR6), .B(_02797__PTR4), .Z(_01892__PTR134) );
  XOR2_X1 U14781 ( .A(P1_P1_PhyAddrPointer_PTR7), .B(_02797__PTR5), .Z(_01892__PTR135) );
  XOR2_X1 U14782 ( .A(P1_P1_PhyAddrPointer_PTR8), .B(_02797__PTR6), .Z(_01892__PTR136) );
  XOR2_X1 U14783 ( .A(P1_P1_PhyAddrPointer_PTR9), .B(_02797__PTR7), .Z(_01892__PTR137) );
  XOR2_X1 U14784 ( .A(P1_P1_PhyAddrPointer_PTR10), .B(_02797__PTR8), .Z(_01892__PTR138) );
  XOR2_X1 U14785 ( .A(P1_P1_PhyAddrPointer_PTR11), .B(_02797__PTR9), .Z(_01892__PTR139) );
  XOR2_X1 U14786 ( .A(P1_P1_PhyAddrPointer_PTR12), .B(_02797__PTR10), .Z(_01892__PTR140) );
  XOR2_X1 U14787 ( .A(P1_P1_PhyAddrPointer_PTR13), .B(_02797__PTR11), .Z(_01892__PTR141) );
  XOR2_X1 U14788 ( .A(P1_P1_PhyAddrPointer_PTR14), .B(_02797__PTR12), .Z(_01892__PTR142) );
  XOR2_X1 U14789 ( .A(P1_P1_PhyAddrPointer_PTR15), .B(_02797__PTR13), .Z(_01892__PTR143) );
  XOR2_X1 U14790 ( .A(P1_P1_PhyAddrPointer_PTR16), .B(_02797__PTR14), .Z(_01892__PTR144) );
  XOR2_X1 U14791 ( .A(P1_P1_PhyAddrPointer_PTR17), .B(_02797__PTR15), .Z(_01892__PTR145) );
  XOR2_X1 U14792 ( .A(P1_P1_PhyAddrPointer_PTR18), .B(_02797__PTR16), .Z(_01892__PTR146) );
  XOR2_X1 U14793 ( .A(P1_P1_PhyAddrPointer_PTR19), .B(_02797__PTR17), .Z(_01892__PTR147) );
  XOR2_X1 U14794 ( .A(P1_P1_PhyAddrPointer_PTR20), .B(_02797__PTR18), .Z(_01892__PTR148) );
  XOR2_X1 U14795 ( .A(P1_P1_PhyAddrPointer_PTR21), .B(_02797__PTR19), .Z(_01892__PTR149) );
  XOR2_X1 U14796 ( .A(P1_P1_PhyAddrPointer_PTR22), .B(_02797__PTR20), .Z(_01892__PTR150) );
  XOR2_X1 U14797 ( .A(P1_P1_PhyAddrPointer_PTR23), .B(_02797__PTR21), .Z(_01892__PTR151) );
  XOR2_X1 U14798 ( .A(P1_P1_PhyAddrPointer_PTR24), .B(_02797__PTR22), .Z(_01892__PTR152) );
  XOR2_X1 U14799 ( .A(P1_P1_PhyAddrPointer_PTR25), .B(_02797__PTR23), .Z(_01892__PTR153) );
  XOR2_X1 U14800 ( .A(P1_P1_PhyAddrPointer_PTR26), .B(_02797__PTR24), .Z(_01892__PTR154) );
  XOR2_X1 U14801 ( .A(P1_P1_PhyAddrPointer_PTR27), .B(_02797__PTR25), .Z(_01892__PTR155) );
  XOR2_X1 U14802 ( .A(P1_P1_PhyAddrPointer_PTR28), .B(_02797__PTR26), .Z(_01892__PTR156) );
  XOR2_X1 U14803 ( .A(P1_P1_PhyAddrPointer_PTR29), .B(_02797__PTR27), .Z(_01892__PTR157) );
  XOR2_X1 U14804 ( .A(P1_P1_PhyAddrPointer_PTR30), .B(_02797__PTR28), .Z(_01892__PTR158) );
  XOR2_X1 U14805 ( .A(P1_P1_PhyAddrPointer_PTR31), .B(_02797__PTR29), .Z(_01892__PTR159) );
  XOR2_X1 U14806 ( .A(P1_P1_PhyAddrPointer_PTR1), .B(_02715__PTR0), .Z(_02946__PTR1) );
  XOR2_X1 U14807 ( .A(_02715__PTR2), .B(_02945__PTR1), .Z(_02946__PTR2) );
  XOR2_X1 U14808 ( .A(_02715__PTR3), .B(_02945__PTR2), .Z(_02946__PTR3) );
  XOR2_X1 U14809 ( .A(_02715__PTR4), .B(_02945__PTR3), .Z(_02946__PTR4) );
  XOR2_X1 U14810 ( .A(_02715__PTR5), .B(_02945__PTR4), .Z(_02946__PTR5) );
  XOR2_X1 U14811 ( .A(_02715__PTR6), .B(_02945__PTR5), .Z(_02946__PTR6) );
  XOR2_X1 U14812 ( .A(_02715__PTR7), .B(_02945__PTR6), .Z(_02946__PTR7) );
  XOR2_X1 U14813 ( .A(_02715__PTR8), .B(_02945__PTR7), .Z(_02946__PTR8) );
  XOR2_X1 U14814 ( .A(_02715__PTR9), .B(_02945__PTR8), .Z(_02946__PTR9) );
  XOR2_X1 U14815 ( .A(_02715__PTR10), .B(_02945__PTR9), .Z(_02946__PTR10) );
  XOR2_X1 U14816 ( .A(_02715__PTR11), .B(_02945__PTR10), .Z(_02946__PTR11) );
  XOR2_X1 U14817 ( .A(_02715__PTR12), .B(_02945__PTR11), .Z(_02946__PTR12) );
  XOR2_X1 U14818 ( .A(_02715__PTR13), .B(_02945__PTR12), .Z(_02946__PTR13) );
  XOR2_X1 U14819 ( .A(_02715__PTR14), .B(_02945__PTR13), .Z(_02946__PTR14) );
  XOR2_X1 U14820 ( .A(_02715__PTR15), .B(_02945__PTR14), .Z(_02946__PTR15) );
  XOR2_X1 U14821 ( .A(_02715__PTR16), .B(_02945__PTR15), .Z(_02946__PTR16) );
  XOR2_X1 U14822 ( .A(_02715__PTR17), .B(_02945__PTR16), .Z(_02946__PTR17) );
  XOR2_X1 U14823 ( .A(_02715__PTR18), .B(_02945__PTR17), .Z(_02946__PTR18) );
  XOR2_X1 U14824 ( .A(_02715__PTR19), .B(_02945__PTR18), .Z(_02946__PTR19) );
  XOR2_X1 U14825 ( .A(_02715__PTR20), .B(_02945__PTR19), .Z(_02946__PTR20) );
  XOR2_X1 U14826 ( .A(_02715__PTR21), .B(_02945__PTR20), .Z(_02946__PTR21) );
  XOR2_X1 U14827 ( .A(_02715__PTR22), .B(_02945__PTR21), .Z(_02946__PTR22) );
  XOR2_X1 U14828 ( .A(_02715__PTR23), .B(_02945__PTR22), .Z(_02946__PTR23) );
  XOR2_X1 U14829 ( .A(_02715__PTR24), .B(_02945__PTR23), .Z(_02946__PTR24) );
  XOR2_X1 U14830 ( .A(_02715__PTR25), .B(_02945__PTR24), .Z(_02946__PTR25) );
  XOR2_X1 U14831 ( .A(_02715__PTR26), .B(_02945__PTR25), .Z(_02946__PTR26) );
  XOR2_X1 U14832 ( .A(_02715__PTR27), .B(_02945__PTR26), .Z(_02946__PTR27) );
  XOR2_X1 U14833 ( .A(_02715__PTR28), .B(_02945__PTR27), .Z(_02946__PTR28) );
  XOR2_X1 U14834 ( .A(_02715__PTR29), .B(_02945__PTR28), .Z(_02946__PTR29) );
  XOR2_X1 U14835 ( .A(_02715__PTR30), .B(_02945__PTR29), .Z(_02946__PTR30) );
  XOR2_X1 U14836 ( .A(_02713__PTR31), .B(_02945__PTR30), .Z(_02946__PTR31) );
  XOR2_X1 U14837 ( .A(P1_P1_PhyAddrPointer_PTR3), .B(P1_P1_PhyAddrPointer_PTR2), .Z(_02796__PTR1) );
  XOR2_X1 U14838 ( .A(P1_P1_PhyAddrPointer_PTR4), .B(_02794__PTR1), .Z(_02796__PTR2) );
  XOR2_X1 U14839 ( .A(P1_P1_PhyAddrPointer_PTR5), .B(_02794__PTR2), .Z(_02796__PTR3) );
  XOR2_X1 U14840 ( .A(P1_P1_PhyAddrPointer_PTR6), .B(_02794__PTR3), .Z(_02796__PTR4) );
  XOR2_X1 U14841 ( .A(P1_P1_PhyAddrPointer_PTR7), .B(_02794__PTR4), .Z(_02796__PTR5) );
  XOR2_X1 U14842 ( .A(P1_P1_PhyAddrPointer_PTR8), .B(_02794__PTR5), .Z(_02796__PTR6) );
  XOR2_X1 U14843 ( .A(P1_P1_PhyAddrPointer_PTR9), .B(_02794__PTR6), .Z(_02796__PTR7) );
  XOR2_X1 U14844 ( .A(P1_P1_PhyAddrPointer_PTR10), .B(_02794__PTR7), .Z(_02796__PTR8) );
  XOR2_X1 U14845 ( .A(P1_P1_PhyAddrPointer_PTR11), .B(_02794__PTR8), .Z(_02796__PTR9) );
  XOR2_X1 U14846 ( .A(P1_P1_PhyAddrPointer_PTR12), .B(_02794__PTR9), .Z(_02796__PTR10) );
  XOR2_X1 U14847 ( .A(P1_P1_PhyAddrPointer_PTR13), .B(_02794__PTR10), .Z(_02796__PTR11) );
  XOR2_X1 U14848 ( .A(P1_P1_PhyAddrPointer_PTR14), .B(_02794__PTR11), .Z(_02796__PTR12) );
  XOR2_X1 U14849 ( .A(P1_P1_PhyAddrPointer_PTR15), .B(_02794__PTR12), .Z(_02796__PTR13) );
  XOR2_X1 U14850 ( .A(P1_P1_PhyAddrPointer_PTR16), .B(_02794__PTR13), .Z(_02796__PTR14) );
  XOR2_X1 U14851 ( .A(P1_P1_PhyAddrPointer_PTR17), .B(_02794__PTR14), .Z(_02796__PTR15) );
  XOR2_X1 U14852 ( .A(P1_P1_PhyAddrPointer_PTR18), .B(_02794__PTR15), .Z(_02796__PTR16) );
  XOR2_X1 U14853 ( .A(P1_P1_PhyAddrPointer_PTR19), .B(_02794__PTR16), .Z(_02796__PTR17) );
  XOR2_X1 U14854 ( .A(P1_P1_PhyAddrPointer_PTR20), .B(_02794__PTR17), .Z(_02796__PTR18) );
  XOR2_X1 U14855 ( .A(P1_P1_PhyAddrPointer_PTR21), .B(_02794__PTR18), .Z(_02796__PTR19) );
  XOR2_X1 U14856 ( .A(P1_P1_PhyAddrPointer_PTR22), .B(_02794__PTR19), .Z(_02796__PTR20) );
  XOR2_X1 U14857 ( .A(P1_P1_PhyAddrPointer_PTR23), .B(_02794__PTR20), .Z(_02796__PTR21) );
  XOR2_X1 U14858 ( .A(P1_P1_PhyAddrPointer_PTR24), .B(_02794__PTR21), .Z(_02796__PTR22) );
  XOR2_X1 U14859 ( .A(P1_P1_PhyAddrPointer_PTR25), .B(_02794__PTR22), .Z(_02796__PTR23) );
  XOR2_X1 U14860 ( .A(P1_P1_PhyAddrPointer_PTR26), .B(_02794__PTR23), .Z(_02796__PTR24) );
  XOR2_X1 U14861 ( .A(P1_P1_PhyAddrPointer_PTR27), .B(_02794__PTR24), .Z(_02796__PTR25) );
  XOR2_X1 U14862 ( .A(P1_P1_PhyAddrPointer_PTR28), .B(_02794__PTR25), .Z(_02796__PTR26) );
  XOR2_X1 U14863 ( .A(P1_P1_PhyAddrPointer_PTR29), .B(_02794__PTR26), .Z(_02796__PTR27) );
  XOR2_X1 U14864 ( .A(P1_P1_PhyAddrPointer_PTR30), .B(_02794__PTR27), .Z(_02796__PTR28) );
  XOR2_X1 U14865 ( .A(P1_P1_PhyAddrPointer_PTR31), .B(_02794__PTR28), .Z(_02796__PTR29) );
  XOR2_X1 U14866 ( .A(P1_P1_InstQueueWr_Addr_PTR1), .B(P1_P1_InstQueueWr_Addr_PTR0), .Z(_01836__PTR1) );
  XOR2_X1 U14867 ( .A(P1_P1_InstQueueWr_Addr_PTR2), .B(_02779__PTR1), .Z(_01836__PTR2) );
  XOR2_X1 U14868 ( .A(P1_P1_InstQueueWr_Addr_PTR3), .B(_02779__PTR2), .Z(_01836__PTR3) );
  XOR2_X1 U14869 ( .A(_01836__PTR1), .B(_01836__PTR0), .Z(_01838__PTR1) );
  XOR2_X1 U14870 ( .A(_01836__PTR2), .B(_02780__PTR1), .Z(_01838__PTR2) );
  XOR2_X1 U14871 ( .A(_01836__PTR3), .B(_02780__PTR2), .Z(_01838__PTR3) );
  XOR2_X1 U14872 ( .A(_01838__PTR1), .B(P1_P1_InstQueueWr_Addr_PTR0), .Z(_01840__PTR1) );
  XOR2_X1 U14873 ( .A(_01838__PTR2), .B(_02785__PTR1), .Z(_01840__PTR2) );
  XOR2_X1 U14874 ( .A(_01838__PTR3), .B(_02785__PTR2), .Z(_01840__PTR3) );
  XOR2_X1 U14875 ( .A(_01840__PTR1), .B(_01836__PTR0), .Z(_02791__PTR1) );
  XOR2_X1 U14876 ( .A(_01840__PTR2), .B(_02790__PTR1), .Z(_02791__PTR2) );
  XOR2_X1 U14877 ( .A(_01840__PTR3), .B(_02790__PTR2), .Z(_02791__PTR3) );
  XOR2_X1 U14878 ( .A(di1_PTR25), .B(_02787__PTR0), .Z(_02789__PTR1) );
  XOR2_X1 U14879 ( .A(di1_PTR26), .B(_02787__PTR1), .Z(_02789__PTR2) );
  XOR2_X1 U14880 ( .A(di1_PTR27), .B(_02787__PTR2), .Z(_02789__PTR3) );
  XOR2_X1 U14881 ( .A(di1_PTR28), .B(_02787__PTR3), .Z(_02789__PTR4) );
  XOR2_X1 U14882 ( .A(di1_PTR29), .B(_02787__PTR4), .Z(_02789__PTR5) );
  XOR2_X1 U14883 ( .A(di1_PTR30), .B(_02787__PTR5), .Z(_02789__PTR6) );
  XOR2_X1 U14884 ( .A(P1_Datai_PTR31), .B(_02787__PTR6), .Z(_02789__PTR7) );
  XOR2_X1 U14885 ( .A(_02786_), .B(di1_PTR24), .Z(_02788__PTR0) );
  AND2_X1 U14886 ( .A1(_02786_), .A2(di1_PTR24), .ZN(_02787__PTR0) );
  XOR2_X1 U14887 ( .A(di1_PTR17), .B(_02782__PTR0), .Z(_02784__PTR1) );
  XOR2_X1 U14888 ( .A(di1_PTR18), .B(_02782__PTR1), .Z(_02784__PTR2) );
  XOR2_X1 U14889 ( .A(di1_PTR19), .B(_02782__PTR2), .Z(_02784__PTR3) );
  XOR2_X1 U14890 ( .A(di1_PTR20), .B(_02782__PTR3), .Z(_02784__PTR4) );
  XOR2_X1 U14891 ( .A(di1_PTR21), .B(_02782__PTR4), .Z(_02784__PTR5) );
  XOR2_X1 U14892 ( .A(di1_PTR22), .B(_02782__PTR5), .Z(_02784__PTR6) );
  XOR2_X1 U14893 ( .A(di1_PTR23), .B(_02782__PTR6), .Z(_02784__PTR7) );
  XOR2_X1 U14894 ( .A(_02781_), .B(di1_PTR16), .Z(_02783__PTR0) );
  AND2_X1 U14895 ( .A1(_02781_), .A2(di1_PTR16), .ZN(_02782__PTR0) );
  XOR2_X1 U14896 ( .A(P1_rEIP_PTR2), .B(_02778__PTR0), .Z(_01880__PTR193) );
  XOR2_X1 U14897 ( .A(P1_rEIP_PTR3), .B(_02778__PTR1), .Z(_01880__PTR194) );
  XOR2_X1 U14898 ( .A(P1_rEIP_PTR4), .B(_02778__PTR2), .Z(_01880__PTR195) );
  XOR2_X1 U14899 ( .A(P1_rEIP_PTR5), .B(_02778__PTR3), .Z(_01880__PTR196) );
  XOR2_X1 U14900 ( .A(P1_rEIP_PTR6), .B(_02778__PTR4), .Z(_01880__PTR197) );
  XOR2_X1 U14901 ( .A(P1_rEIP_PTR7), .B(_02778__PTR5), .Z(_01880__PTR198) );
  XOR2_X1 U14902 ( .A(P1_rEIP_PTR8), .B(_02778__PTR6), .Z(_01880__PTR199) );
  XOR2_X1 U14903 ( .A(P1_rEIP_PTR9), .B(_02778__PTR7), .Z(_01880__PTR200) );
  XOR2_X1 U14904 ( .A(P1_rEIP_PTR10), .B(_02778__PTR8), .Z(_01880__PTR201) );
  XOR2_X1 U14905 ( .A(P1_rEIP_PTR11), .B(_02778__PTR9), .Z(_01880__PTR202) );
  XOR2_X1 U14906 ( .A(P1_rEIP_PTR12), .B(_02778__PTR10), .Z(_01880__PTR203) );
  XOR2_X1 U14907 ( .A(P1_rEIP_PTR13), .B(_02778__PTR11), .Z(_01880__PTR204) );
  XOR2_X1 U14908 ( .A(P1_rEIP_PTR14), .B(_02778__PTR12), .Z(_01880__PTR205) );
  XOR2_X1 U14909 ( .A(P1_rEIP_PTR15), .B(_02778__PTR13), .Z(_01880__PTR206) );
  XOR2_X1 U14910 ( .A(P1_rEIP_PTR16), .B(_02778__PTR14), .Z(_01880__PTR207) );
  XOR2_X1 U14911 ( .A(P1_rEIP_PTR17), .B(_02778__PTR15), .Z(_01880__PTR208) );
  XOR2_X1 U14912 ( .A(P1_rEIP_PTR18), .B(_02778__PTR16), .Z(_01880__PTR209) );
  XOR2_X1 U14913 ( .A(P1_rEIP_PTR19), .B(_02778__PTR17), .Z(_01880__PTR210) );
  XOR2_X1 U14914 ( .A(P1_rEIP_PTR20), .B(_02778__PTR18), .Z(_01880__PTR211) );
  XOR2_X1 U14915 ( .A(P1_rEIP_PTR21), .B(_02778__PTR19), .Z(_01880__PTR212) );
  XOR2_X1 U14916 ( .A(P1_rEIP_PTR22), .B(_02778__PTR20), .Z(_01880__PTR213) );
  XOR2_X1 U14917 ( .A(P1_rEIP_PTR23), .B(_02778__PTR21), .Z(_01880__PTR214) );
  XOR2_X1 U14918 ( .A(P1_rEIP_PTR24), .B(_02778__PTR22), .Z(_01880__PTR215) );
  XOR2_X1 U14919 ( .A(P1_rEIP_PTR25), .B(_02778__PTR23), .Z(_01880__PTR216) );
  XOR2_X1 U14920 ( .A(P1_rEIP_PTR26), .B(_02778__PTR24), .Z(_01880__PTR217) );
  XOR2_X1 U14921 ( .A(P1_rEIP_PTR27), .B(_02778__PTR25), .Z(_01880__PTR218) );
  XOR2_X1 U14922 ( .A(P1_rEIP_PTR28), .B(_02778__PTR26), .Z(_01880__PTR219) );
  XOR2_X1 U14923 ( .A(P1_rEIP_PTR29), .B(_02778__PTR27), .Z(_01880__PTR220) );
  XOR2_X1 U14924 ( .A(P1_rEIP_PTR30), .B(_02778__PTR28), .Z(_01880__PTR221) );
  XOR2_X1 U14925 ( .A(_02777_), .B(P1_rEIP_PTR1), .Z(_01880__PTR192) );
  AND2_X1 U14926 ( .A1(_02777_), .A2(P1_rEIP_PTR1), .ZN(_02778__PTR0) );
  XOR2_X1 U14927 ( .A(P1_rEIP_PTR3), .B(_02793__PTR0), .Z(_01880__PTR65) );
  XOR2_X1 U14928 ( .A(P1_rEIP_PTR4), .B(_02793__PTR1), .Z(_01880__PTR66) );
  XOR2_X1 U14929 ( .A(P1_rEIP_PTR5), .B(_02793__PTR2), .Z(_01880__PTR67) );
  XOR2_X1 U14930 ( .A(P1_rEIP_PTR6), .B(_02793__PTR3), .Z(_01880__PTR68) );
  XOR2_X1 U14931 ( .A(P1_rEIP_PTR7), .B(_02793__PTR4), .Z(_01880__PTR69) );
  XOR2_X1 U14932 ( .A(P1_rEIP_PTR8), .B(_02793__PTR5), .Z(_01880__PTR70) );
  XOR2_X1 U14933 ( .A(P1_rEIP_PTR9), .B(_02793__PTR6), .Z(_01880__PTR71) );
  XOR2_X1 U14934 ( .A(P1_rEIP_PTR10), .B(_02793__PTR7), .Z(_01880__PTR72) );
  XOR2_X1 U14935 ( .A(P1_rEIP_PTR11), .B(_02793__PTR8), .Z(_01880__PTR73) );
  XOR2_X1 U14936 ( .A(P1_rEIP_PTR12), .B(_02793__PTR9), .Z(_01880__PTR74) );
  XOR2_X1 U14937 ( .A(P1_rEIP_PTR13), .B(_02793__PTR10), .Z(_01880__PTR75) );
  XOR2_X1 U14938 ( .A(P1_rEIP_PTR14), .B(_02793__PTR11), .Z(_01880__PTR76) );
  XOR2_X1 U14939 ( .A(P1_rEIP_PTR15), .B(_02793__PTR12), .Z(_01880__PTR77) );
  XOR2_X1 U14940 ( .A(P1_rEIP_PTR16), .B(_02793__PTR13), .Z(_01880__PTR78) );
  XOR2_X1 U14941 ( .A(P1_rEIP_PTR17), .B(_02793__PTR14), .Z(_01880__PTR79) );
  XOR2_X1 U14942 ( .A(P1_rEIP_PTR18), .B(_02793__PTR15), .Z(_01880__PTR80) );
  XOR2_X1 U14943 ( .A(P1_rEIP_PTR19), .B(_02793__PTR16), .Z(_01880__PTR81) );
  XOR2_X1 U14944 ( .A(P1_rEIP_PTR20), .B(_02793__PTR17), .Z(_01880__PTR82) );
  XOR2_X1 U14945 ( .A(P1_rEIP_PTR21), .B(_02793__PTR18), .Z(_01880__PTR83) );
  XOR2_X1 U14946 ( .A(P1_rEIP_PTR22), .B(_02793__PTR19), .Z(_01880__PTR84) );
  XOR2_X1 U14947 ( .A(P1_rEIP_PTR23), .B(_02793__PTR20), .Z(_01880__PTR85) );
  XOR2_X1 U14948 ( .A(P1_rEIP_PTR24), .B(_02793__PTR21), .Z(_01880__PTR86) );
  XOR2_X1 U14949 ( .A(P1_rEIP_PTR25), .B(_02793__PTR22), .Z(_01880__PTR87) );
  XOR2_X1 U14950 ( .A(P1_rEIP_PTR26), .B(_02793__PTR23), .Z(_01880__PTR88) );
  XOR2_X1 U14951 ( .A(P1_rEIP_PTR27), .B(_02793__PTR24), .Z(_01880__PTR89) );
  XOR2_X1 U14952 ( .A(P1_rEIP_PTR28), .B(_02793__PTR25), .Z(_01880__PTR90) );
  XOR2_X1 U14953 ( .A(P1_rEIP_PTR29), .B(_02793__PTR26), .Z(_01880__PTR91) );
  XOR2_X1 U14954 ( .A(P1_rEIP_PTR30), .B(_02793__PTR27), .Z(_01880__PTR92) );
  XOR2_X1 U14955 ( .A(P1_rEIP_PTR31), .B(_02793__PTR28), .Z(_01880__PTR93) );
  XOR2_X1 U14956 ( .A(_02792_), .B(P1_rEIP_PTR2), .Z(_01880__PTR64) );
  AND2_X1 U14957 ( .A1(_02792_), .A2(P1_rEIP_PTR2), .ZN(_02793__PTR0) );
  XOR2_X1 U14958 ( .A(P2_P1_InstQueueRd_Addr_PTR1), .B(P2_P1_InstQueueRd_Addr_PTR0), .Z(_02176__PTR4) );
  XOR2_X1 U14959 ( .A(_03188__PTR4), .B(_03189__PTR3), .Z(_02991__PTR4) );
  XOR2_X1 U14960 ( .A(_03074__PTR1), .B(P2_P1_InstAddrPointer_PTR0), .Z(_03076__PTR1) );
  XOR2_X1 U14961 ( .A(_02373__PTR33), .B(_02373__PTR0), .Z(_03194__PTR1) );
  XOR2_X1 U14962 ( .A(_03186__PTR4), .B(_03187__PTR3), .Z(_02984__PTR4) );
  XOR2_X1 U14963 ( .A(_02224__PTR40), .B(_02129__PTR0), .Z(_02982__PTR0) );
  XOR2_X1 U14964 ( .A(_02224__PTR41), .B(_02980__PTR1), .Z(_02982__PTR1) );
  XOR2_X1 U14965 ( .A(_02224__PTR42), .B(_02980__PTR2), .Z(_02982__PTR2) );
  XOR2_X1 U14966 ( .A(_02224__PTR43), .B(_02980__PTR3), .Z(_02982__PTR3) );
  XOR2_X1 U14967 ( .A(_02224__PTR44), .B(_02980__PTR4), .Z(_02982__PTR4) );
  AND2_X1 U14968 ( .A1(_02224__PTR40), .A2(_02129__PTR0), .ZN(_02983__PTR0) );
  AND2_X1 U14969 ( .A1(_02224__PTR41), .A2(_02980__PTR1), .ZN(_02983__PTR1) );
  AND2_X1 U14970 ( .A1(_02224__PTR42), .A2(_02980__PTR2), .ZN(_02983__PTR2) );
  AND2_X1 U14971 ( .A1(_02224__PTR43), .A2(_02980__PTR3), .ZN(_02983__PTR3) );
  AND2_X1 U14972 ( .A1(_02224__PTR44), .A2(_02980__PTR4), .ZN(_02983__PTR4) );
  XOR2_X1 U14973 ( .A(P2_EBX_PTR1), .B(P2_EBX_PTR0), .Z(_02389__PTR33) );
  XOR2_X1 U14974 ( .A(P2_EBX_PTR2), .B(_03073__PTR1), .Z(_02389__PTR34) );
  XOR2_X1 U14975 ( .A(P2_EBX_PTR3), .B(_03073__PTR2), .Z(_02389__PTR35) );
  XOR2_X1 U14976 ( .A(P2_EBX_PTR4), .B(_03073__PTR3), .Z(_02389__PTR36) );
  XOR2_X1 U14977 ( .A(P2_EBX_PTR5), .B(_03073__PTR4), .Z(_02389__PTR37) );
  XOR2_X1 U14978 ( .A(P2_EBX_PTR6), .B(_03073__PTR5), .Z(_02389__PTR38) );
  XOR2_X1 U14979 ( .A(P2_EBX_PTR7), .B(_03073__PTR6), .Z(_02389__PTR39) );
  XOR2_X1 U14980 ( .A(P2_EBX_PTR8), .B(_03073__PTR7), .Z(_02389__PTR40) );
  XOR2_X1 U14981 ( .A(P2_EBX_PTR9), .B(_03073__PTR8), .Z(_02389__PTR41) );
  XOR2_X1 U14982 ( .A(P2_EBX_PTR10), .B(_03073__PTR9), .Z(_02389__PTR42) );
  XOR2_X1 U14983 ( .A(P2_EBX_PTR11), .B(_03073__PTR10), .Z(_02389__PTR43) );
  XOR2_X1 U14984 ( .A(P2_EBX_PTR12), .B(_03073__PTR11), .Z(_02389__PTR44) );
  XOR2_X1 U14985 ( .A(P2_EBX_PTR13), .B(_03073__PTR12), .Z(_02389__PTR45) );
  XOR2_X1 U14986 ( .A(P2_EBX_PTR14), .B(_03073__PTR13), .Z(_02389__PTR46) );
  XOR2_X1 U14987 ( .A(P2_EBX_PTR15), .B(_03073__PTR14), .Z(_02389__PTR47) );
  XOR2_X1 U14988 ( .A(P2_EBX_PTR16), .B(_03073__PTR15), .Z(_02389__PTR48) );
  XOR2_X1 U14989 ( .A(P2_EBX_PTR17), .B(_03073__PTR16), .Z(_02389__PTR49) );
  XOR2_X1 U14990 ( .A(P2_EBX_PTR18), .B(_03073__PTR17), .Z(_02389__PTR50) );
  XOR2_X1 U14991 ( .A(P2_EBX_PTR19), .B(_03073__PTR18), .Z(_02389__PTR51) );
  XOR2_X1 U14992 ( .A(P2_EBX_PTR20), .B(_03073__PTR19), .Z(_02389__PTR52) );
  XOR2_X1 U14993 ( .A(P2_EBX_PTR21), .B(_03073__PTR20), .Z(_02389__PTR53) );
  XOR2_X1 U14994 ( .A(P2_EBX_PTR22), .B(_03073__PTR21), .Z(_02389__PTR54) );
  XOR2_X1 U14995 ( .A(P2_EBX_PTR23), .B(_03073__PTR22), .Z(_02389__PTR55) );
  XOR2_X1 U14996 ( .A(P2_EBX_PTR24), .B(_03073__PTR23), .Z(_02389__PTR56) );
  XOR2_X1 U14997 ( .A(P2_EBX_PTR25), .B(_03073__PTR24), .Z(_02389__PTR57) );
  XOR2_X1 U14998 ( .A(P2_EBX_PTR26), .B(_03073__PTR25), .Z(_02389__PTR58) );
  XOR2_X1 U14999 ( .A(P2_EBX_PTR27), .B(_03073__PTR26), .Z(_02389__PTR59) );
  XOR2_X1 U15000 ( .A(P2_EBX_PTR28), .B(_03073__PTR27), .Z(_02389__PTR60) );
  XOR2_X1 U15001 ( .A(P2_EBX_PTR29), .B(_03073__PTR28), .Z(_02389__PTR61) );
  XOR2_X1 U15002 ( .A(P2_EBX_PTR30), .B(_03073__PTR29), .Z(_02389__PTR62) );
  XOR2_X1 U15003 ( .A(P2_EBX_PTR31), .B(_03073__PTR30), .Z(_02389__PTR63) );
  XOR2_X1 U15004 ( .A(P2_EAX_PTR1), .B(P2_EAX_PTR0), .Z(_02385__PTR33) );
  XOR2_X1 U15005 ( .A(P2_EAX_PTR2), .B(_03072__PTR1), .Z(_02385__PTR34) );
  XOR2_X1 U15006 ( .A(P2_EAX_PTR3), .B(_03072__PTR2), .Z(_02385__PTR35) );
  XOR2_X1 U15007 ( .A(P2_EAX_PTR4), .B(_03072__PTR3), .Z(_02385__PTR36) );
  XOR2_X1 U15008 ( .A(P2_EAX_PTR5), .B(_03072__PTR4), .Z(_02385__PTR37) );
  XOR2_X1 U15009 ( .A(P2_EAX_PTR6), .B(_03072__PTR5), .Z(_02385__PTR38) );
  XOR2_X1 U15010 ( .A(P2_EAX_PTR7), .B(_03072__PTR6), .Z(_02385__PTR39) );
  XOR2_X1 U15011 ( .A(P2_EAX_PTR8), .B(_03072__PTR7), .Z(_02385__PTR40) );
  XOR2_X1 U15012 ( .A(P2_EAX_PTR9), .B(_03072__PTR8), .Z(_02385__PTR41) );
  XOR2_X1 U15013 ( .A(P2_EAX_PTR10), .B(_03072__PTR9), .Z(_02385__PTR42) );
  XOR2_X1 U15014 ( .A(P2_EAX_PTR11), .B(_03072__PTR10), .Z(_02385__PTR43) );
  XOR2_X1 U15015 ( .A(P2_EAX_PTR12), .B(_03072__PTR11), .Z(_02385__PTR44) );
  XOR2_X1 U15016 ( .A(P2_EAX_PTR13), .B(_03072__PTR12), .Z(_02385__PTR45) );
  XOR2_X1 U15017 ( .A(P2_EAX_PTR14), .B(_03072__PTR13), .Z(_02385__PTR46) );
  XOR2_X1 U15018 ( .A(P2_EAX_PTR15), .B(_03072__PTR14), .Z(_02385__PTR47) );
  XOR2_X1 U15019 ( .A(P2_EAX_PTR16), .B(_03072__PTR15), .Z(_02385__PTR48) );
  XOR2_X1 U15020 ( .A(P2_EAX_PTR17), .B(_03072__PTR16), .Z(_02385__PTR49) );
  XOR2_X1 U15021 ( .A(P2_EAX_PTR18), .B(_03072__PTR17), .Z(_02385__PTR50) );
  XOR2_X1 U15022 ( .A(P2_EAX_PTR19), .B(_03072__PTR18), .Z(_02385__PTR51) );
  XOR2_X1 U15023 ( .A(P2_EAX_PTR20), .B(_03072__PTR19), .Z(_02385__PTR52) );
  XOR2_X1 U15024 ( .A(P2_EAX_PTR21), .B(_03072__PTR20), .Z(_02385__PTR53) );
  XOR2_X1 U15025 ( .A(P2_EAX_PTR22), .B(_03072__PTR21), .Z(_02385__PTR54) );
  XOR2_X1 U15026 ( .A(P2_EAX_PTR23), .B(_03072__PTR22), .Z(_02385__PTR55) );
  XOR2_X1 U15027 ( .A(P2_EAX_PTR24), .B(_03072__PTR23), .Z(_02385__PTR56) );
  XOR2_X1 U15028 ( .A(P2_EAX_PTR25), .B(_03072__PTR24), .Z(_02385__PTR57) );
  XOR2_X1 U15029 ( .A(P2_EAX_PTR26), .B(_03072__PTR25), .Z(_02385__PTR58) );
  XOR2_X1 U15030 ( .A(P2_EAX_PTR27), .B(_03072__PTR26), .Z(_02385__PTR59) );
  XOR2_X1 U15031 ( .A(P2_EAX_PTR28), .B(_03072__PTR27), .Z(_02385__PTR60) );
  XOR2_X1 U15032 ( .A(P2_EAX_PTR29), .B(_03072__PTR28), .Z(_02385__PTR61) );
  XOR2_X1 U15033 ( .A(P2_EAX_PTR30), .B(_03072__PTR29), .Z(_02385__PTR62) );
  XOR2_X1 U15034 ( .A(P2_EAX_PTR31), .B(_03072__PTR30), .Z(_02385__PTR63) );
  XOR2_X1 U15035 ( .A(P2_EAX_PTR17), .B(_03069__PTR0), .Z(_03071__PTR1) );
  XOR2_X1 U15036 ( .A(P2_EAX_PTR18), .B(_03069__PTR1), .Z(_03071__PTR2) );
  XOR2_X1 U15037 ( .A(P2_EAX_PTR19), .B(_03069__PTR2), .Z(_03071__PTR3) );
  XOR2_X1 U15038 ( .A(P2_EAX_PTR20), .B(_03069__PTR3), .Z(_03071__PTR4) );
  XOR2_X1 U15039 ( .A(P2_EAX_PTR21), .B(_03069__PTR4), .Z(_03071__PTR5) );
  XOR2_X1 U15040 ( .A(P2_EAX_PTR22), .B(_03069__PTR5), .Z(_03071__PTR6) );
  XOR2_X1 U15041 ( .A(P2_EAX_PTR23), .B(_03069__PTR6), .Z(_03071__PTR7) );
  XOR2_X1 U15042 ( .A(P2_EAX_PTR24), .B(_03069__PTR7), .Z(_03071__PTR8) );
  XOR2_X1 U15043 ( .A(P2_EAX_PTR25), .B(_03069__PTR8), .Z(_03071__PTR9) );
  XOR2_X1 U15044 ( .A(P2_EAX_PTR26), .B(_03069__PTR9), .Z(_03071__PTR10) );
  XOR2_X1 U15045 ( .A(P2_EAX_PTR27), .B(_03069__PTR10), .Z(_03071__PTR11) );
  XOR2_X1 U15046 ( .A(P2_EAX_PTR28), .B(_03069__PTR11), .Z(_03071__PTR12) );
  XOR2_X1 U15047 ( .A(P2_EAX_PTR29), .B(_03069__PTR12), .Z(_03071__PTR13) );
  XOR2_X1 U15048 ( .A(P2_EAX_PTR30), .B(_03069__PTR13), .Z(_03071__PTR14) );
  XOR2_X1 U15049 ( .A(_03068_), .B(P2_EAX_PTR16), .Z(_03070__PTR0) );
  AND2_X1 U15050 ( .A1(_03068_), .A2(P2_EAX_PTR16), .ZN(_03069__PTR0) );
  XOR2_X1 U15051 ( .A(P2_rEIP_PTR2), .B(P2_rEIP_PTR1), .Z(_03067__PTR1) );
  XOR2_X1 U15052 ( .A(P2_rEIP_PTR3), .B(_03066__PTR1), .Z(_03067__PTR2) );
  XOR2_X1 U15053 ( .A(P2_rEIP_PTR4), .B(_03066__PTR2), .Z(_03067__PTR3) );
  XOR2_X1 U15054 ( .A(P2_rEIP_PTR5), .B(_03066__PTR3), .Z(_03067__PTR4) );
  XOR2_X1 U15055 ( .A(P2_rEIP_PTR6), .B(_03066__PTR4), .Z(_03067__PTR5) );
  XOR2_X1 U15056 ( .A(P2_rEIP_PTR7), .B(_03066__PTR5), .Z(_03067__PTR6) );
  XOR2_X1 U15057 ( .A(P2_rEIP_PTR8), .B(_03066__PTR6), .Z(_03067__PTR7) );
  XOR2_X1 U15058 ( .A(P2_rEIP_PTR9), .B(_03066__PTR7), .Z(_03067__PTR8) );
  XOR2_X1 U15059 ( .A(P2_rEIP_PTR10), .B(_03066__PTR8), .Z(_03067__PTR9) );
  XOR2_X1 U15060 ( .A(P2_rEIP_PTR11), .B(_03066__PTR9), .Z(_03067__PTR10) );
  XOR2_X1 U15061 ( .A(P2_rEIP_PTR12), .B(_03066__PTR10), .Z(_03067__PTR11) );
  XOR2_X1 U15062 ( .A(P2_rEIP_PTR13), .B(_03066__PTR11), .Z(_03067__PTR12) );
  XOR2_X1 U15063 ( .A(P2_rEIP_PTR14), .B(_03066__PTR12), .Z(_03067__PTR13) );
  XOR2_X1 U15064 ( .A(P2_rEIP_PTR15), .B(_03066__PTR13), .Z(_03067__PTR14) );
  XOR2_X1 U15065 ( .A(P2_rEIP_PTR16), .B(_03066__PTR14), .Z(_03067__PTR15) );
  XOR2_X1 U15066 ( .A(P2_rEIP_PTR17), .B(_03066__PTR15), .Z(_03067__PTR16) );
  XOR2_X1 U15067 ( .A(P2_rEIP_PTR18), .B(_03066__PTR16), .Z(_03067__PTR17) );
  XOR2_X1 U15068 ( .A(P2_rEIP_PTR19), .B(_03066__PTR17), .Z(_03067__PTR18) );
  XOR2_X1 U15069 ( .A(P2_rEIP_PTR20), .B(_03066__PTR18), .Z(_03067__PTR19) );
  XOR2_X1 U15070 ( .A(P2_rEIP_PTR21), .B(_03066__PTR19), .Z(_03067__PTR20) );
  XOR2_X1 U15071 ( .A(P2_rEIP_PTR22), .B(_03066__PTR20), .Z(_03067__PTR21) );
  XOR2_X1 U15072 ( .A(P2_rEIP_PTR23), .B(_03066__PTR21), .Z(_03067__PTR22) );
  XOR2_X1 U15073 ( .A(P2_rEIP_PTR24), .B(_03066__PTR22), .Z(_03067__PTR23) );
  XOR2_X1 U15074 ( .A(P2_rEIP_PTR25), .B(_03066__PTR23), .Z(_03067__PTR24) );
  XOR2_X1 U15075 ( .A(P2_rEIP_PTR26), .B(_03066__PTR24), .Z(_03067__PTR25) );
  XOR2_X1 U15076 ( .A(P2_rEIP_PTR27), .B(_03066__PTR25), .Z(_03067__PTR26) );
  XOR2_X1 U15077 ( .A(P2_rEIP_PTR28), .B(_03066__PTR26), .Z(_03067__PTR27) );
  XOR2_X1 U15078 ( .A(P2_rEIP_PTR29), .B(_03066__PTR27), .Z(_03067__PTR28) );
  XOR2_X1 U15079 ( .A(P2_rEIP_PTR30), .B(_03066__PTR28), .Z(_03067__PTR29) );
  XOR2_X1 U15080 ( .A(P2_rEIP_PTR31), .B(_03066__PTR29), .Z(_03067__PTR30) );
  XOR2_X1 U15081 ( .A(_02979__PTR1), .B(_02389__PTR32), .Z(_03193__PTR1) );
  XOR2_X1 U15082 ( .A(_02979__PTR2), .B(_03192__PTR1), .Z(_03193__PTR2) );
  XOR2_X1 U15083 ( .A(_02979__PTR3), .B(_03192__PTR2), .Z(_03193__PTR3) );
  XOR2_X1 U15084 ( .A(_02979__PTR4), .B(_03192__PTR3), .Z(_03193__PTR4) );
  XOR2_X1 U15085 ( .A(_02979__PTR5), .B(_03192__PTR4), .Z(_03193__PTR5) );
  XOR2_X1 U15086 ( .A(_02979__PTR6), .B(_03192__PTR5), .Z(_03193__PTR6) );
  XOR2_X1 U15087 ( .A(_02979__PTR7), .B(_03192__PTR6), .Z(_03193__PTR7) );
  XOR2_X1 U15088 ( .A(_02979__PTR8), .B(_03192__PTR7), .Z(_03193__PTR8) );
  XOR2_X1 U15089 ( .A(_02979__PTR9), .B(_03192__PTR8), .Z(_03193__PTR9) );
  XOR2_X1 U15090 ( .A(_02979__PTR10), .B(_03192__PTR9), .Z(_03193__PTR10) );
  XOR2_X1 U15091 ( .A(_02979__PTR11), .B(_03192__PTR10), .Z(_03193__PTR11) );
  XOR2_X1 U15092 ( .A(_02979__PTR12), .B(_03192__PTR11), .Z(_03193__PTR12) );
  XOR2_X1 U15093 ( .A(_02979__PTR13), .B(_03192__PTR12), .Z(_03193__PTR13) );
  XOR2_X1 U15094 ( .A(_02979__PTR14), .B(_03192__PTR13), .Z(_03193__PTR14) );
  XOR2_X1 U15095 ( .A(_02979__PTR15), .B(_03192__PTR14), .Z(_03193__PTR15) );
  XOR2_X1 U15096 ( .A(_02979__PTR16), .B(_03192__PTR15), .Z(_03193__PTR16) );
  XOR2_X1 U15097 ( .A(_02979__PTR17), .B(_03192__PTR16), .Z(_03193__PTR17) );
  XOR2_X1 U15098 ( .A(_02979__PTR18), .B(_03192__PTR17), .Z(_03193__PTR18) );
  XOR2_X1 U15099 ( .A(_02979__PTR19), .B(_03192__PTR18), .Z(_03193__PTR19) );
  XOR2_X1 U15100 ( .A(_02979__PTR20), .B(_03192__PTR19), .Z(_03193__PTR20) );
  XOR2_X1 U15101 ( .A(_02979__PTR21), .B(_03192__PTR20), .Z(_03193__PTR21) );
  XOR2_X1 U15102 ( .A(_02979__PTR22), .B(_03192__PTR21), .Z(_03193__PTR22) );
  XOR2_X1 U15103 ( .A(_02979__PTR23), .B(_03192__PTR22), .Z(_03193__PTR23) );
  XOR2_X1 U15104 ( .A(_02979__PTR24), .B(_03192__PTR23), .Z(_03193__PTR24) );
  XOR2_X1 U15105 ( .A(_02979__PTR25), .B(_03192__PTR24), .Z(_03193__PTR25) );
  XOR2_X1 U15106 ( .A(_02979__PTR26), .B(_03192__PTR25), .Z(_03193__PTR26) );
  XOR2_X1 U15107 ( .A(_02979__PTR27), .B(_03192__PTR26), .Z(_03193__PTR27) );
  XOR2_X1 U15108 ( .A(_02979__PTR28), .B(_03192__PTR27), .Z(_03193__PTR28) );
  XOR2_X1 U15109 ( .A(_02979__PTR29), .B(_03192__PTR28), .Z(_03193__PTR29) );
  XOR2_X1 U15110 ( .A(_02979__PTR30), .B(_03192__PTR29), .Z(_03193__PTR30) );
  XOR2_X1 U15111 ( .A(_02977__PTR31), .B(_03192__PTR30), .Z(_03193__PTR31) );
  XOR2_X1 U15112 ( .A(_03177__PTR1), .B(_03176__PTR0), .Z(_02962__PTR1) );
  XOR2_X1 U15113 ( .A(_03177__PTR2), .B(_03176__PTR1), .Z(_02962__PTR2) );
  XOR2_X1 U15114 ( .A(_03177__PTR3), .B(_03176__PTR2), .Z(_02962__PTR3) );
  XOR2_X1 U15115 ( .A(_03177__PTR4), .B(_03176__PTR3), .Z(_02962__PTR4) );
  XOR2_X1 U15116 ( .A(P2_P1_InstQueueWr_Addr_PTR0), .B(_02176__PTR3), .Z(_02963__PTR0) );
  XOR2_X1 U15117 ( .A(P2_P1_InstQueueWr_Addr_PTR1), .B(_02182__PTR4), .Z(_03177__PTR1) );
  XOR2_X1 U15118 ( .A(P2_P1_InstQueueWr_Addr_PTR2), .B(_02178__PTR5), .Z(_03177__PTR2) );
  XOR2_X1 U15119 ( .A(P2_P1_InstQueueWr_Addr_PTR3), .B(_03175__PTR3), .Z(_03177__PTR3) );
  XOR2_X1 U15120 ( .A(P2_P1_InstQueueWr_Addr_PTR4), .B(_02996__PTR4), .Z(_03177__PTR4) );
  AND2_X1 U15121 ( .A1(P2_P1_InstQueueWr_Addr_PTR0), .A2(_02176__PTR3), .ZN(_03178__PTR0) );
  AND2_X1 U15122 ( .A1(P2_P1_InstQueueWr_Addr_PTR1), .A2(_02182__PTR4), .ZN(_03178__PTR1) );
  AND2_X1 U15123 ( .A1(P2_P1_InstQueueWr_Addr_PTR2), .A2(_02178__PTR5), .ZN(_03178__PTR2) );
  AND2_X1 U15124 ( .A1(P2_P1_InstQueueWr_Addr_PTR3), .A2(_03175__PTR3), .ZN(_03178__PTR3) );
  AND2_X1 U15125 ( .A1(P2_P1_InstQueueWr_Addr_PTR4), .A2(_02996__PTR4), .ZN(_03178__PTR4) );
  XOR2_X1 U15126 ( .A(_02178__PTR5), .B(_02995__PTR1), .Z(_03065__PTR2) );
  XOR2_X1 U15127 ( .A(P2_P1_InstQueueRd_Addr_PTR3), .B(_03064__PTR2), .Z(_03065__PTR3) );
  XOR2_X1 U15128 ( .A(P2_P1_InstQueueRd_Addr_PTR2), .B(P2_P1_InstQueueRd_Addr_PTR1), .Z(_02182__PTR5) );
  XOR2_X1 U15129 ( .A(P2_P1_InstQueueRd_Addr_PTR3), .B(_03062__PTR1), .Z(_02182__PTR6) );
  XOR2_X1 U15130 ( .A(P2_P1_InstQueueRd_Addr_PTR4), .B(_03062__PTR2), .Z(_03063__PTR3) );
  XOR2_X1 U15131 ( .A(_02179__PTR1), .B(_03059__PTR0), .Z(_03061__PTR1) );
  XOR2_X1 U15132 ( .A(_02179__PTR2), .B(_03059__PTR1), .Z(_03061__PTR2) );
  XOR2_X1 U15133 ( .A(_02179__PTR3), .B(_03059__PTR2), .Z(_03061__PTR3) );
  XOR2_X1 U15134 ( .A(_02179__PTR4), .B(_03059__PTR3), .Z(_03061__PTR4) );
  XOR2_X1 U15135 ( .A(_02179__PTR5), .B(_03059__PTR4), .Z(_03061__PTR5) );
  XOR2_X1 U15136 ( .A(_02179__PTR6), .B(_03059__PTR5), .Z(_03061__PTR6) );
  XOR2_X1 U15137 ( .A(_02179__PTR7), .B(_03059__PTR6), .Z(_03061__PTR7) );
  XOR2_X1 U15138 ( .A(_02179__PTR0), .B(_02181__PTR7), .Z(_03060__PTR0) );
  AND2_X1 U15139 ( .A1(_02179__PTR0), .A2(_02181__PTR7), .ZN(_03059__PTR0) );
  XOR2_X1 U15140 ( .A(_02182__PTR4), .B(P2_P1_InstQueueRd_Addr_PTR0), .Z(_02180__PTR4) );
  XOR2_X1 U15141 ( .A(P2_P1_InstQueueRd_Addr_PTR2), .B(_03058__PTR1), .Z(_02180__PTR5) );
  XOR2_X1 U15142 ( .A(P2_P1_InstQueueRd_Addr_PTR3), .B(_03058__PTR2), .Z(_02180__PTR6) );
  XOR2_X1 U15143 ( .A(P2_P1_InstQueueRd_Addr_PTR3), .B(P2_P1_InstQueueRd_Addr_PTR2), .Z(_02178__PTR6) );
  XOR2_X1 U15144 ( .A(P2_P1_InstAddrPointer_PTR1), .B(P2_P1_InstAddrPointer_PTR0), .Z(_02373__PTR1) );
  XOR2_X1 U15145 ( .A(_02990__PTR2), .B(_03043__PTR1), .Z(_03052__PTR2) );
  XOR2_X1 U15146 ( .A(P2_P1_InstAddrPointer_PTR3), .B(_03051__PTR2), .Z(_03052__PTR3) );
  XOR2_X1 U15147 ( .A(P2_P1_InstAddrPointer_PTR4), .B(_03051__PTR3), .Z(_03052__PTR4) );
  XOR2_X1 U15148 ( .A(P2_P1_InstAddrPointer_PTR5), .B(_03051__PTR4), .Z(_03052__PTR5) );
  XOR2_X1 U15149 ( .A(P2_P1_InstAddrPointer_PTR6), .B(_03051__PTR5), .Z(_03052__PTR6) );
  XOR2_X1 U15150 ( .A(P2_P1_InstAddrPointer_PTR7), .B(_03051__PTR6), .Z(_03052__PTR7) );
  XOR2_X1 U15151 ( .A(P2_P1_InstAddrPointer_PTR8), .B(_03051__PTR7), .Z(_03052__PTR8) );
  XOR2_X1 U15152 ( .A(P2_P1_InstAddrPointer_PTR9), .B(_03051__PTR8), .Z(_03052__PTR9) );
  XOR2_X1 U15153 ( .A(P2_P1_InstAddrPointer_PTR10), .B(_03051__PTR9), .Z(_03052__PTR10) );
  XOR2_X1 U15154 ( .A(P2_P1_InstAddrPointer_PTR11), .B(_03051__PTR10), .Z(_03052__PTR11) );
  XOR2_X1 U15155 ( .A(P2_P1_InstAddrPointer_PTR12), .B(_03051__PTR11), .Z(_03052__PTR12) );
  XOR2_X1 U15156 ( .A(P2_P1_InstAddrPointer_PTR13), .B(_03051__PTR12), .Z(_03052__PTR13) );
  XOR2_X1 U15157 ( .A(P2_P1_InstAddrPointer_PTR14), .B(_03051__PTR13), .Z(_03052__PTR14) );
  XOR2_X1 U15158 ( .A(P2_P1_InstAddrPointer_PTR15), .B(_03051__PTR14), .Z(_03052__PTR15) );
  XOR2_X1 U15159 ( .A(P2_P1_InstAddrPointer_PTR16), .B(_03051__PTR15), .Z(_03052__PTR16) );
  XOR2_X1 U15160 ( .A(P2_P1_InstAddrPointer_PTR17), .B(_03051__PTR16), .Z(_03052__PTR17) );
  XOR2_X1 U15161 ( .A(P2_P1_InstAddrPointer_PTR18), .B(_03051__PTR17), .Z(_03052__PTR18) );
  XOR2_X1 U15162 ( .A(P2_P1_InstAddrPointer_PTR19), .B(_03051__PTR18), .Z(_03052__PTR19) );
  XOR2_X1 U15163 ( .A(P2_P1_InstAddrPointer_PTR20), .B(_03051__PTR19), .Z(_03052__PTR20) );
  XOR2_X1 U15164 ( .A(P2_P1_InstAddrPointer_PTR21), .B(_03051__PTR20), .Z(_03052__PTR21) );
  XOR2_X1 U15165 ( .A(P2_P1_InstAddrPointer_PTR22), .B(_03051__PTR21), .Z(_03052__PTR22) );
  XOR2_X1 U15166 ( .A(P2_P1_InstAddrPointer_PTR23), .B(_03051__PTR22), .Z(_03052__PTR23) );
  XOR2_X1 U15167 ( .A(P2_P1_InstAddrPointer_PTR24), .B(_03051__PTR23), .Z(_03052__PTR24) );
  XOR2_X1 U15168 ( .A(P2_P1_InstAddrPointer_PTR25), .B(_03051__PTR24), .Z(_03052__PTR25) );
  XOR2_X1 U15169 ( .A(P2_P1_InstAddrPointer_PTR26), .B(_03051__PTR25), .Z(_03052__PTR26) );
  XOR2_X1 U15170 ( .A(P2_P1_InstAddrPointer_PTR27), .B(_03051__PTR26), .Z(_03052__PTR27) );
  XOR2_X1 U15171 ( .A(P2_P1_InstAddrPointer_PTR28), .B(_03051__PTR27), .Z(_03052__PTR28) );
  XOR2_X1 U15172 ( .A(P2_P1_InstAddrPointer_PTR29), .B(_03051__PTR28), .Z(_03052__PTR29) );
  XOR2_X1 U15173 ( .A(P2_P1_InstAddrPointer_PTR30), .B(_03051__PTR29), .Z(_03052__PTR30) );
  XOR2_X1 U15174 ( .A(P2_P1_InstAddrPointer_PTR31), .B(_03051__PTR30), .Z(_03052__PTR31) );
  XOR2_X1 U15175 ( .A(_03054__PTR1), .B(_03053__PTR0), .Z(_03055__PTR1) );
  XOR2_X1 U15176 ( .A(_03054__PTR2), .B(_03053__PTR1), .Z(_03055__PTR2) );
  XOR2_X1 U15177 ( .A(_03054__PTR3), .B(_03053__PTR2), .Z(_03055__PTR3) );
  XOR2_X1 U15178 ( .A(_03054__PTR4), .B(_03053__PTR3), .Z(_03055__PTR4) );
  XOR2_X1 U15179 ( .A(_03054__PTR5), .B(_03053__PTR4), .Z(_03055__PTR5) );
  XOR2_X1 U15180 ( .A(_03054__PTR6), .B(_03053__PTR5), .Z(_03055__PTR6) );
  XOR2_X1 U15181 ( .A(_03054__PTR7), .B(_03053__PTR6), .Z(_03055__PTR7) );
  XOR2_X1 U15182 ( .A(_03052__PTR8), .B(_03053__PTR7), .Z(_03055__PTR8) );
  XOR2_X1 U15183 ( .A(_03052__PTR9), .B(_03053__PTR8), .Z(_03055__PTR9) );
  XOR2_X1 U15184 ( .A(_03052__PTR10), .B(_03053__PTR9), .Z(_03055__PTR10) );
  XOR2_X1 U15185 ( .A(_03052__PTR11), .B(_03053__PTR10), .Z(_03055__PTR11) );
  XOR2_X1 U15186 ( .A(_03052__PTR12), .B(_03053__PTR11), .Z(_03055__PTR12) );
  XOR2_X1 U15187 ( .A(_03052__PTR13), .B(_03053__PTR12), .Z(_03055__PTR13) );
  XOR2_X1 U15188 ( .A(_03052__PTR14), .B(_03053__PTR13), .Z(_03055__PTR14) );
  XOR2_X1 U15189 ( .A(_03052__PTR15), .B(_03053__PTR14), .Z(_03055__PTR15) );
  XOR2_X1 U15190 ( .A(_03052__PTR16), .B(_03053__PTR15), .Z(_03055__PTR16) );
  XOR2_X1 U15191 ( .A(_03052__PTR17), .B(_03053__PTR16), .Z(_03055__PTR17) );
  XOR2_X1 U15192 ( .A(_03052__PTR18), .B(_03053__PTR17), .Z(_03055__PTR18) );
  XOR2_X1 U15193 ( .A(_03052__PTR19), .B(_03053__PTR18), .Z(_03055__PTR19) );
  XOR2_X1 U15194 ( .A(_03052__PTR20), .B(_03053__PTR19), .Z(_03055__PTR20) );
  XOR2_X1 U15195 ( .A(_03052__PTR21), .B(_03053__PTR20), .Z(_03055__PTR21) );
  XOR2_X1 U15196 ( .A(_03052__PTR22), .B(_03053__PTR21), .Z(_03055__PTR22) );
  XOR2_X1 U15197 ( .A(_03052__PTR23), .B(_03053__PTR22), .Z(_03055__PTR23) );
  XOR2_X1 U15198 ( .A(_03052__PTR24), .B(_03053__PTR23), .Z(_03055__PTR24) );
  XOR2_X1 U15199 ( .A(_03052__PTR25), .B(_03053__PTR24), .Z(_03055__PTR25) );
  XOR2_X1 U15200 ( .A(_03052__PTR26), .B(_03053__PTR25), .Z(_03055__PTR26) );
  XOR2_X1 U15201 ( .A(_03052__PTR27), .B(_03053__PTR26), .Z(_03055__PTR27) );
  XOR2_X1 U15202 ( .A(_03052__PTR28), .B(_03053__PTR27), .Z(_03055__PTR28) );
  XOR2_X1 U15203 ( .A(_03052__PTR29), .B(_03053__PTR28), .Z(_03055__PTR29) );
  XOR2_X1 U15204 ( .A(_03052__PTR30), .B(_03053__PTR29), .Z(_03055__PTR30) );
  XOR2_X1 U15205 ( .A(_03052__PTR31), .B(_03053__PTR30), .Z(_03055__PTR31) );
  XOR2_X1 U15206 ( .A(_02373__PTR0), .B(_02177__PTR0), .Z(_03054__PTR0) );
  XOR2_X1 U15207 ( .A(_03052__PTR2), .B(_02177__PTR2), .Z(_03054__PTR2) );
  XOR2_X1 U15208 ( .A(_03052__PTR3), .B(_02177__PTR3), .Z(_03054__PTR3) );
  XOR2_X1 U15209 ( .A(_03052__PTR4), .B(_02177__PTR4), .Z(_03054__PTR4) );
  XOR2_X1 U15210 ( .A(_03052__PTR5), .B(_02177__PTR5), .Z(_03054__PTR5) );
  XOR2_X1 U15211 ( .A(_03052__PTR6), .B(_02177__PTR6), .Z(_03054__PTR6) );
  XOR2_X1 U15212 ( .A(_03052__PTR7), .B(_02177__PTR7), .Z(_03054__PTR7) );
  AND2_X1 U15213 ( .A1(_02373__PTR0), .A2(_02177__PTR0), .ZN(_03053__PTR0) );
  AND2_X1 U15214 ( .A1(_02373__PTR1), .A2(_02177__PTR1), .ZN(_03056__PTR1) );
  AND2_X1 U15215 ( .A1(_03052__PTR2), .A2(_02177__PTR2), .ZN(_03056__PTR2) );
  AND2_X1 U15216 ( .A1(_03052__PTR3), .A2(_02177__PTR3), .ZN(_03056__PTR3) );
  AND2_X1 U15217 ( .A1(_03052__PTR4), .A2(_02177__PTR4), .ZN(_03056__PTR4) );
  AND2_X1 U15218 ( .A1(_03052__PTR5), .A2(_02177__PTR5), .ZN(_03056__PTR5) );
  AND2_X1 U15219 ( .A1(_03052__PTR6), .A2(_02177__PTR6), .ZN(_03056__PTR6) );
  AND2_X1 U15220 ( .A1(_03052__PTR7), .A2(_02177__PTR7), .ZN(_03056__PTR7) );
  XOR2_X1 U15221 ( .A(P2_P1_InstAddrPointer_PTR2), .B(P2_P1_InstAddrPointer_PTR1), .Z(_02373__PTR34) );
  XOR2_X1 U15222 ( .A(P2_P1_InstAddrPointer_PTR3), .B(_03046__PTR1), .Z(_02373__PTR35) );
  XOR2_X1 U15223 ( .A(P2_P1_InstAddrPointer_PTR4), .B(_03046__PTR2), .Z(_02373__PTR36) );
  XOR2_X1 U15224 ( .A(P2_P1_InstAddrPointer_PTR5), .B(_03046__PTR3), .Z(_02373__PTR37) );
  XOR2_X1 U15225 ( .A(P2_P1_InstAddrPointer_PTR6), .B(_03046__PTR4), .Z(_02373__PTR38) );
  XOR2_X1 U15226 ( .A(P2_P1_InstAddrPointer_PTR7), .B(_03046__PTR5), .Z(_02373__PTR39) );
  XOR2_X1 U15227 ( .A(P2_P1_InstAddrPointer_PTR8), .B(_03046__PTR6), .Z(_02373__PTR40) );
  XOR2_X1 U15228 ( .A(P2_P1_InstAddrPointer_PTR9), .B(_03046__PTR7), .Z(_02373__PTR41) );
  XOR2_X1 U15229 ( .A(P2_P1_InstAddrPointer_PTR10), .B(_03046__PTR8), .Z(_02373__PTR42) );
  XOR2_X1 U15230 ( .A(P2_P1_InstAddrPointer_PTR11), .B(_03046__PTR9), .Z(_02373__PTR43) );
  XOR2_X1 U15231 ( .A(P2_P1_InstAddrPointer_PTR12), .B(_03046__PTR10), .Z(_02373__PTR44) );
  XOR2_X1 U15232 ( .A(P2_P1_InstAddrPointer_PTR13), .B(_03046__PTR11), .Z(_02373__PTR45) );
  XOR2_X1 U15233 ( .A(P2_P1_InstAddrPointer_PTR14), .B(_03046__PTR12), .Z(_02373__PTR46) );
  XOR2_X1 U15234 ( .A(P2_P1_InstAddrPointer_PTR15), .B(_03046__PTR13), .Z(_02373__PTR47) );
  XOR2_X1 U15235 ( .A(P2_P1_InstAddrPointer_PTR16), .B(_03046__PTR14), .Z(_02373__PTR48) );
  XOR2_X1 U15236 ( .A(P2_P1_InstAddrPointer_PTR17), .B(_03046__PTR15), .Z(_02373__PTR49) );
  XOR2_X1 U15237 ( .A(P2_P1_InstAddrPointer_PTR18), .B(_03046__PTR16), .Z(_02373__PTR50) );
  XOR2_X1 U15238 ( .A(P2_P1_InstAddrPointer_PTR19), .B(_03046__PTR17), .Z(_02373__PTR51) );
  XOR2_X1 U15239 ( .A(P2_P1_InstAddrPointer_PTR20), .B(_03046__PTR18), .Z(_02373__PTR52) );
  XOR2_X1 U15240 ( .A(P2_P1_InstAddrPointer_PTR21), .B(_03046__PTR19), .Z(_02373__PTR53) );
  XOR2_X1 U15241 ( .A(P2_P1_InstAddrPointer_PTR22), .B(_03046__PTR20), .Z(_02373__PTR54) );
  XOR2_X1 U15242 ( .A(P2_P1_InstAddrPointer_PTR23), .B(_03046__PTR21), .Z(_02373__PTR55) );
  XOR2_X1 U15243 ( .A(P2_P1_InstAddrPointer_PTR24), .B(_03046__PTR22), .Z(_02373__PTR56) );
  XOR2_X1 U15244 ( .A(P2_P1_InstAddrPointer_PTR25), .B(_03046__PTR23), .Z(_02373__PTR57) );
  XOR2_X1 U15245 ( .A(P2_P1_InstAddrPointer_PTR26), .B(_03046__PTR24), .Z(_02373__PTR58) );
  XOR2_X1 U15246 ( .A(P2_P1_InstAddrPointer_PTR27), .B(_03046__PTR25), .Z(_02373__PTR59) );
  XOR2_X1 U15247 ( .A(P2_P1_InstAddrPointer_PTR28), .B(_03046__PTR26), .Z(_02373__PTR60) );
  XOR2_X1 U15248 ( .A(P2_P1_InstAddrPointer_PTR29), .B(_03046__PTR27), .Z(_02373__PTR61) );
  XOR2_X1 U15249 ( .A(P2_P1_InstAddrPointer_PTR30), .B(_03046__PTR28), .Z(_02373__PTR62) );
  XOR2_X1 U15250 ( .A(P2_P1_InstAddrPointer_PTR31), .B(_03046__PTR29), .Z(_02373__PTR63) );
  XOR2_X1 U15251 ( .A(_03048__PTR1), .B(_03047__PTR0), .Z(_03049__PTR1) );
  XOR2_X1 U15252 ( .A(_03048__PTR2), .B(_03047__PTR1), .Z(_03049__PTR2) );
  XOR2_X1 U15253 ( .A(_03048__PTR3), .B(_03047__PTR2), .Z(_03049__PTR3) );
  XOR2_X1 U15254 ( .A(_03048__PTR4), .B(_03047__PTR3), .Z(_03049__PTR4) );
  XOR2_X1 U15255 ( .A(_03048__PTR5), .B(_03047__PTR4), .Z(_03049__PTR5) );
  XOR2_X1 U15256 ( .A(_03048__PTR6), .B(_03047__PTR5), .Z(_03049__PTR6) );
  XOR2_X1 U15257 ( .A(_03048__PTR7), .B(_03047__PTR6), .Z(_03049__PTR7) );
  XOR2_X1 U15258 ( .A(_02373__PTR40), .B(_03047__PTR7), .Z(_03049__PTR8) );
  XOR2_X1 U15259 ( .A(_02373__PTR41), .B(_03047__PTR8), .Z(_03049__PTR9) );
  XOR2_X1 U15260 ( .A(_02373__PTR42), .B(_03047__PTR9), .Z(_03049__PTR10) );
  XOR2_X1 U15261 ( .A(_02373__PTR43), .B(_03047__PTR10), .Z(_03049__PTR11) );
  XOR2_X1 U15262 ( .A(_02373__PTR44), .B(_03047__PTR11), .Z(_03049__PTR12) );
  XOR2_X1 U15263 ( .A(_02373__PTR45), .B(_03047__PTR12), .Z(_03049__PTR13) );
  XOR2_X1 U15264 ( .A(_02373__PTR46), .B(_03047__PTR13), .Z(_03049__PTR14) );
  XOR2_X1 U15265 ( .A(_02373__PTR47), .B(_03047__PTR14), .Z(_03049__PTR15) );
  XOR2_X1 U15266 ( .A(_02373__PTR48), .B(_03047__PTR15), .Z(_03049__PTR16) );
  XOR2_X1 U15267 ( .A(_02373__PTR49), .B(_03047__PTR16), .Z(_03049__PTR17) );
  XOR2_X1 U15268 ( .A(_02373__PTR50), .B(_03047__PTR17), .Z(_03049__PTR18) );
  XOR2_X1 U15269 ( .A(_02373__PTR51), .B(_03047__PTR18), .Z(_03049__PTR19) );
  XOR2_X1 U15270 ( .A(_02373__PTR52), .B(_03047__PTR19), .Z(_03049__PTR20) );
  XOR2_X1 U15271 ( .A(_02373__PTR53), .B(_03047__PTR20), .Z(_03049__PTR21) );
  XOR2_X1 U15272 ( .A(_02373__PTR54), .B(_03047__PTR21), .Z(_03049__PTR22) );
  XOR2_X1 U15273 ( .A(_02373__PTR55), .B(_03047__PTR22), .Z(_03049__PTR23) );
  XOR2_X1 U15274 ( .A(_02373__PTR56), .B(_03047__PTR23), .Z(_03049__PTR24) );
  XOR2_X1 U15275 ( .A(_02373__PTR57), .B(_03047__PTR24), .Z(_03049__PTR25) );
  XOR2_X1 U15276 ( .A(_02373__PTR58), .B(_03047__PTR25), .Z(_03049__PTR26) );
  XOR2_X1 U15277 ( .A(_02373__PTR59), .B(_03047__PTR26), .Z(_03049__PTR27) );
  XOR2_X1 U15278 ( .A(_02373__PTR60), .B(_03047__PTR27), .Z(_03049__PTR28) );
  XOR2_X1 U15279 ( .A(_02373__PTR61), .B(_03047__PTR28), .Z(_03049__PTR29) );
  XOR2_X1 U15280 ( .A(_02373__PTR62), .B(_03047__PTR29), .Z(_03049__PTR30) );
  XOR2_X1 U15281 ( .A(_02373__PTR63), .B(_03047__PTR30), .Z(_03049__PTR31) );
  XOR2_X1 U15282 ( .A(P2_P1_InstAddrPointer_PTR0), .B(_02177__PTR0), .Z(_03048__PTR0) );
  XOR2_X1 U15283 ( .A(_02373__PTR33), .B(_02177__PTR1), .Z(_03048__PTR1) );
  XOR2_X1 U15284 ( .A(_02373__PTR34), .B(_02177__PTR2), .Z(_03048__PTR2) );
  XOR2_X1 U15285 ( .A(_02373__PTR35), .B(_02177__PTR3), .Z(_03048__PTR3) );
  XOR2_X1 U15286 ( .A(_02373__PTR36), .B(_02177__PTR4), .Z(_03048__PTR4) );
  XOR2_X1 U15287 ( .A(_02373__PTR37), .B(_02177__PTR5), .Z(_03048__PTR5) );
  XOR2_X1 U15288 ( .A(_02373__PTR38), .B(_02177__PTR6), .Z(_03048__PTR6) );
  XOR2_X1 U15289 ( .A(_02373__PTR39), .B(_02177__PTR7), .Z(_03048__PTR7) );
  AND2_X1 U15290 ( .A1(P2_P1_InstAddrPointer_PTR0), .A2(_02177__PTR0), .ZN(_03047__PTR0) );
  AND2_X1 U15291 ( .A1(_02373__PTR33), .A2(_02177__PTR1), .ZN(_03050__PTR1) );
  AND2_X1 U15292 ( .A1(_02373__PTR34), .A2(_02177__PTR2), .ZN(_03050__PTR2) );
  AND2_X1 U15293 ( .A1(_02373__PTR35), .A2(_02177__PTR3), .ZN(_03050__PTR3) );
  AND2_X1 U15294 ( .A1(_02373__PTR36), .A2(_02177__PTR4), .ZN(_03050__PTR4) );
  AND2_X1 U15295 ( .A1(_02373__PTR37), .A2(_02177__PTR5), .ZN(_03050__PTR5) );
  AND2_X1 U15296 ( .A1(_02373__PTR38), .A2(_02177__PTR6), .ZN(_03050__PTR6) );
  AND2_X1 U15297 ( .A1(_02373__PTR39), .A2(_02177__PTR7), .ZN(_03050__PTR7) );
  XOR2_X1 U15298 ( .A(_02177__PTR5), .B(_02969__PTR4), .Z(_02970__PTR5) );
  XOR2_X1 U15299 ( .A(_02177__PTR6), .B(_02969__PTR5), .Z(_02970__PTR6) );
  XOR2_X1 U15300 ( .A(_02177__PTR7), .B(_02969__PTR6), .Z(_03180__PTR7) );
  XOR2_X1 U15301 ( .A(P2_P1_InstAddrPointer_PTR2), .B(_03043__PTR1), .Z(_02373__PTR2) );
  XOR2_X1 U15302 ( .A(P2_P1_InstAddrPointer_PTR3), .B(_03043__PTR2), .Z(_02373__PTR3) );
  XOR2_X1 U15303 ( .A(P2_P1_InstAddrPointer_PTR4), .B(_03043__PTR3), .Z(_02373__PTR4) );
  XOR2_X1 U15304 ( .A(P2_P1_InstAddrPointer_PTR5), .B(_03043__PTR4), .Z(_02373__PTR5) );
  XOR2_X1 U15305 ( .A(P2_P1_InstAddrPointer_PTR6), .B(_03043__PTR5), .Z(_02373__PTR6) );
  XOR2_X1 U15306 ( .A(P2_P1_InstAddrPointer_PTR7), .B(_03043__PTR6), .Z(_02373__PTR7) );
  XOR2_X1 U15307 ( .A(P2_P1_InstAddrPointer_PTR8), .B(_03043__PTR7), .Z(_02373__PTR8) );
  XOR2_X1 U15308 ( .A(P2_P1_InstAddrPointer_PTR9), .B(_03043__PTR8), .Z(_02373__PTR9) );
  XOR2_X1 U15309 ( .A(P2_P1_InstAddrPointer_PTR10), .B(_03043__PTR9), .Z(_02373__PTR10) );
  XOR2_X1 U15310 ( .A(P2_P1_InstAddrPointer_PTR11), .B(_03043__PTR10), .Z(_02373__PTR11) );
  XOR2_X1 U15311 ( .A(P2_P1_InstAddrPointer_PTR12), .B(_03043__PTR11), .Z(_02373__PTR12) );
  XOR2_X1 U15312 ( .A(P2_P1_InstAddrPointer_PTR13), .B(_03043__PTR12), .Z(_02373__PTR13) );
  XOR2_X1 U15313 ( .A(P2_P1_InstAddrPointer_PTR14), .B(_03043__PTR13), .Z(_02373__PTR14) );
  XOR2_X1 U15314 ( .A(P2_P1_InstAddrPointer_PTR15), .B(_03043__PTR14), .Z(_02373__PTR15) );
  XOR2_X1 U15315 ( .A(P2_P1_InstAddrPointer_PTR16), .B(_03043__PTR15), .Z(_02373__PTR16) );
  XOR2_X1 U15316 ( .A(P2_P1_InstAddrPointer_PTR17), .B(_03043__PTR16), .Z(_02373__PTR17) );
  XOR2_X1 U15317 ( .A(P2_P1_InstAddrPointer_PTR18), .B(_03043__PTR17), .Z(_02373__PTR18) );
  XOR2_X1 U15318 ( .A(P2_P1_InstAddrPointer_PTR19), .B(_03043__PTR18), .Z(_02373__PTR19) );
  XOR2_X1 U15319 ( .A(P2_P1_InstAddrPointer_PTR20), .B(_03043__PTR19), .Z(_02373__PTR20) );
  XOR2_X1 U15320 ( .A(P2_P1_InstAddrPointer_PTR21), .B(_03043__PTR20), .Z(_02373__PTR21) );
  XOR2_X1 U15321 ( .A(P2_P1_InstAddrPointer_PTR22), .B(_03043__PTR21), .Z(_02373__PTR22) );
  XOR2_X1 U15322 ( .A(P2_P1_InstAddrPointer_PTR23), .B(_03043__PTR22), .Z(_02373__PTR23) );
  XOR2_X1 U15323 ( .A(P2_P1_InstAddrPointer_PTR24), .B(_03043__PTR23), .Z(_02373__PTR24) );
  XOR2_X1 U15324 ( .A(P2_P1_InstAddrPointer_PTR25), .B(_03043__PTR24), .Z(_02373__PTR25) );
  XOR2_X1 U15325 ( .A(P2_P1_InstAddrPointer_PTR26), .B(_03043__PTR25), .Z(_02373__PTR26) );
  XOR2_X1 U15326 ( .A(P2_P1_InstAddrPointer_PTR27), .B(_03043__PTR26), .Z(_02373__PTR27) );
  XOR2_X1 U15327 ( .A(P2_P1_InstAddrPointer_PTR28), .B(_03043__PTR27), .Z(_02373__PTR28) );
  XOR2_X1 U15328 ( .A(P2_P1_InstAddrPointer_PTR29), .B(_03043__PTR28), .Z(_02373__PTR29) );
  XOR2_X1 U15329 ( .A(P2_P1_InstAddrPointer_PTR30), .B(_03043__PTR29), .Z(_02373__PTR30) );
  XOR2_X1 U15330 ( .A(P2_P1_InstAddrPointer_PTR31), .B(_03043__PTR30), .Z(_02373__PTR31) );
  XOR2_X1 U15331 ( .A(_03054__PTR1), .B(_03182__PTR0), .Z(_03184__PTR1) );
  XOR2_X1 U15332 ( .A(_03183__PTR2), .B(_03182__PTR1), .Z(_03184__PTR2) );
  XOR2_X1 U15333 ( .A(_03183__PTR3), .B(_03182__PTR2), .Z(_03184__PTR3) );
  XOR2_X1 U15334 ( .A(_03183__PTR4), .B(_03182__PTR3), .Z(_03184__PTR4) );
  XOR2_X1 U15335 ( .A(_03183__PTR5), .B(_03182__PTR4), .Z(_03184__PTR5) );
  XOR2_X1 U15336 ( .A(_03183__PTR6), .B(_03182__PTR5), .Z(_03184__PTR6) );
  XOR2_X1 U15337 ( .A(_03183__PTR7), .B(_03182__PTR6), .Z(_03184__PTR7) );
  XOR2_X1 U15338 ( .A(_03183__PTR8), .B(_03182__PTR7), .Z(_03184__PTR8) );
  XOR2_X1 U15339 ( .A(_03183__PTR9), .B(_03182__PTR8), .Z(_03184__PTR9) );
  XOR2_X1 U15340 ( .A(_03183__PTR10), .B(_03182__PTR9), .Z(_03184__PTR10) );
  XOR2_X1 U15341 ( .A(_03183__PTR11), .B(_03182__PTR10), .Z(_03184__PTR11) );
  XOR2_X1 U15342 ( .A(_03183__PTR12), .B(_03182__PTR11), .Z(_03184__PTR12) );
  XOR2_X1 U15343 ( .A(_03183__PTR13), .B(_03182__PTR12), .Z(_03184__PTR13) );
  XOR2_X1 U15344 ( .A(_03183__PTR14), .B(_03182__PTR13), .Z(_03184__PTR14) );
  XOR2_X1 U15345 ( .A(_03183__PTR15), .B(_03182__PTR14), .Z(_03184__PTR15) );
  XOR2_X1 U15346 ( .A(_03183__PTR16), .B(_03182__PTR15), .Z(_03184__PTR16) );
  XOR2_X1 U15347 ( .A(_03183__PTR17), .B(_03182__PTR16), .Z(_03184__PTR17) );
  XOR2_X1 U15348 ( .A(_03183__PTR18), .B(_03182__PTR17), .Z(_03184__PTR18) );
  XOR2_X1 U15349 ( .A(_03183__PTR19), .B(_03182__PTR18), .Z(_03184__PTR19) );
  XOR2_X1 U15350 ( .A(_03183__PTR20), .B(_03182__PTR19), .Z(_03184__PTR20) );
  XOR2_X1 U15351 ( .A(_03183__PTR21), .B(_03182__PTR20), .Z(_03184__PTR21) );
  XOR2_X1 U15352 ( .A(_03183__PTR22), .B(_03182__PTR21), .Z(_03184__PTR22) );
  XOR2_X1 U15353 ( .A(_03183__PTR23), .B(_03182__PTR22), .Z(_03184__PTR23) );
  XOR2_X1 U15354 ( .A(_03183__PTR24), .B(_03182__PTR23), .Z(_03184__PTR24) );
  XOR2_X1 U15355 ( .A(_03183__PTR25), .B(_03182__PTR24), .Z(_03184__PTR25) );
  XOR2_X1 U15356 ( .A(_03183__PTR26), .B(_03182__PTR25), .Z(_03184__PTR26) );
  XOR2_X1 U15357 ( .A(_03183__PTR27), .B(_03182__PTR26), .Z(_03184__PTR27) );
  XOR2_X1 U15358 ( .A(_03183__PTR28), .B(_03182__PTR27), .Z(_03184__PTR28) );
  XOR2_X1 U15359 ( .A(_03183__PTR29), .B(_03182__PTR28), .Z(_03184__PTR29) );
  XOR2_X1 U15360 ( .A(_03183__PTR30), .B(_03182__PTR29), .Z(_03184__PTR30) );
  XOR2_X1 U15361 ( .A(_03183__PTR32), .B(_03182__PTR30), .Z(_03184__PTR31) );
  XOR2_X1 U15362 ( .A(_02373__PTR1), .B(_02177__PTR1), .Z(_03054__PTR1) );
  XOR2_X1 U15363 ( .A(_02373__PTR2), .B(_02177__PTR2), .Z(_03183__PTR2) );
  XOR2_X1 U15364 ( .A(_02373__PTR3), .B(_02177__PTR3), .Z(_03183__PTR3) );
  XOR2_X1 U15365 ( .A(_02373__PTR4), .B(_03181__PTR4), .Z(_03183__PTR4) );
  XOR2_X1 U15366 ( .A(_02373__PTR5), .B(_03181__PTR5), .Z(_03183__PTR5) );
  XOR2_X1 U15367 ( .A(_02373__PTR6), .B(_03181__PTR6), .Z(_03183__PTR6) );
  XOR2_X1 U15368 ( .A(_02373__PTR7), .B(_03181__PTR7), .Z(_03183__PTR7) );
  XOR2_X1 U15369 ( .A(_02373__PTR8), .B(_03179__PTR8), .Z(_03183__PTR8) );
  XOR2_X1 U15370 ( .A(_02373__PTR9), .B(_03179__PTR8), .Z(_03183__PTR9) );
  XOR2_X1 U15371 ( .A(_02373__PTR10), .B(_03179__PTR8), .Z(_03183__PTR10) );
  XOR2_X1 U15372 ( .A(_02373__PTR11), .B(_03179__PTR8), .Z(_03183__PTR11) );
  XOR2_X1 U15373 ( .A(_02373__PTR12), .B(_03179__PTR8), .Z(_03183__PTR12) );
  XOR2_X1 U15374 ( .A(_02373__PTR13), .B(_03179__PTR8), .Z(_03183__PTR13) );
  XOR2_X1 U15375 ( .A(_02373__PTR14), .B(_03179__PTR8), .Z(_03183__PTR14) );
  XOR2_X1 U15376 ( .A(_02373__PTR15), .B(_03179__PTR8), .Z(_03183__PTR15) );
  XOR2_X1 U15377 ( .A(_02373__PTR16), .B(_03179__PTR8), .Z(_03183__PTR16) );
  XOR2_X1 U15378 ( .A(_02373__PTR17), .B(_03179__PTR8), .Z(_03183__PTR17) );
  XOR2_X1 U15379 ( .A(_02373__PTR18), .B(_03179__PTR8), .Z(_03183__PTR18) );
  XOR2_X1 U15380 ( .A(_02373__PTR19), .B(_03179__PTR8), .Z(_03183__PTR19) );
  XOR2_X1 U15381 ( .A(_02373__PTR20), .B(_03179__PTR8), .Z(_03183__PTR20) );
  XOR2_X1 U15382 ( .A(_02373__PTR21), .B(_03179__PTR8), .Z(_03183__PTR21) );
  XOR2_X1 U15383 ( .A(_02373__PTR22), .B(_03179__PTR8), .Z(_03183__PTR22) );
  XOR2_X1 U15384 ( .A(_02373__PTR23), .B(_03179__PTR8), .Z(_03183__PTR23) );
  XOR2_X1 U15385 ( .A(_02373__PTR24), .B(_03179__PTR8), .Z(_03183__PTR24) );
  XOR2_X1 U15386 ( .A(_02373__PTR25), .B(_03179__PTR8), .Z(_03183__PTR25) );
  XOR2_X1 U15387 ( .A(_02373__PTR26), .B(_03179__PTR8), .Z(_03183__PTR26) );
  XOR2_X1 U15388 ( .A(_02373__PTR27), .B(_03179__PTR8), .Z(_03183__PTR27) );
  XOR2_X1 U15389 ( .A(_02373__PTR28), .B(_03179__PTR8), .Z(_03183__PTR28) );
  XOR2_X1 U15390 ( .A(_02373__PTR29), .B(_03179__PTR8), .Z(_03183__PTR29) );
  XOR2_X1 U15391 ( .A(_02373__PTR30), .B(_03179__PTR8), .Z(_03183__PTR30) );
  XOR2_X1 U15392 ( .A(_02373__PTR31), .B(_03179__PTR8), .Z(_03183__PTR32) );
  AND2_X1 U15393 ( .A1(_02373__PTR2), .A2(_02177__PTR2), .ZN(_03185__PTR2) );
  AND2_X1 U15394 ( .A1(_02373__PTR3), .A2(_02177__PTR3), .ZN(_03185__PTR3) );
  AND2_X1 U15395 ( .A1(_02373__PTR4), .A2(_03181__PTR4), .ZN(_03185__PTR4) );
  AND2_X1 U15396 ( .A1(_02373__PTR5), .A2(_03181__PTR5), .ZN(_03185__PTR5) );
  AND2_X1 U15397 ( .A1(_02373__PTR6), .A2(_03181__PTR6), .ZN(_03185__PTR6) );
  AND2_X1 U15398 ( .A1(_02373__PTR7), .A2(_03181__PTR7), .ZN(_03185__PTR7) );
  AND2_X1 U15399 ( .A1(_02373__PTR8), .A2(_03179__PTR8), .ZN(_03185__PTR8) );
  AND2_X1 U15400 ( .A1(_02373__PTR9), .A2(_03179__PTR8), .ZN(_03185__PTR9) );
  AND2_X1 U15401 ( .A1(_02373__PTR10), .A2(_03179__PTR8), .ZN(_03185__PTR10) );
  AND2_X1 U15402 ( .A1(_02373__PTR11), .A2(_03179__PTR8), .ZN(_03185__PTR11) );
  AND2_X1 U15403 ( .A1(_02373__PTR12), .A2(_03179__PTR8), .ZN(_03185__PTR12) );
  AND2_X1 U15404 ( .A1(_02373__PTR13), .A2(_03179__PTR8), .ZN(_03185__PTR13) );
  AND2_X1 U15405 ( .A1(_02373__PTR14), .A2(_03179__PTR8), .ZN(_03185__PTR14) );
  AND2_X1 U15406 ( .A1(_02373__PTR15), .A2(_03179__PTR8), .ZN(_03185__PTR15) );
  AND2_X1 U15407 ( .A1(_02373__PTR16), .A2(_03179__PTR8), .ZN(_03185__PTR16) );
  AND2_X1 U15408 ( .A1(_02373__PTR17), .A2(_03179__PTR8), .ZN(_03185__PTR17) );
  AND2_X1 U15409 ( .A1(_02373__PTR18), .A2(_03179__PTR8), .ZN(_03185__PTR18) );
  AND2_X1 U15410 ( .A1(_02373__PTR19), .A2(_03179__PTR8), .ZN(_03185__PTR19) );
  AND2_X1 U15411 ( .A1(_02373__PTR20), .A2(_03179__PTR8), .ZN(_03185__PTR20) );
  AND2_X1 U15412 ( .A1(_02373__PTR21), .A2(_03179__PTR8), .ZN(_03185__PTR21) );
  AND2_X1 U15413 ( .A1(_02373__PTR22), .A2(_03179__PTR8), .ZN(_03185__PTR22) );
  AND2_X1 U15414 ( .A1(_02373__PTR23), .A2(_03179__PTR8), .ZN(_03185__PTR23) );
  AND2_X1 U15415 ( .A1(_02373__PTR24), .A2(_03179__PTR8), .ZN(_03185__PTR24) );
  AND2_X1 U15416 ( .A1(_02373__PTR25), .A2(_03179__PTR8), .ZN(_03185__PTR25) );
  AND2_X1 U15417 ( .A1(_02373__PTR26), .A2(_03179__PTR8), .ZN(_03185__PTR26) );
  AND2_X1 U15418 ( .A1(_02373__PTR27), .A2(_03179__PTR8), .ZN(_03185__PTR27) );
  AND2_X1 U15419 ( .A1(_02373__PTR28), .A2(_03179__PTR8), .ZN(_03185__PTR28) );
  AND2_X1 U15420 ( .A1(_02373__PTR29), .A2(_03179__PTR8), .ZN(_03185__PTR29) );
  AND2_X1 U15421 ( .A1(_02373__PTR30), .A2(_03179__PTR8), .ZN(_03185__PTR30) );
  XOR2_X1 U15422 ( .A(_02177__PTR4), .B(_02969__PTR3), .Z(_02970__PTR4) );
  XOR2_X1 U15423 ( .A(P2_P1_InstQueueRd_Addr_PTR2), .B(_02995__PTR1), .Z(_02176__PTR5) );
  XOR2_X1 U15424 ( .A(P2_P1_InstQueueRd_Addr_PTR3), .B(_02995__PTR2), .Z(_02176__PTR6) );
  XOR2_X1 U15425 ( .A(P2_P1_InstQueueRd_Addr_PTR4), .B(_02995__PTR3), .Z(_03045__PTR4) );
  XOR2_X1 U15426 ( .A(P2_P1_PhyAddrPointer_PTR2), .B(P2_P1_PhyAddrPointer_PTR1), .Z(_02184__PTR130) );
  XOR2_X1 U15427 ( .A(P2_P1_PhyAddrPointer_PTR3), .B(_03042__PTR1), .Z(_02184__PTR131) );
  XOR2_X1 U15428 ( .A(P2_P1_PhyAddrPointer_PTR4), .B(_03042__PTR2), .Z(_02184__PTR132) );
  XOR2_X1 U15429 ( .A(P2_P1_PhyAddrPointer_PTR5), .B(_03042__PTR3), .Z(_02184__PTR133) );
  XOR2_X1 U15430 ( .A(P2_P1_PhyAddrPointer_PTR6), .B(_03042__PTR4), .Z(_02184__PTR134) );
  XOR2_X1 U15431 ( .A(P2_P1_PhyAddrPointer_PTR7), .B(_03042__PTR5), .Z(_02184__PTR135) );
  XOR2_X1 U15432 ( .A(P2_P1_PhyAddrPointer_PTR8), .B(_03042__PTR6), .Z(_02184__PTR136) );
  XOR2_X1 U15433 ( .A(P2_P1_PhyAddrPointer_PTR9), .B(_03042__PTR7), .Z(_02184__PTR137) );
  XOR2_X1 U15434 ( .A(P2_P1_PhyAddrPointer_PTR10), .B(_03042__PTR8), .Z(_02184__PTR138) );
  XOR2_X1 U15435 ( .A(P2_P1_PhyAddrPointer_PTR11), .B(_03042__PTR9), .Z(_02184__PTR139) );
  XOR2_X1 U15436 ( .A(P2_P1_PhyAddrPointer_PTR12), .B(_03042__PTR10), .Z(_02184__PTR140) );
  XOR2_X1 U15437 ( .A(P2_P1_PhyAddrPointer_PTR13), .B(_03042__PTR11), .Z(_02184__PTR141) );
  XOR2_X1 U15438 ( .A(P2_P1_PhyAddrPointer_PTR14), .B(_03042__PTR12), .Z(_02184__PTR142) );
  XOR2_X1 U15439 ( .A(P2_P1_PhyAddrPointer_PTR15), .B(_03042__PTR13), .Z(_02184__PTR143) );
  XOR2_X1 U15440 ( .A(P2_P1_PhyAddrPointer_PTR16), .B(_03042__PTR14), .Z(_02184__PTR144) );
  XOR2_X1 U15441 ( .A(P2_P1_PhyAddrPointer_PTR17), .B(_03042__PTR15), .Z(_02184__PTR145) );
  XOR2_X1 U15442 ( .A(P2_P1_PhyAddrPointer_PTR18), .B(_03042__PTR16), .Z(_02184__PTR146) );
  XOR2_X1 U15443 ( .A(P2_P1_PhyAddrPointer_PTR19), .B(_03042__PTR17), .Z(_02184__PTR147) );
  XOR2_X1 U15444 ( .A(P2_P1_PhyAddrPointer_PTR20), .B(_03042__PTR18), .Z(_02184__PTR148) );
  XOR2_X1 U15445 ( .A(P2_P1_PhyAddrPointer_PTR21), .B(_03042__PTR19), .Z(_02184__PTR149) );
  XOR2_X1 U15446 ( .A(P2_P1_PhyAddrPointer_PTR22), .B(_03042__PTR20), .Z(_02184__PTR150) );
  XOR2_X1 U15447 ( .A(P2_P1_PhyAddrPointer_PTR23), .B(_03042__PTR21), .Z(_02184__PTR151) );
  XOR2_X1 U15448 ( .A(P2_P1_PhyAddrPointer_PTR24), .B(_03042__PTR22), .Z(_02184__PTR152) );
  XOR2_X1 U15449 ( .A(P2_P1_PhyAddrPointer_PTR25), .B(_03042__PTR23), .Z(_02184__PTR153) );
  XOR2_X1 U15450 ( .A(P2_P1_PhyAddrPointer_PTR26), .B(_03042__PTR24), .Z(_02184__PTR154) );
  XOR2_X1 U15451 ( .A(P2_P1_PhyAddrPointer_PTR27), .B(_03042__PTR25), .Z(_02184__PTR155) );
  XOR2_X1 U15452 ( .A(P2_P1_PhyAddrPointer_PTR28), .B(_03042__PTR26), .Z(_02184__PTR156) );
  XOR2_X1 U15453 ( .A(P2_P1_PhyAddrPointer_PTR29), .B(_03042__PTR27), .Z(_02184__PTR157) );
  XOR2_X1 U15454 ( .A(P2_P1_PhyAddrPointer_PTR30), .B(_03042__PTR28), .Z(_02184__PTR158) );
  XOR2_X1 U15455 ( .A(P2_P1_PhyAddrPointer_PTR31), .B(_03042__PTR29), .Z(_02184__PTR159) );
  XOR2_X1 U15456 ( .A(P2_P1_PhyAddrPointer_PTR1), .B(_02960__PTR0), .Z(_03191__PTR1) );
  XOR2_X1 U15457 ( .A(_02960__PTR2), .B(_03190__PTR1), .Z(_03191__PTR2) );
  XOR2_X1 U15458 ( .A(_02960__PTR3), .B(_03190__PTR2), .Z(_03191__PTR3) );
  XOR2_X1 U15459 ( .A(_02960__PTR4), .B(_03190__PTR3), .Z(_03191__PTR4) );
  XOR2_X1 U15460 ( .A(_02960__PTR5), .B(_03190__PTR4), .Z(_03191__PTR5) );
  XOR2_X1 U15461 ( .A(_02960__PTR6), .B(_03190__PTR5), .Z(_03191__PTR6) );
  XOR2_X1 U15462 ( .A(_02960__PTR7), .B(_03190__PTR6), .Z(_03191__PTR7) );
  XOR2_X1 U15463 ( .A(_02960__PTR8), .B(_03190__PTR7), .Z(_03191__PTR8) );
  XOR2_X1 U15464 ( .A(_02960__PTR9), .B(_03190__PTR8), .Z(_03191__PTR9) );
  XOR2_X1 U15465 ( .A(_02960__PTR10), .B(_03190__PTR9), .Z(_03191__PTR10) );
  XOR2_X1 U15466 ( .A(_02960__PTR11), .B(_03190__PTR10), .Z(_03191__PTR11) );
  XOR2_X1 U15467 ( .A(_02960__PTR12), .B(_03190__PTR11), .Z(_03191__PTR12) );
  XOR2_X1 U15468 ( .A(_02960__PTR13), .B(_03190__PTR12), .Z(_03191__PTR13) );
  XOR2_X1 U15469 ( .A(_02960__PTR14), .B(_03190__PTR13), .Z(_03191__PTR14) );
  XOR2_X1 U15470 ( .A(_02960__PTR15), .B(_03190__PTR14), .Z(_03191__PTR15) );
  XOR2_X1 U15471 ( .A(_02960__PTR16), .B(_03190__PTR15), .Z(_03191__PTR16) );
  XOR2_X1 U15472 ( .A(_02960__PTR17), .B(_03190__PTR16), .Z(_03191__PTR17) );
  XOR2_X1 U15473 ( .A(_02960__PTR18), .B(_03190__PTR17), .Z(_03191__PTR18) );
  XOR2_X1 U15474 ( .A(_02960__PTR19), .B(_03190__PTR18), .Z(_03191__PTR19) );
  XOR2_X1 U15475 ( .A(_02960__PTR20), .B(_03190__PTR19), .Z(_03191__PTR20) );
  XOR2_X1 U15476 ( .A(_02960__PTR21), .B(_03190__PTR20), .Z(_03191__PTR21) );
  XOR2_X1 U15477 ( .A(_02960__PTR22), .B(_03190__PTR21), .Z(_03191__PTR22) );
  XOR2_X1 U15478 ( .A(_02960__PTR23), .B(_03190__PTR22), .Z(_03191__PTR23) );
  XOR2_X1 U15479 ( .A(_02960__PTR24), .B(_03190__PTR23), .Z(_03191__PTR24) );
  XOR2_X1 U15480 ( .A(_02960__PTR25), .B(_03190__PTR24), .Z(_03191__PTR25) );
  XOR2_X1 U15481 ( .A(_02960__PTR26), .B(_03190__PTR25), .Z(_03191__PTR26) );
  XOR2_X1 U15482 ( .A(_02960__PTR27), .B(_03190__PTR26), .Z(_03191__PTR27) );
  XOR2_X1 U15483 ( .A(_02960__PTR28), .B(_03190__PTR27), .Z(_03191__PTR28) );
  XOR2_X1 U15484 ( .A(_02960__PTR29), .B(_03190__PTR28), .Z(_03191__PTR29) );
  XOR2_X1 U15485 ( .A(_02960__PTR30), .B(_03190__PTR29), .Z(_03191__PTR30) );
  XOR2_X1 U15486 ( .A(_02958__PTR31), .B(_03190__PTR30), .Z(_03191__PTR31) );
  XOR2_X1 U15487 ( .A(P2_P1_PhyAddrPointer_PTR3), .B(P2_P1_PhyAddrPointer_PTR2), .Z(_03041__PTR1) );
  XOR2_X1 U15488 ( .A(P2_P1_PhyAddrPointer_PTR4), .B(_03039__PTR1), .Z(_03041__PTR2) );
  XOR2_X1 U15489 ( .A(P2_P1_PhyAddrPointer_PTR5), .B(_03039__PTR2), .Z(_03041__PTR3) );
  XOR2_X1 U15490 ( .A(P2_P1_PhyAddrPointer_PTR6), .B(_03039__PTR3), .Z(_03041__PTR4) );
  XOR2_X1 U15491 ( .A(P2_P1_PhyAddrPointer_PTR7), .B(_03039__PTR4), .Z(_03041__PTR5) );
  XOR2_X1 U15492 ( .A(P2_P1_PhyAddrPointer_PTR8), .B(_03039__PTR5), .Z(_03041__PTR6) );
  XOR2_X1 U15493 ( .A(P2_P1_PhyAddrPointer_PTR9), .B(_03039__PTR6), .Z(_03041__PTR7) );
  XOR2_X1 U15494 ( .A(P2_P1_PhyAddrPointer_PTR10), .B(_03039__PTR7), .Z(_03041__PTR8) );
  XOR2_X1 U15495 ( .A(P2_P1_PhyAddrPointer_PTR11), .B(_03039__PTR8), .Z(_03041__PTR9) );
  XOR2_X1 U15496 ( .A(P2_P1_PhyAddrPointer_PTR12), .B(_03039__PTR9), .Z(_03041__PTR10) );
  XOR2_X1 U15497 ( .A(P2_P1_PhyAddrPointer_PTR13), .B(_03039__PTR10), .Z(_03041__PTR11) );
  XOR2_X1 U15498 ( .A(P2_P1_PhyAddrPointer_PTR14), .B(_03039__PTR11), .Z(_03041__PTR12) );
  XOR2_X1 U15499 ( .A(P2_P1_PhyAddrPointer_PTR15), .B(_03039__PTR12), .Z(_03041__PTR13) );
  XOR2_X1 U15500 ( .A(P2_P1_PhyAddrPointer_PTR16), .B(_03039__PTR13), .Z(_03041__PTR14) );
  XOR2_X1 U15501 ( .A(P2_P1_PhyAddrPointer_PTR17), .B(_03039__PTR14), .Z(_03041__PTR15) );
  XOR2_X1 U15502 ( .A(P2_P1_PhyAddrPointer_PTR18), .B(_03039__PTR15), .Z(_03041__PTR16) );
  XOR2_X1 U15503 ( .A(P2_P1_PhyAddrPointer_PTR19), .B(_03039__PTR16), .Z(_03041__PTR17) );
  XOR2_X1 U15504 ( .A(P2_P1_PhyAddrPointer_PTR20), .B(_03039__PTR17), .Z(_03041__PTR18) );
  XOR2_X1 U15505 ( .A(P2_P1_PhyAddrPointer_PTR21), .B(_03039__PTR18), .Z(_03041__PTR19) );
  XOR2_X1 U15506 ( .A(P2_P1_PhyAddrPointer_PTR22), .B(_03039__PTR19), .Z(_03041__PTR20) );
  XOR2_X1 U15507 ( .A(P2_P1_PhyAddrPointer_PTR23), .B(_03039__PTR20), .Z(_03041__PTR21) );
  XOR2_X1 U15508 ( .A(P2_P1_PhyAddrPointer_PTR24), .B(_03039__PTR21), .Z(_03041__PTR22) );
  XOR2_X1 U15509 ( .A(P2_P1_PhyAddrPointer_PTR25), .B(_03039__PTR22), .Z(_03041__PTR23) );
  XOR2_X1 U15510 ( .A(P2_P1_PhyAddrPointer_PTR26), .B(_03039__PTR23), .Z(_03041__PTR24) );
  XOR2_X1 U15511 ( .A(P2_P1_PhyAddrPointer_PTR27), .B(_03039__PTR24), .Z(_03041__PTR25) );
  XOR2_X1 U15512 ( .A(P2_P1_PhyAddrPointer_PTR28), .B(_03039__PTR25), .Z(_03041__PTR26) );
  XOR2_X1 U15513 ( .A(P2_P1_PhyAddrPointer_PTR29), .B(_03039__PTR26), .Z(_03041__PTR27) );
  XOR2_X1 U15514 ( .A(P2_P1_PhyAddrPointer_PTR30), .B(_03039__PTR27), .Z(_03041__PTR28) );
  XOR2_X1 U15515 ( .A(P2_P1_PhyAddrPointer_PTR31), .B(_03039__PTR28), .Z(_03041__PTR29) );
  XOR2_X1 U15516 ( .A(P2_P1_InstQueueWr_Addr_PTR1), .B(P2_P1_InstQueueWr_Addr_PTR0), .Z(_02129__PTR1) );
  XOR2_X1 U15517 ( .A(P2_P1_InstQueueWr_Addr_PTR2), .B(_03024__PTR1), .Z(_02129__PTR2) );
  XOR2_X1 U15518 ( .A(P2_P1_InstQueueWr_Addr_PTR3), .B(_03024__PTR2), .Z(_02129__PTR3) );
  XOR2_X1 U15519 ( .A(_02129__PTR1), .B(_02129__PTR0), .Z(_02131__PTR1) );
  XOR2_X1 U15520 ( .A(_02129__PTR2), .B(_03025__PTR1), .Z(_02131__PTR2) );
  XOR2_X1 U15521 ( .A(_02129__PTR3), .B(_03025__PTR2), .Z(_02131__PTR3) );
  XOR2_X1 U15522 ( .A(_02131__PTR1), .B(P2_P1_InstQueueWr_Addr_PTR0), .Z(_02133__PTR1) );
  XOR2_X1 U15523 ( .A(_02131__PTR2), .B(_03030__PTR1), .Z(_02133__PTR2) );
  XOR2_X1 U15524 ( .A(_02131__PTR3), .B(_03030__PTR2), .Z(_02133__PTR3) );
  XOR2_X1 U15525 ( .A(_02133__PTR1), .B(_02129__PTR0), .Z(_03036__PTR1) );
  XOR2_X1 U15526 ( .A(_02133__PTR2), .B(_03035__PTR1), .Z(_03036__PTR2) );
  XOR2_X1 U15527 ( .A(_02133__PTR3), .B(_03035__PTR2), .Z(_03036__PTR3) );
  XOR2_X1 U15528 ( .A(di2_PTR25), .B(_03032__PTR0), .Z(_03034__PTR1) );
  XOR2_X1 U15529 ( .A(di2_PTR26), .B(_03032__PTR1), .Z(_03034__PTR2) );
  XOR2_X1 U15530 ( .A(di2_PTR27), .B(_03032__PTR2), .Z(_03034__PTR3) );
  XOR2_X1 U15531 ( .A(di2_PTR28), .B(_03032__PTR3), .Z(_03034__PTR4) );
  XOR2_X1 U15532 ( .A(di2_PTR29), .B(_03032__PTR4), .Z(_03034__PTR5) );
  XOR2_X1 U15533 ( .A(di2_PTR30), .B(_03032__PTR5), .Z(_03034__PTR6) );
  XOR2_X1 U15534 ( .A(P2_Datai_PTR31), .B(_03032__PTR6), .Z(_03034__PTR7) );
  XOR2_X1 U15535 ( .A(_03031_), .B(di2_PTR24), .Z(_03033__PTR0) );
  AND2_X1 U15536 ( .A1(_03031_), .A2(di2_PTR24), .ZN(_03032__PTR0) );
  XOR2_X1 U15537 ( .A(di2_PTR17), .B(_03027__PTR0), .Z(_03029__PTR1) );
  XOR2_X1 U15538 ( .A(di2_PTR18), .B(_03027__PTR1), .Z(_03029__PTR2) );
  XOR2_X1 U15539 ( .A(di2_PTR19), .B(_03027__PTR2), .Z(_03029__PTR3) );
  XOR2_X1 U15540 ( .A(di2_PTR20), .B(_03027__PTR3), .Z(_03029__PTR4) );
  XOR2_X1 U15541 ( .A(di2_PTR21), .B(_03027__PTR4), .Z(_03029__PTR5) );
  XOR2_X1 U15542 ( .A(di2_PTR22), .B(_03027__PTR5), .Z(_03029__PTR6) );
  XOR2_X1 U15543 ( .A(di2_PTR23), .B(_03027__PTR6), .Z(_03029__PTR7) );
  XOR2_X1 U15544 ( .A(_03026_), .B(di2_PTR16), .Z(_03028__PTR0) );
  AND2_X1 U15545 ( .A1(_03026_), .A2(di2_PTR16), .ZN(_03027__PTR0) );
  XOR2_X1 U15546 ( .A(P2_rEIP_PTR2), .B(_03023__PTR0), .Z(_02172__PTR193) );
  XOR2_X1 U15547 ( .A(P2_rEIP_PTR3), .B(_03023__PTR1), .Z(_02172__PTR194) );
  XOR2_X1 U15548 ( .A(P2_rEIP_PTR4), .B(_03023__PTR2), .Z(_02172__PTR195) );
  XOR2_X1 U15549 ( .A(P2_rEIP_PTR5), .B(_03023__PTR3), .Z(_02172__PTR196) );
  XOR2_X1 U15550 ( .A(P2_rEIP_PTR6), .B(_03023__PTR4), .Z(_02172__PTR197) );
  XOR2_X1 U15551 ( .A(P2_rEIP_PTR7), .B(_03023__PTR5), .Z(_02172__PTR198) );
  XOR2_X1 U15552 ( .A(P2_rEIP_PTR8), .B(_03023__PTR6), .Z(_02172__PTR199) );
  XOR2_X1 U15553 ( .A(P2_rEIP_PTR9), .B(_03023__PTR7), .Z(_02172__PTR200) );
  XOR2_X1 U15554 ( .A(P2_rEIP_PTR10), .B(_03023__PTR8), .Z(_02172__PTR201) );
  XOR2_X1 U15555 ( .A(P2_rEIP_PTR11), .B(_03023__PTR9), .Z(_02172__PTR202) );
  XOR2_X1 U15556 ( .A(P2_rEIP_PTR12), .B(_03023__PTR10), .Z(_02172__PTR203) );
  XOR2_X1 U15557 ( .A(P2_rEIP_PTR13), .B(_03023__PTR11), .Z(_02172__PTR204) );
  XOR2_X1 U15558 ( .A(P2_rEIP_PTR14), .B(_03023__PTR12), .Z(_02172__PTR205) );
  XOR2_X1 U15559 ( .A(P2_rEIP_PTR15), .B(_03023__PTR13), .Z(_02172__PTR206) );
  XOR2_X1 U15560 ( .A(P2_rEIP_PTR16), .B(_03023__PTR14), .Z(_02172__PTR207) );
  XOR2_X1 U15561 ( .A(P2_rEIP_PTR17), .B(_03023__PTR15), .Z(_02172__PTR208) );
  XOR2_X1 U15562 ( .A(P2_rEIP_PTR18), .B(_03023__PTR16), .Z(_02172__PTR209) );
  XOR2_X1 U15563 ( .A(P2_rEIP_PTR19), .B(_03023__PTR17), .Z(_02172__PTR210) );
  XOR2_X1 U15564 ( .A(P2_rEIP_PTR20), .B(_03023__PTR18), .Z(_02172__PTR211) );
  XOR2_X1 U15565 ( .A(P2_rEIP_PTR21), .B(_03023__PTR19), .Z(_02172__PTR212) );
  XOR2_X1 U15566 ( .A(P2_rEIP_PTR22), .B(_03023__PTR20), .Z(_02172__PTR213) );
  XOR2_X1 U15567 ( .A(P2_rEIP_PTR23), .B(_03023__PTR21), .Z(_02172__PTR214) );
  XOR2_X1 U15568 ( .A(P2_rEIP_PTR24), .B(_03023__PTR22), .Z(_02172__PTR215) );
  XOR2_X1 U15569 ( .A(P2_rEIP_PTR25), .B(_03023__PTR23), .Z(_02172__PTR216) );
  XOR2_X1 U15570 ( .A(P2_rEIP_PTR26), .B(_03023__PTR24), .Z(_02172__PTR217) );
  XOR2_X1 U15571 ( .A(P2_rEIP_PTR27), .B(_03023__PTR25), .Z(_02172__PTR218) );
  XOR2_X1 U15572 ( .A(P2_rEIP_PTR28), .B(_03023__PTR26), .Z(_02172__PTR219) );
  XOR2_X1 U15573 ( .A(P2_rEIP_PTR29), .B(_03023__PTR27), .Z(_02172__PTR220) );
  XOR2_X1 U15574 ( .A(P2_rEIP_PTR30), .B(_03023__PTR28), .Z(_02172__PTR221) );
  XOR2_X1 U15575 ( .A(_03022_), .B(P2_rEIP_PTR1), .Z(_02172__PTR192) );
  AND2_X1 U15576 ( .A1(_03022_), .A2(P2_rEIP_PTR1), .ZN(_03023__PTR0) );
  XOR2_X1 U15577 ( .A(P2_rEIP_PTR3), .B(_03038__PTR0), .Z(_02172__PTR65) );
  XOR2_X1 U15578 ( .A(P2_rEIP_PTR4), .B(_03038__PTR1), .Z(_02172__PTR66) );
  XOR2_X1 U15579 ( .A(P2_rEIP_PTR5), .B(_03038__PTR2), .Z(_02172__PTR67) );
  XOR2_X1 U15580 ( .A(P2_rEIP_PTR6), .B(_03038__PTR3), .Z(_02172__PTR68) );
  XOR2_X1 U15581 ( .A(P2_rEIP_PTR7), .B(_03038__PTR4), .Z(_02172__PTR69) );
  XOR2_X1 U15582 ( .A(P2_rEIP_PTR8), .B(_03038__PTR5), .Z(_02172__PTR70) );
  XOR2_X1 U15583 ( .A(P2_rEIP_PTR9), .B(_03038__PTR6), .Z(_02172__PTR71) );
  XOR2_X1 U15584 ( .A(P2_rEIP_PTR10), .B(_03038__PTR7), .Z(_02172__PTR72) );
  XOR2_X1 U15585 ( .A(P2_rEIP_PTR11), .B(_03038__PTR8), .Z(_02172__PTR73) );
  XOR2_X1 U15586 ( .A(P2_rEIP_PTR12), .B(_03038__PTR9), .Z(_02172__PTR74) );
  XOR2_X1 U15587 ( .A(P2_rEIP_PTR13), .B(_03038__PTR10), .Z(_02172__PTR75) );
  XOR2_X1 U15588 ( .A(P2_rEIP_PTR14), .B(_03038__PTR11), .Z(_02172__PTR76) );
  XOR2_X1 U15589 ( .A(P2_rEIP_PTR15), .B(_03038__PTR12), .Z(_02172__PTR77) );
  XOR2_X1 U15590 ( .A(P2_rEIP_PTR16), .B(_03038__PTR13), .Z(_02172__PTR78) );
  XOR2_X1 U15591 ( .A(P2_rEIP_PTR17), .B(_03038__PTR14), .Z(_02172__PTR79) );
  XOR2_X1 U15592 ( .A(P2_rEIP_PTR18), .B(_03038__PTR15), .Z(_02172__PTR80) );
  XOR2_X1 U15593 ( .A(P2_rEIP_PTR19), .B(_03038__PTR16), .Z(_02172__PTR81) );
  XOR2_X1 U15594 ( .A(P2_rEIP_PTR20), .B(_03038__PTR17), .Z(_02172__PTR82) );
  XOR2_X1 U15595 ( .A(P2_rEIP_PTR21), .B(_03038__PTR18), .Z(_02172__PTR83) );
  XOR2_X1 U15596 ( .A(P2_rEIP_PTR22), .B(_03038__PTR19), .Z(_02172__PTR84) );
  XOR2_X1 U15597 ( .A(P2_rEIP_PTR23), .B(_03038__PTR20), .Z(_02172__PTR85) );
  XOR2_X1 U15598 ( .A(P2_rEIP_PTR24), .B(_03038__PTR21), .Z(_02172__PTR86) );
  XOR2_X1 U15599 ( .A(P2_rEIP_PTR25), .B(_03038__PTR22), .Z(_02172__PTR87) );
  XOR2_X1 U15600 ( .A(P2_rEIP_PTR26), .B(_03038__PTR23), .Z(_02172__PTR88) );
  XOR2_X1 U15601 ( .A(P2_rEIP_PTR27), .B(_03038__PTR24), .Z(_02172__PTR89) );
  XOR2_X1 U15602 ( .A(P2_rEIP_PTR28), .B(_03038__PTR25), .Z(_02172__PTR90) );
  XOR2_X1 U15603 ( .A(P2_rEIP_PTR29), .B(_03038__PTR26), .Z(_02172__PTR91) );
  XOR2_X1 U15604 ( .A(P2_rEIP_PTR30), .B(_03038__PTR27), .Z(_02172__PTR92) );
  XOR2_X1 U15605 ( .A(P2_rEIP_PTR31), .B(_03038__PTR28), .Z(_02172__PTR93) );
  XOR2_X1 U15606 ( .A(_03037_), .B(P2_rEIP_PTR2), .Z(_02172__PTR64) );
  AND2_X1 U15607 ( .A1(_03037_), .A2(P2_rEIP_PTR2), .ZN(_03038__PTR0) );
  XOR2_X1 U15608 ( .A(_03433__PTR4), .B(_03434__PTR3), .Z(_03236__PTR4) );
  XOR2_X1 U15609 ( .A(_03319__PTR1), .B(P3_P1_InstAddrPointer_PTR0), .Z(_03321__PTR1) );
  XOR2_X1 U15610 ( .A(_02662__PTR33), .B(_02662__PTR0), .Z(_03439__PTR1) );
  XOR2_X1 U15611 ( .A(_03431__PTR4), .B(_03432__PTR3), .Z(_03229__PTR4) );
  XOR2_X1 U15612 ( .A(_02513__PTR40), .B(_02418__PTR0), .Z(_03227__PTR0) );
  XOR2_X1 U15613 ( .A(_02513__PTR41), .B(_03225__PTR1), .Z(_03227__PTR1) );
  XOR2_X1 U15614 ( .A(_02513__PTR42), .B(_03225__PTR2), .Z(_03227__PTR2) );
  XOR2_X1 U15615 ( .A(_02513__PTR43), .B(_03225__PTR3), .Z(_03227__PTR3) );
  XOR2_X1 U15616 ( .A(_02513__PTR44), .B(_03225__PTR4), .Z(_03227__PTR4) );
  AND2_X1 U15617 ( .A1(_02513__PTR40), .A2(_02418__PTR0), .ZN(_03228__PTR0) );
  AND2_X1 U15618 ( .A1(_02513__PTR41), .A2(_03225__PTR1), .ZN(_03228__PTR1) );
  AND2_X1 U15619 ( .A1(_02513__PTR42), .A2(_03225__PTR2), .ZN(_03228__PTR2) );
  AND2_X1 U15620 ( .A1(_02513__PTR43), .A2(_03225__PTR3), .ZN(_03228__PTR3) );
  AND2_X1 U15621 ( .A1(_02513__PTR44), .A2(_03225__PTR4), .ZN(_03228__PTR4) );
  XOR2_X1 U15622 ( .A(P3_EBX_PTR1), .B(P3_EBX_PTR0), .Z(_02678__PTR33) );
  XOR2_X1 U15623 ( .A(P3_EBX_PTR2), .B(_03318__PTR1), .Z(_02678__PTR34) );
  XOR2_X1 U15624 ( .A(P3_EBX_PTR3), .B(_03318__PTR2), .Z(_02678__PTR35) );
  XOR2_X1 U15625 ( .A(P3_EBX_PTR4), .B(_03318__PTR3), .Z(_02678__PTR36) );
  XOR2_X1 U15626 ( .A(P3_EBX_PTR5), .B(_03318__PTR4), .Z(_02678__PTR37) );
  XOR2_X1 U15627 ( .A(P3_EBX_PTR6), .B(_03318__PTR5), .Z(_02678__PTR38) );
  XOR2_X1 U15628 ( .A(P3_EBX_PTR7), .B(_03318__PTR6), .Z(_02678__PTR39) );
  XOR2_X1 U15629 ( .A(P3_EBX_PTR8), .B(_03318__PTR7), .Z(_02678__PTR40) );
  XOR2_X1 U15630 ( .A(P3_EBX_PTR9), .B(_03318__PTR8), .Z(_02678__PTR41) );
  XOR2_X1 U15631 ( .A(P3_EBX_PTR10), .B(_03318__PTR9), .Z(_02678__PTR42) );
  XOR2_X1 U15632 ( .A(P3_EBX_PTR11), .B(_03318__PTR10), .Z(_02678__PTR43) );
  XOR2_X1 U15633 ( .A(P3_EBX_PTR12), .B(_03318__PTR11), .Z(_02678__PTR44) );
  XOR2_X1 U15634 ( .A(P3_EBX_PTR13), .B(_03318__PTR12), .Z(_02678__PTR45) );
  XOR2_X1 U15635 ( .A(P3_EBX_PTR14), .B(_03318__PTR13), .Z(_02678__PTR46) );
  XOR2_X1 U15636 ( .A(P3_EBX_PTR15), .B(_03318__PTR14), .Z(_02678__PTR47) );
  XOR2_X1 U15637 ( .A(P3_EBX_PTR16), .B(_03318__PTR15), .Z(_02678__PTR48) );
  XOR2_X1 U15638 ( .A(P3_EBX_PTR17), .B(_03318__PTR16), .Z(_02678__PTR49) );
  XOR2_X1 U15639 ( .A(P3_EBX_PTR18), .B(_03318__PTR17), .Z(_02678__PTR50) );
  XOR2_X1 U15640 ( .A(P3_EBX_PTR19), .B(_03318__PTR18), .Z(_02678__PTR51) );
  XOR2_X1 U15641 ( .A(P3_EBX_PTR20), .B(_03318__PTR19), .Z(_02678__PTR52) );
  XOR2_X1 U15642 ( .A(P3_EBX_PTR21), .B(_03318__PTR20), .Z(_02678__PTR53) );
  XOR2_X1 U15643 ( .A(P3_EBX_PTR22), .B(_03318__PTR21), .Z(_02678__PTR54) );
  XOR2_X1 U15644 ( .A(P3_EBX_PTR23), .B(_03318__PTR22), .Z(_02678__PTR55) );
  XOR2_X1 U15645 ( .A(P3_EBX_PTR24), .B(_03318__PTR23), .Z(_02678__PTR56) );
  XOR2_X1 U15646 ( .A(P3_EBX_PTR25), .B(_03318__PTR24), .Z(_02678__PTR57) );
  XOR2_X1 U15647 ( .A(P3_EBX_PTR26), .B(_03318__PTR25), .Z(_02678__PTR58) );
  XOR2_X1 U15648 ( .A(P3_EBX_PTR27), .B(_03318__PTR26), .Z(_02678__PTR59) );
  XOR2_X1 U15649 ( .A(P3_EBX_PTR28), .B(_03318__PTR27), .Z(_02678__PTR60) );
  XOR2_X1 U15650 ( .A(P3_EBX_PTR29), .B(_03318__PTR28), .Z(_02678__PTR61) );
  XOR2_X1 U15651 ( .A(P3_EBX_PTR30), .B(_03318__PTR29), .Z(_02678__PTR62) );
  XOR2_X1 U15652 ( .A(P3_EBX_PTR31), .B(_03318__PTR30), .Z(_02678__PTR63) );
  XOR2_X1 U15653 ( .A(P3_EAX_PTR1), .B(P3_EAX_PTR0), .Z(_02674__PTR33) );
  XOR2_X1 U15654 ( .A(P3_EAX_PTR2), .B(_03317__PTR1), .Z(_02674__PTR34) );
  XOR2_X1 U15655 ( .A(P3_EAX_PTR3), .B(_03317__PTR2), .Z(_02674__PTR35) );
  XOR2_X1 U15656 ( .A(P3_EAX_PTR4), .B(_03317__PTR3), .Z(_02674__PTR36) );
  XOR2_X1 U15657 ( .A(P3_EAX_PTR5), .B(_03317__PTR4), .Z(_02674__PTR37) );
  XOR2_X1 U15658 ( .A(P3_EAX_PTR6), .B(_03317__PTR5), .Z(_02674__PTR38) );
  XOR2_X1 U15659 ( .A(P3_EAX_PTR7), .B(_03317__PTR6), .Z(_02674__PTR39) );
  XOR2_X1 U15660 ( .A(P3_EAX_PTR8), .B(_03317__PTR7), .Z(_02674__PTR40) );
  XOR2_X1 U15661 ( .A(P3_EAX_PTR9), .B(_03317__PTR8), .Z(_02674__PTR41) );
  XOR2_X1 U15662 ( .A(P3_EAX_PTR10), .B(_03317__PTR9), .Z(_02674__PTR42) );
  XOR2_X1 U15663 ( .A(P3_EAX_PTR11), .B(_03317__PTR10), .Z(_02674__PTR43) );
  XOR2_X1 U15664 ( .A(P3_EAX_PTR12), .B(_03317__PTR11), .Z(_02674__PTR44) );
  XOR2_X1 U15665 ( .A(P3_EAX_PTR13), .B(_03317__PTR12), .Z(_02674__PTR45) );
  XOR2_X1 U15666 ( .A(P3_EAX_PTR14), .B(_03317__PTR13), .Z(_02674__PTR46) );
  XOR2_X1 U15667 ( .A(P3_EAX_PTR15), .B(_03317__PTR14), .Z(_02674__PTR47) );
  XOR2_X1 U15668 ( .A(P3_EAX_PTR16), .B(_03317__PTR15), .Z(_02674__PTR48) );
  XOR2_X1 U15669 ( .A(P3_EAX_PTR17), .B(_03317__PTR16), .Z(_02674__PTR49) );
  XOR2_X1 U15670 ( .A(P3_EAX_PTR18), .B(_03317__PTR17), .Z(_02674__PTR50) );
  XOR2_X1 U15671 ( .A(P3_EAX_PTR19), .B(_03317__PTR18), .Z(_02674__PTR51) );
  XOR2_X1 U15672 ( .A(P3_EAX_PTR20), .B(_03317__PTR19), .Z(_02674__PTR52) );
  XOR2_X1 U15673 ( .A(P3_EAX_PTR21), .B(_03317__PTR20), .Z(_02674__PTR53) );
  XOR2_X1 U15674 ( .A(P3_EAX_PTR22), .B(_03317__PTR21), .Z(_02674__PTR54) );
  XOR2_X1 U15675 ( .A(P3_EAX_PTR23), .B(_03317__PTR22), .Z(_02674__PTR55) );
  XOR2_X1 U15676 ( .A(P3_EAX_PTR24), .B(_03317__PTR23), .Z(_02674__PTR56) );
  XOR2_X1 U15677 ( .A(P3_EAX_PTR25), .B(_03317__PTR24), .Z(_02674__PTR57) );
  XOR2_X1 U15678 ( .A(P3_EAX_PTR26), .B(_03317__PTR25), .Z(_02674__PTR58) );
  XOR2_X1 U15679 ( .A(P3_EAX_PTR27), .B(_03317__PTR26), .Z(_02674__PTR59) );
  XOR2_X1 U15680 ( .A(P3_EAX_PTR28), .B(_03317__PTR27), .Z(_02674__PTR60) );
  XOR2_X1 U15681 ( .A(P3_EAX_PTR29), .B(_03317__PTR28), .Z(_02674__PTR61) );
  XOR2_X1 U15682 ( .A(P3_EAX_PTR30), .B(_03317__PTR29), .Z(_02674__PTR62) );
  XOR2_X1 U15683 ( .A(P3_EAX_PTR31), .B(_03317__PTR30), .Z(_02674__PTR63) );
  XOR2_X1 U15684 ( .A(P3_EAX_PTR17), .B(_03314__PTR0), .Z(_03316__PTR1) );
  XOR2_X1 U15685 ( .A(P3_EAX_PTR18), .B(_03314__PTR1), .Z(_03316__PTR2) );
  XOR2_X1 U15686 ( .A(P3_EAX_PTR19), .B(_03314__PTR2), .Z(_03316__PTR3) );
  XOR2_X1 U15687 ( .A(P3_EAX_PTR20), .B(_03314__PTR3), .Z(_03316__PTR4) );
  XOR2_X1 U15688 ( .A(P3_EAX_PTR21), .B(_03314__PTR4), .Z(_03316__PTR5) );
  XOR2_X1 U15689 ( .A(P3_EAX_PTR22), .B(_03314__PTR5), .Z(_03316__PTR6) );
  XOR2_X1 U15690 ( .A(P3_EAX_PTR23), .B(_03314__PTR6), .Z(_03316__PTR7) );
  XOR2_X1 U15691 ( .A(P3_EAX_PTR24), .B(_03314__PTR7), .Z(_03316__PTR8) );
  XOR2_X1 U15692 ( .A(P3_EAX_PTR25), .B(_03314__PTR8), .Z(_03316__PTR9) );
  XOR2_X1 U15693 ( .A(P3_EAX_PTR26), .B(_03314__PTR9), .Z(_03316__PTR10) );
  XOR2_X1 U15694 ( .A(P3_EAX_PTR27), .B(_03314__PTR10), .Z(_03316__PTR11) );
  XOR2_X1 U15695 ( .A(P3_EAX_PTR28), .B(_03314__PTR11), .Z(_03316__PTR12) );
  XOR2_X1 U15696 ( .A(P3_EAX_PTR29), .B(_03314__PTR12), .Z(_03316__PTR13) );
  XOR2_X1 U15697 ( .A(P3_EAX_PTR30), .B(_03314__PTR13), .Z(_03316__PTR14) );
  XOR2_X1 U15698 ( .A(_03313_), .B(P3_EAX_PTR16), .Z(_03315__PTR0) );
  AND2_X1 U15699 ( .A1(_03313_), .A2(P3_EAX_PTR16), .ZN(_03314__PTR0) );
  XOR2_X1 U15700 ( .A(P3_rEIP_PTR2), .B(P3_rEIP_PTR1), .Z(_03312__PTR1) );
  XOR2_X1 U15701 ( .A(P3_rEIP_PTR3), .B(_03311__PTR1), .Z(_03312__PTR2) );
  XOR2_X1 U15702 ( .A(P3_rEIP_PTR4), .B(_03311__PTR2), .Z(_03312__PTR3) );
  XOR2_X1 U15703 ( .A(P3_rEIP_PTR5), .B(_03311__PTR3), .Z(_03312__PTR4) );
  XOR2_X1 U15704 ( .A(P3_rEIP_PTR6), .B(_03311__PTR4), .Z(_03312__PTR5) );
  XOR2_X1 U15705 ( .A(P3_rEIP_PTR7), .B(_03311__PTR5), .Z(_03312__PTR6) );
  XOR2_X1 U15706 ( .A(P3_rEIP_PTR8), .B(_03311__PTR6), .Z(_03312__PTR7) );
  XOR2_X1 U15707 ( .A(P3_rEIP_PTR9), .B(_03311__PTR7), .Z(_03312__PTR8) );
  XOR2_X1 U15708 ( .A(P3_rEIP_PTR10), .B(_03311__PTR8), .Z(_03312__PTR9) );
  XOR2_X1 U15709 ( .A(P3_rEIP_PTR11), .B(_03311__PTR9), .Z(_03312__PTR10) );
  XOR2_X1 U15710 ( .A(P3_rEIP_PTR12), .B(_03311__PTR10), .Z(_03312__PTR11) );
  XOR2_X1 U15711 ( .A(P3_rEIP_PTR13), .B(_03311__PTR11), .Z(_03312__PTR12) );
  XOR2_X1 U15712 ( .A(P3_rEIP_PTR14), .B(_03311__PTR12), .Z(_03312__PTR13) );
  XOR2_X1 U15713 ( .A(P3_rEIP_PTR15), .B(_03311__PTR13), .Z(_03312__PTR14) );
  XOR2_X1 U15714 ( .A(P3_rEIP_PTR16), .B(_03311__PTR14), .Z(_03312__PTR15) );
  XOR2_X1 U15715 ( .A(P3_rEIP_PTR17), .B(_03311__PTR15), .Z(_03312__PTR16) );
  XOR2_X1 U15716 ( .A(P3_rEIP_PTR18), .B(_03311__PTR16), .Z(_03312__PTR17) );
  XOR2_X1 U15717 ( .A(P3_rEIP_PTR19), .B(_03311__PTR17), .Z(_03312__PTR18) );
  XOR2_X1 U15718 ( .A(P3_rEIP_PTR20), .B(_03311__PTR18), .Z(_03312__PTR19) );
  XOR2_X1 U15719 ( .A(P3_rEIP_PTR21), .B(_03311__PTR19), .Z(_03312__PTR20) );
  XOR2_X1 U15720 ( .A(P3_rEIP_PTR22), .B(_03311__PTR20), .Z(_03312__PTR21) );
  XOR2_X1 U15721 ( .A(P3_rEIP_PTR23), .B(_03311__PTR21), .Z(_03312__PTR22) );
  XOR2_X1 U15722 ( .A(P3_rEIP_PTR24), .B(_03311__PTR22), .Z(_03312__PTR23) );
  XOR2_X1 U15723 ( .A(P3_rEIP_PTR25), .B(_03311__PTR23), .Z(_03312__PTR24) );
  XOR2_X1 U15724 ( .A(P3_rEIP_PTR26), .B(_03311__PTR24), .Z(_03312__PTR25) );
  XOR2_X1 U15725 ( .A(P3_rEIP_PTR27), .B(_03311__PTR25), .Z(_03312__PTR26) );
  XOR2_X1 U15726 ( .A(P3_rEIP_PTR28), .B(_03311__PTR26), .Z(_03312__PTR27) );
  XOR2_X1 U15727 ( .A(P3_rEIP_PTR29), .B(_03311__PTR27), .Z(_03312__PTR28) );
  XOR2_X1 U15728 ( .A(P3_rEIP_PTR30), .B(_03311__PTR28), .Z(_03312__PTR29) );
  XOR2_X1 U15729 ( .A(P3_rEIP_PTR31), .B(_03311__PTR29), .Z(_03312__PTR30) );
  XOR2_X1 U15730 ( .A(_03224__PTR1), .B(_02678__PTR32), .Z(_03438__PTR1) );
  XOR2_X1 U15731 ( .A(_03224__PTR2), .B(_03437__PTR1), .Z(_03438__PTR2) );
  XOR2_X1 U15732 ( .A(_03224__PTR3), .B(_03437__PTR2), .Z(_03438__PTR3) );
  XOR2_X1 U15733 ( .A(_03224__PTR4), .B(_03437__PTR3), .Z(_03438__PTR4) );
  XOR2_X1 U15734 ( .A(_03224__PTR5), .B(_03437__PTR4), .Z(_03438__PTR5) );
  XOR2_X1 U15735 ( .A(_03224__PTR6), .B(_03437__PTR5), .Z(_03438__PTR6) );
  XOR2_X1 U15736 ( .A(_03224__PTR7), .B(_03437__PTR6), .Z(_03438__PTR7) );
  XOR2_X1 U15737 ( .A(_03224__PTR8), .B(_03437__PTR7), .Z(_03438__PTR8) );
  XOR2_X1 U15738 ( .A(_03224__PTR9), .B(_03437__PTR8), .Z(_03438__PTR9) );
  XOR2_X1 U15739 ( .A(_03224__PTR10), .B(_03437__PTR9), .Z(_03438__PTR10) );
  XOR2_X1 U15740 ( .A(_03224__PTR11), .B(_03437__PTR10), .Z(_03438__PTR11) );
  XOR2_X1 U15741 ( .A(_03224__PTR12), .B(_03437__PTR11), .Z(_03438__PTR12) );
  XOR2_X1 U15742 ( .A(_03224__PTR13), .B(_03437__PTR12), .Z(_03438__PTR13) );
  XOR2_X1 U15743 ( .A(_03224__PTR14), .B(_03437__PTR13), .Z(_03438__PTR14) );
  XOR2_X1 U15744 ( .A(_03224__PTR15), .B(_03437__PTR14), .Z(_03438__PTR15) );
  XOR2_X1 U15745 ( .A(_03224__PTR16), .B(_03437__PTR15), .Z(_03438__PTR16) );
  XOR2_X1 U15746 ( .A(_03224__PTR17), .B(_03437__PTR16), .Z(_03438__PTR17) );
  XOR2_X1 U15747 ( .A(_03224__PTR18), .B(_03437__PTR17), .Z(_03438__PTR18) );
  XOR2_X1 U15748 ( .A(_03224__PTR19), .B(_03437__PTR18), .Z(_03438__PTR19) );
  XOR2_X1 U15749 ( .A(_03224__PTR20), .B(_03437__PTR19), .Z(_03438__PTR20) );
  XOR2_X1 U15750 ( .A(_03224__PTR21), .B(_03437__PTR20), .Z(_03438__PTR21) );
  XOR2_X1 U15751 ( .A(_03224__PTR22), .B(_03437__PTR21), .Z(_03438__PTR22) );
  XOR2_X1 U15752 ( .A(_03224__PTR23), .B(_03437__PTR22), .Z(_03438__PTR23) );
  XOR2_X1 U15753 ( .A(_03224__PTR24), .B(_03437__PTR23), .Z(_03438__PTR24) );
  XOR2_X1 U15754 ( .A(_03224__PTR25), .B(_03437__PTR24), .Z(_03438__PTR25) );
  XOR2_X1 U15755 ( .A(_03224__PTR26), .B(_03437__PTR25), .Z(_03438__PTR26) );
  XOR2_X1 U15756 ( .A(_03224__PTR27), .B(_03437__PTR26), .Z(_03438__PTR27) );
  XOR2_X1 U15757 ( .A(_03224__PTR28), .B(_03437__PTR27), .Z(_03438__PTR28) );
  XOR2_X1 U15758 ( .A(_03224__PTR29), .B(_03437__PTR28), .Z(_03438__PTR29) );
  XOR2_X1 U15759 ( .A(_03224__PTR30), .B(_03437__PTR29), .Z(_03438__PTR30) );
  XOR2_X1 U15760 ( .A(_03222__PTR31), .B(_03437__PTR30), .Z(_03438__PTR31) );
  XOR2_X1 U15761 ( .A(_03422__PTR1), .B(_03421__PTR0), .Z(_03207__PTR1) );
  XOR2_X1 U15762 ( .A(_03422__PTR2), .B(_03421__PTR1), .Z(_03207__PTR2) );
  XOR2_X1 U15763 ( .A(_03422__PTR3), .B(_03421__PTR2), .Z(_03207__PTR3) );
  XOR2_X1 U15764 ( .A(_03422__PTR4), .B(_03421__PTR3), .Z(_03207__PTR4) );
  XOR2_X1 U15765 ( .A(P3_P1_InstQueueWr_Addr_PTR0), .B(_02465__PTR3), .Z(_03208__PTR0) );
  XOR2_X1 U15766 ( .A(P3_P1_InstQueueWr_Addr_PTR1), .B(_02471__PTR4), .Z(_03422__PTR1) );
  XOR2_X1 U15767 ( .A(P3_P1_InstQueueWr_Addr_PTR2), .B(_02467__PTR5), .Z(_03422__PTR2) );
  XOR2_X1 U15768 ( .A(P3_P1_InstQueueWr_Addr_PTR3), .B(_03420__PTR3), .Z(_03422__PTR3) );
  XOR2_X1 U15769 ( .A(P3_P1_InstQueueWr_Addr_PTR4), .B(_03241__PTR4), .Z(_03422__PTR4) );
  AND2_X1 U15770 ( .A1(P3_P1_InstQueueWr_Addr_PTR0), .A2(_02465__PTR3), .ZN(_03423__PTR0) );
  AND2_X1 U15771 ( .A1(P3_P1_InstQueueWr_Addr_PTR1), .A2(_02471__PTR4), .ZN(_03423__PTR1) );
  AND2_X1 U15772 ( .A1(P3_P1_InstQueueWr_Addr_PTR2), .A2(_02467__PTR5), .ZN(_03423__PTR2) );
  AND2_X1 U15773 ( .A1(P3_P1_InstQueueWr_Addr_PTR3), .A2(_03420__PTR3), .ZN(_03423__PTR3) );
  AND2_X1 U15774 ( .A1(P3_P1_InstQueueWr_Addr_PTR4), .A2(_03241__PTR4), .ZN(_03423__PTR4) );
  XOR2_X1 U15775 ( .A(P3_P1_InstQueueRd_Addr_PTR1), .B(P3_P1_InstQueueRd_Addr_PTR0), .Z(_02465__PTR4) );
  XOR2_X1 U15776 ( .A(_02467__PTR5), .B(_03240__PTR1), .Z(_03310__PTR2) );
  XOR2_X1 U15777 ( .A(P3_P1_InstQueueRd_Addr_PTR3), .B(_03309__PTR2), .Z(_03310__PTR3) );
  XOR2_X1 U15778 ( .A(P3_P1_InstQueueRd_Addr_PTR2), .B(P3_P1_InstQueueRd_Addr_PTR1), .Z(_02471__PTR5) );
  XOR2_X1 U15779 ( .A(P3_P1_InstQueueRd_Addr_PTR3), .B(_03307__PTR1), .Z(_02471__PTR6) );
  XOR2_X1 U15780 ( .A(P3_P1_InstQueueRd_Addr_PTR4), .B(_03307__PTR2), .Z(_03308__PTR3) );
  XOR2_X1 U15781 ( .A(_02468__PTR1), .B(_03304__PTR0), .Z(_03306__PTR1) );
  XOR2_X1 U15782 ( .A(_02468__PTR2), .B(_03304__PTR1), .Z(_03306__PTR2) );
  XOR2_X1 U15783 ( .A(_02468__PTR3), .B(_03304__PTR2), .Z(_03306__PTR3) );
  XOR2_X1 U15784 ( .A(_02468__PTR4), .B(_03304__PTR3), .Z(_03306__PTR4) );
  XOR2_X1 U15785 ( .A(_02468__PTR5), .B(_03304__PTR4), .Z(_03306__PTR5) );
  XOR2_X1 U15786 ( .A(_02468__PTR6), .B(_03304__PTR5), .Z(_03306__PTR6) );
  XOR2_X1 U15787 ( .A(_02468__PTR7), .B(_03304__PTR6), .Z(_03306__PTR7) );
  XOR2_X1 U15788 ( .A(_02468__PTR0), .B(_02470__PTR7), .Z(_03305__PTR0) );
  AND2_X1 U15789 ( .A1(_02468__PTR0), .A2(_02470__PTR7), .ZN(_03304__PTR0) );
  XOR2_X1 U15790 ( .A(_02471__PTR4), .B(P3_P1_InstQueueRd_Addr_PTR0), .Z(_02469__PTR4) );
  XOR2_X1 U15791 ( .A(P3_P1_InstQueueRd_Addr_PTR2), .B(_03303__PTR1), .Z(_02469__PTR5) );
  XOR2_X1 U15792 ( .A(P3_P1_InstQueueRd_Addr_PTR3), .B(_03303__PTR2), .Z(_02469__PTR6) );
  XOR2_X1 U15793 ( .A(P3_P1_InstQueueRd_Addr_PTR3), .B(P3_P1_InstQueueRd_Addr_PTR2), .Z(_02467__PTR6) );
  XOR2_X1 U15794 ( .A(P3_P1_InstAddrPointer_PTR1), .B(P3_P1_InstAddrPointer_PTR0), .Z(_02662__PTR1) );
  XOR2_X1 U15795 ( .A(_03235__PTR2), .B(_03288__PTR1), .Z(_03297__PTR2) );
  XOR2_X1 U15796 ( .A(P3_P1_InstAddrPointer_PTR3), .B(_03296__PTR2), .Z(_03297__PTR3) );
  XOR2_X1 U15797 ( .A(P3_P1_InstAddrPointer_PTR4), .B(_03296__PTR3), .Z(_03297__PTR4) );
  XOR2_X1 U15798 ( .A(P3_P1_InstAddrPointer_PTR5), .B(_03296__PTR4), .Z(_03297__PTR5) );
  XOR2_X1 U15799 ( .A(P3_P1_InstAddrPointer_PTR6), .B(_03296__PTR5), .Z(_03297__PTR6) );
  XOR2_X1 U15800 ( .A(P3_P1_InstAddrPointer_PTR7), .B(_03296__PTR6), .Z(_03297__PTR7) );
  XOR2_X1 U15801 ( .A(P3_P1_InstAddrPointer_PTR8), .B(_03296__PTR7), .Z(_03297__PTR8) );
  XOR2_X1 U15802 ( .A(P3_P1_InstAddrPointer_PTR9), .B(_03296__PTR8), .Z(_03297__PTR9) );
  XOR2_X1 U15803 ( .A(P3_P1_InstAddrPointer_PTR10), .B(_03296__PTR9), .Z(_03297__PTR10) );
  XOR2_X1 U15804 ( .A(P3_P1_InstAddrPointer_PTR11), .B(_03296__PTR10), .Z(_03297__PTR11) );
  XOR2_X1 U15805 ( .A(P3_P1_InstAddrPointer_PTR12), .B(_03296__PTR11), .Z(_03297__PTR12) );
  XOR2_X1 U15806 ( .A(P3_P1_InstAddrPointer_PTR13), .B(_03296__PTR12), .Z(_03297__PTR13) );
  XOR2_X1 U15807 ( .A(P3_P1_InstAddrPointer_PTR14), .B(_03296__PTR13), .Z(_03297__PTR14) );
  XOR2_X1 U15808 ( .A(P3_P1_InstAddrPointer_PTR15), .B(_03296__PTR14), .Z(_03297__PTR15) );
  XOR2_X1 U15809 ( .A(P3_P1_InstAddrPointer_PTR16), .B(_03296__PTR15), .Z(_03297__PTR16) );
  XOR2_X1 U15810 ( .A(P3_P1_InstAddrPointer_PTR17), .B(_03296__PTR16), .Z(_03297__PTR17) );
  XOR2_X1 U15811 ( .A(P3_P1_InstAddrPointer_PTR18), .B(_03296__PTR17), .Z(_03297__PTR18) );
  XOR2_X1 U15812 ( .A(P3_P1_InstAddrPointer_PTR19), .B(_03296__PTR18), .Z(_03297__PTR19) );
  XOR2_X1 U15813 ( .A(P3_P1_InstAddrPointer_PTR20), .B(_03296__PTR19), .Z(_03297__PTR20) );
  XOR2_X1 U15814 ( .A(P3_P1_InstAddrPointer_PTR21), .B(_03296__PTR20), .Z(_03297__PTR21) );
  XOR2_X1 U15815 ( .A(P3_P1_InstAddrPointer_PTR22), .B(_03296__PTR21), .Z(_03297__PTR22) );
  XOR2_X1 U15816 ( .A(P3_P1_InstAddrPointer_PTR23), .B(_03296__PTR22), .Z(_03297__PTR23) );
  XOR2_X1 U15817 ( .A(P3_P1_InstAddrPointer_PTR24), .B(_03296__PTR23), .Z(_03297__PTR24) );
  XOR2_X1 U15818 ( .A(P3_P1_InstAddrPointer_PTR25), .B(_03296__PTR24), .Z(_03297__PTR25) );
  XOR2_X1 U15819 ( .A(P3_P1_InstAddrPointer_PTR26), .B(_03296__PTR25), .Z(_03297__PTR26) );
  XOR2_X1 U15820 ( .A(P3_P1_InstAddrPointer_PTR27), .B(_03296__PTR26), .Z(_03297__PTR27) );
  XOR2_X1 U15821 ( .A(P3_P1_InstAddrPointer_PTR28), .B(_03296__PTR27), .Z(_03297__PTR28) );
  XOR2_X1 U15822 ( .A(P3_P1_InstAddrPointer_PTR29), .B(_03296__PTR28), .Z(_03297__PTR29) );
  XOR2_X1 U15823 ( .A(P3_P1_InstAddrPointer_PTR30), .B(_03296__PTR29), .Z(_03297__PTR30) );
  XOR2_X1 U15824 ( .A(P3_P1_InstAddrPointer_PTR31), .B(_03296__PTR30), .Z(_03297__PTR31) );
  XOR2_X1 U15825 ( .A(_03299__PTR1), .B(_03298__PTR0), .Z(_03300__PTR1) );
  XOR2_X1 U15826 ( .A(_03299__PTR2), .B(_03298__PTR1), .Z(_03300__PTR2) );
  XOR2_X1 U15827 ( .A(_03299__PTR3), .B(_03298__PTR2), .Z(_03300__PTR3) );
  XOR2_X1 U15828 ( .A(_03299__PTR4), .B(_03298__PTR3), .Z(_03300__PTR4) );
  XOR2_X1 U15829 ( .A(_03299__PTR5), .B(_03298__PTR4), .Z(_03300__PTR5) );
  XOR2_X1 U15830 ( .A(_03299__PTR6), .B(_03298__PTR5), .Z(_03300__PTR6) );
  XOR2_X1 U15831 ( .A(_03299__PTR7), .B(_03298__PTR6), .Z(_03300__PTR7) );
  XOR2_X1 U15832 ( .A(_03297__PTR8), .B(_03298__PTR7), .Z(_03300__PTR8) );
  XOR2_X1 U15833 ( .A(_03297__PTR9), .B(_03298__PTR8), .Z(_03300__PTR9) );
  XOR2_X1 U15834 ( .A(_03297__PTR10), .B(_03298__PTR9), .Z(_03300__PTR10) );
  XOR2_X1 U15835 ( .A(_03297__PTR11), .B(_03298__PTR10), .Z(_03300__PTR11) );
  XOR2_X1 U15836 ( .A(_03297__PTR12), .B(_03298__PTR11), .Z(_03300__PTR12) );
  XOR2_X1 U15837 ( .A(_03297__PTR13), .B(_03298__PTR12), .Z(_03300__PTR13) );
  XOR2_X1 U15838 ( .A(_03297__PTR14), .B(_03298__PTR13), .Z(_03300__PTR14) );
  XOR2_X1 U15839 ( .A(_03297__PTR15), .B(_03298__PTR14), .Z(_03300__PTR15) );
  XOR2_X1 U15840 ( .A(_03297__PTR16), .B(_03298__PTR15), .Z(_03300__PTR16) );
  XOR2_X1 U15841 ( .A(_03297__PTR17), .B(_03298__PTR16), .Z(_03300__PTR17) );
  XOR2_X1 U15842 ( .A(_03297__PTR18), .B(_03298__PTR17), .Z(_03300__PTR18) );
  XOR2_X1 U15843 ( .A(_03297__PTR19), .B(_03298__PTR18), .Z(_03300__PTR19) );
  XOR2_X1 U15844 ( .A(_03297__PTR20), .B(_03298__PTR19), .Z(_03300__PTR20) );
  XOR2_X1 U15845 ( .A(_03297__PTR21), .B(_03298__PTR20), .Z(_03300__PTR21) );
  XOR2_X1 U15846 ( .A(_03297__PTR22), .B(_03298__PTR21), .Z(_03300__PTR22) );
  XOR2_X1 U15847 ( .A(_03297__PTR23), .B(_03298__PTR22), .Z(_03300__PTR23) );
  XOR2_X1 U15848 ( .A(_03297__PTR24), .B(_03298__PTR23), .Z(_03300__PTR24) );
  XOR2_X1 U15849 ( .A(_03297__PTR25), .B(_03298__PTR24), .Z(_03300__PTR25) );
  XOR2_X1 U15850 ( .A(_03297__PTR26), .B(_03298__PTR25), .Z(_03300__PTR26) );
  XOR2_X1 U15851 ( .A(_03297__PTR27), .B(_03298__PTR26), .Z(_03300__PTR27) );
  XOR2_X1 U15852 ( .A(_03297__PTR28), .B(_03298__PTR27), .Z(_03300__PTR28) );
  XOR2_X1 U15853 ( .A(_03297__PTR29), .B(_03298__PTR28), .Z(_03300__PTR29) );
  XOR2_X1 U15854 ( .A(_03297__PTR30), .B(_03298__PTR29), .Z(_03300__PTR30) );
  XOR2_X1 U15855 ( .A(_03297__PTR31), .B(_03298__PTR30), .Z(_03300__PTR31) );
  XOR2_X1 U15856 ( .A(_02662__PTR0), .B(_02466__PTR0), .Z(_03299__PTR0) );
  XOR2_X1 U15857 ( .A(_03297__PTR2), .B(_02466__PTR2), .Z(_03299__PTR2) );
  XOR2_X1 U15858 ( .A(_03297__PTR3), .B(_02466__PTR3), .Z(_03299__PTR3) );
  XOR2_X1 U15859 ( .A(_03297__PTR4), .B(_02466__PTR4), .Z(_03299__PTR4) );
  XOR2_X1 U15860 ( .A(_03297__PTR5), .B(_02466__PTR5), .Z(_03299__PTR5) );
  XOR2_X1 U15861 ( .A(_03297__PTR6), .B(_02466__PTR6), .Z(_03299__PTR6) );
  XOR2_X1 U15862 ( .A(_03297__PTR7), .B(_02466__PTR7), .Z(_03299__PTR7) );
  AND2_X1 U15863 ( .A1(_02662__PTR1), .A2(_02466__PTR1), .ZN(_03301__PTR1) );
  AND2_X1 U15864 ( .A1(_03297__PTR2), .A2(_02466__PTR2), .ZN(_03301__PTR2) );
  AND2_X1 U15865 ( .A1(_03297__PTR3), .A2(_02466__PTR3), .ZN(_03301__PTR3) );
  AND2_X1 U15866 ( .A1(_03297__PTR4), .A2(_02466__PTR4), .ZN(_03301__PTR4) );
  AND2_X1 U15867 ( .A1(_03297__PTR5), .A2(_02466__PTR5), .ZN(_03301__PTR5) );
  AND2_X1 U15868 ( .A1(_03297__PTR6), .A2(_02466__PTR6), .ZN(_03301__PTR6) );
  AND2_X1 U15869 ( .A1(_03297__PTR7), .A2(_02466__PTR7), .ZN(_03301__PTR7) );
  XOR2_X1 U15870 ( .A(P3_P1_InstAddrPointer_PTR2), .B(P3_P1_InstAddrPointer_PTR1), .Z(_02662__PTR34) );
  XOR2_X1 U15871 ( .A(P3_P1_InstAddrPointer_PTR3), .B(_03291__PTR1), .Z(_02662__PTR35) );
  XOR2_X1 U15872 ( .A(P3_P1_InstAddrPointer_PTR4), .B(_03291__PTR2), .Z(_02662__PTR36) );
  XOR2_X1 U15873 ( .A(P3_P1_InstAddrPointer_PTR5), .B(_03291__PTR3), .Z(_02662__PTR37) );
  XOR2_X1 U15874 ( .A(P3_P1_InstAddrPointer_PTR6), .B(_03291__PTR4), .Z(_02662__PTR38) );
  XOR2_X1 U15875 ( .A(P3_P1_InstAddrPointer_PTR7), .B(_03291__PTR5), .Z(_02662__PTR39) );
  XOR2_X1 U15876 ( .A(P3_P1_InstAddrPointer_PTR8), .B(_03291__PTR6), .Z(_02662__PTR40) );
  XOR2_X1 U15877 ( .A(P3_P1_InstAddrPointer_PTR9), .B(_03291__PTR7), .Z(_02662__PTR41) );
  XOR2_X1 U15878 ( .A(P3_P1_InstAddrPointer_PTR10), .B(_03291__PTR8), .Z(_02662__PTR42) );
  XOR2_X1 U15879 ( .A(P3_P1_InstAddrPointer_PTR11), .B(_03291__PTR9), .Z(_02662__PTR43) );
  XOR2_X1 U15880 ( .A(P3_P1_InstAddrPointer_PTR12), .B(_03291__PTR10), .Z(_02662__PTR44) );
  XOR2_X1 U15881 ( .A(P3_P1_InstAddrPointer_PTR13), .B(_03291__PTR11), .Z(_02662__PTR45) );
  XOR2_X1 U15882 ( .A(P3_P1_InstAddrPointer_PTR14), .B(_03291__PTR12), .Z(_02662__PTR46) );
  XOR2_X1 U15883 ( .A(P3_P1_InstAddrPointer_PTR15), .B(_03291__PTR13), .Z(_02662__PTR47) );
  XOR2_X1 U15884 ( .A(P3_P1_InstAddrPointer_PTR16), .B(_03291__PTR14), .Z(_02662__PTR48) );
  XOR2_X1 U15885 ( .A(P3_P1_InstAddrPointer_PTR17), .B(_03291__PTR15), .Z(_02662__PTR49) );
  XOR2_X1 U15886 ( .A(P3_P1_InstAddrPointer_PTR18), .B(_03291__PTR16), .Z(_02662__PTR50) );
  XOR2_X1 U15887 ( .A(P3_P1_InstAddrPointer_PTR19), .B(_03291__PTR17), .Z(_02662__PTR51) );
  XOR2_X1 U15888 ( .A(P3_P1_InstAddrPointer_PTR20), .B(_03291__PTR18), .Z(_02662__PTR52) );
  XOR2_X1 U15889 ( .A(P3_P1_InstAddrPointer_PTR21), .B(_03291__PTR19), .Z(_02662__PTR53) );
  XOR2_X1 U15890 ( .A(P3_P1_InstAddrPointer_PTR22), .B(_03291__PTR20), .Z(_02662__PTR54) );
  XOR2_X1 U15891 ( .A(P3_P1_InstAddrPointer_PTR23), .B(_03291__PTR21), .Z(_02662__PTR55) );
  XOR2_X1 U15892 ( .A(P3_P1_InstAddrPointer_PTR24), .B(_03291__PTR22), .Z(_02662__PTR56) );
  XOR2_X1 U15893 ( .A(P3_P1_InstAddrPointer_PTR25), .B(_03291__PTR23), .Z(_02662__PTR57) );
  XOR2_X1 U15894 ( .A(P3_P1_InstAddrPointer_PTR26), .B(_03291__PTR24), .Z(_02662__PTR58) );
  XOR2_X1 U15895 ( .A(P3_P1_InstAddrPointer_PTR27), .B(_03291__PTR25), .Z(_02662__PTR59) );
  XOR2_X1 U15896 ( .A(P3_P1_InstAddrPointer_PTR28), .B(_03291__PTR26), .Z(_02662__PTR60) );
  XOR2_X1 U15897 ( .A(P3_P1_InstAddrPointer_PTR29), .B(_03291__PTR27), .Z(_02662__PTR61) );
  XOR2_X1 U15898 ( .A(P3_P1_InstAddrPointer_PTR30), .B(_03291__PTR28), .Z(_02662__PTR62) );
  XOR2_X1 U15899 ( .A(P3_P1_InstAddrPointer_PTR31), .B(_03291__PTR29), .Z(_02662__PTR63) );
  XOR2_X1 U15900 ( .A(_03293__PTR1), .B(_03292__PTR0), .Z(_03294__PTR1) );
  XOR2_X1 U15901 ( .A(_03293__PTR2), .B(_03292__PTR1), .Z(_03294__PTR2) );
  XOR2_X1 U15902 ( .A(_03293__PTR3), .B(_03292__PTR2), .Z(_03294__PTR3) );
  XOR2_X1 U15903 ( .A(_03293__PTR4), .B(_03292__PTR3), .Z(_03294__PTR4) );
  XOR2_X1 U15904 ( .A(_03293__PTR5), .B(_03292__PTR4), .Z(_03294__PTR5) );
  XOR2_X1 U15905 ( .A(_03293__PTR6), .B(_03292__PTR5), .Z(_03294__PTR6) );
  XOR2_X1 U15906 ( .A(_03293__PTR7), .B(_03292__PTR6), .Z(_03294__PTR7) );
  XOR2_X1 U15907 ( .A(_02662__PTR40), .B(_03292__PTR7), .Z(_03294__PTR8) );
  XOR2_X1 U15908 ( .A(_02662__PTR41), .B(_03292__PTR8), .Z(_03294__PTR9) );
  XOR2_X1 U15909 ( .A(_02662__PTR42), .B(_03292__PTR9), .Z(_03294__PTR10) );
  XOR2_X1 U15910 ( .A(_02662__PTR43), .B(_03292__PTR10), .Z(_03294__PTR11) );
  XOR2_X1 U15911 ( .A(_02662__PTR44), .B(_03292__PTR11), .Z(_03294__PTR12) );
  XOR2_X1 U15912 ( .A(_02662__PTR45), .B(_03292__PTR12), .Z(_03294__PTR13) );
  XOR2_X1 U15913 ( .A(_02662__PTR46), .B(_03292__PTR13), .Z(_03294__PTR14) );
  XOR2_X1 U15914 ( .A(_02662__PTR47), .B(_03292__PTR14), .Z(_03294__PTR15) );
  XOR2_X1 U15915 ( .A(_02662__PTR48), .B(_03292__PTR15), .Z(_03294__PTR16) );
  XOR2_X1 U15916 ( .A(_02662__PTR49), .B(_03292__PTR16), .Z(_03294__PTR17) );
  XOR2_X1 U15917 ( .A(_02662__PTR50), .B(_03292__PTR17), .Z(_03294__PTR18) );
  XOR2_X1 U15918 ( .A(_02662__PTR51), .B(_03292__PTR18), .Z(_03294__PTR19) );
  XOR2_X1 U15919 ( .A(_02662__PTR52), .B(_03292__PTR19), .Z(_03294__PTR20) );
  XOR2_X1 U15920 ( .A(_02662__PTR53), .B(_03292__PTR20), .Z(_03294__PTR21) );
  XOR2_X1 U15921 ( .A(_02662__PTR54), .B(_03292__PTR21), .Z(_03294__PTR22) );
  XOR2_X1 U15922 ( .A(_02662__PTR55), .B(_03292__PTR22), .Z(_03294__PTR23) );
  XOR2_X1 U15923 ( .A(_02662__PTR56), .B(_03292__PTR23), .Z(_03294__PTR24) );
  XOR2_X1 U15924 ( .A(_02662__PTR57), .B(_03292__PTR24), .Z(_03294__PTR25) );
  XOR2_X1 U15925 ( .A(_02662__PTR58), .B(_03292__PTR25), .Z(_03294__PTR26) );
  XOR2_X1 U15926 ( .A(_02662__PTR59), .B(_03292__PTR26), .Z(_03294__PTR27) );
  XOR2_X1 U15927 ( .A(_02662__PTR60), .B(_03292__PTR27), .Z(_03294__PTR28) );
  XOR2_X1 U15928 ( .A(_02662__PTR61), .B(_03292__PTR28), .Z(_03294__PTR29) );
  XOR2_X1 U15929 ( .A(_02662__PTR62), .B(_03292__PTR29), .Z(_03294__PTR30) );
  XOR2_X1 U15930 ( .A(_02662__PTR63), .B(_03292__PTR30), .Z(_03294__PTR31) );
  XOR2_X1 U15931 ( .A(P3_P1_InstAddrPointer_PTR0), .B(_02466__PTR0), .Z(_03293__PTR0) );
  XOR2_X1 U15932 ( .A(_02662__PTR33), .B(_02466__PTR1), .Z(_03293__PTR1) );
  XOR2_X1 U15933 ( .A(_02662__PTR34), .B(_02466__PTR2), .Z(_03293__PTR2) );
  XOR2_X1 U15934 ( .A(_02662__PTR35), .B(_02466__PTR3), .Z(_03293__PTR3) );
  XOR2_X1 U15935 ( .A(_02662__PTR36), .B(_02466__PTR4), .Z(_03293__PTR4) );
  XOR2_X1 U15936 ( .A(_02662__PTR37), .B(_02466__PTR5), .Z(_03293__PTR5) );
  XOR2_X1 U15937 ( .A(_02662__PTR38), .B(_02466__PTR6), .Z(_03293__PTR6) );
  XOR2_X1 U15938 ( .A(_02662__PTR39), .B(_02466__PTR7), .Z(_03293__PTR7) );
  AND2_X1 U15939 ( .A1(P3_P1_InstAddrPointer_PTR0), .A2(_02466__PTR0), .ZN(_03292__PTR0) );
  AND2_X1 U15940 ( .A1(_02662__PTR33), .A2(_02466__PTR1), .ZN(_03295__PTR1) );
  AND2_X1 U15941 ( .A1(_02662__PTR34), .A2(_02466__PTR2), .ZN(_03295__PTR2) );
  AND2_X1 U15942 ( .A1(_02662__PTR35), .A2(_02466__PTR3), .ZN(_03295__PTR3) );
  AND2_X1 U15943 ( .A1(_02662__PTR36), .A2(_02466__PTR4), .ZN(_03295__PTR4) );
  AND2_X1 U15944 ( .A1(_02662__PTR37), .A2(_02466__PTR5), .ZN(_03295__PTR5) );
  AND2_X1 U15945 ( .A1(_02662__PTR38), .A2(_02466__PTR6), .ZN(_03295__PTR6) );
  AND2_X1 U15946 ( .A1(_02662__PTR39), .A2(_02466__PTR7), .ZN(_03295__PTR7) );
  XOR2_X1 U15947 ( .A(_02466__PTR4), .B(_03214__PTR3), .Z(_03215__PTR4) );
  XOR2_X1 U15948 ( .A(_02466__PTR6), .B(_03214__PTR5), .Z(_03215__PTR6) );
  XOR2_X1 U15949 ( .A(_02466__PTR7), .B(_03214__PTR6), .Z(_03425__PTR7) );
  XOR2_X1 U15950 ( .A(P3_P1_InstAddrPointer_PTR2), .B(_03288__PTR1), .Z(_02662__PTR2) );
  XOR2_X1 U15951 ( .A(P3_P1_InstAddrPointer_PTR3), .B(_03288__PTR2), .Z(_02662__PTR3) );
  XOR2_X1 U15952 ( .A(P3_P1_InstAddrPointer_PTR4), .B(_03288__PTR3), .Z(_02662__PTR4) );
  XOR2_X1 U15953 ( .A(P3_P1_InstAddrPointer_PTR5), .B(_03288__PTR4), .Z(_02662__PTR5) );
  XOR2_X1 U15954 ( .A(P3_P1_InstAddrPointer_PTR6), .B(_03288__PTR5), .Z(_02662__PTR6) );
  XOR2_X1 U15955 ( .A(P3_P1_InstAddrPointer_PTR7), .B(_03288__PTR6), .Z(_02662__PTR7) );
  XOR2_X1 U15956 ( .A(P3_P1_InstAddrPointer_PTR8), .B(_03288__PTR7), .Z(_02662__PTR8) );
  XOR2_X1 U15957 ( .A(P3_P1_InstAddrPointer_PTR9), .B(_03288__PTR8), .Z(_02662__PTR9) );
  XOR2_X1 U15958 ( .A(P3_P1_InstAddrPointer_PTR10), .B(_03288__PTR9), .Z(_02662__PTR10) );
  XOR2_X1 U15959 ( .A(P3_P1_InstAddrPointer_PTR11), .B(_03288__PTR10), .Z(_02662__PTR11) );
  XOR2_X1 U15960 ( .A(P3_P1_InstAddrPointer_PTR12), .B(_03288__PTR11), .Z(_02662__PTR12) );
  XOR2_X1 U15961 ( .A(P3_P1_InstAddrPointer_PTR13), .B(_03288__PTR12), .Z(_02662__PTR13) );
  XOR2_X1 U15962 ( .A(P3_P1_InstAddrPointer_PTR14), .B(_03288__PTR13), .Z(_02662__PTR14) );
  XOR2_X1 U15963 ( .A(P3_P1_InstAddrPointer_PTR15), .B(_03288__PTR14), .Z(_02662__PTR15) );
  XOR2_X1 U15964 ( .A(P3_P1_InstAddrPointer_PTR16), .B(_03288__PTR15), .Z(_02662__PTR16) );
  XOR2_X1 U15965 ( .A(P3_P1_InstAddrPointer_PTR17), .B(_03288__PTR16), .Z(_02662__PTR17) );
  XOR2_X1 U15966 ( .A(P3_P1_InstAddrPointer_PTR18), .B(_03288__PTR17), .Z(_02662__PTR18) );
  XOR2_X1 U15967 ( .A(P3_P1_InstAddrPointer_PTR19), .B(_03288__PTR18), .Z(_02662__PTR19) );
  XOR2_X1 U15968 ( .A(P3_P1_InstAddrPointer_PTR20), .B(_03288__PTR19), .Z(_02662__PTR20) );
  XOR2_X1 U15969 ( .A(P3_P1_InstAddrPointer_PTR21), .B(_03288__PTR20), .Z(_02662__PTR21) );
  XOR2_X1 U15970 ( .A(P3_P1_InstAddrPointer_PTR22), .B(_03288__PTR21), .Z(_02662__PTR22) );
  XOR2_X1 U15971 ( .A(P3_P1_InstAddrPointer_PTR23), .B(_03288__PTR22), .Z(_02662__PTR23) );
  XOR2_X1 U15972 ( .A(P3_P1_InstAddrPointer_PTR24), .B(_03288__PTR23), .Z(_02662__PTR24) );
  XOR2_X1 U15973 ( .A(P3_P1_InstAddrPointer_PTR25), .B(_03288__PTR24), .Z(_02662__PTR25) );
  XOR2_X1 U15974 ( .A(P3_P1_InstAddrPointer_PTR26), .B(_03288__PTR25), .Z(_02662__PTR26) );
  XOR2_X1 U15975 ( .A(P3_P1_InstAddrPointer_PTR27), .B(_03288__PTR26), .Z(_02662__PTR27) );
  XOR2_X1 U15976 ( .A(P3_P1_InstAddrPointer_PTR28), .B(_03288__PTR27), .Z(_02662__PTR28) );
  XOR2_X1 U15977 ( .A(P3_P1_InstAddrPointer_PTR29), .B(_03288__PTR28), .Z(_02662__PTR29) );
  XOR2_X1 U15978 ( .A(P3_P1_InstAddrPointer_PTR30), .B(_03288__PTR29), .Z(_02662__PTR30) );
  XOR2_X1 U15979 ( .A(P3_P1_InstAddrPointer_PTR31), .B(_03288__PTR30), .Z(_02662__PTR31) );
  XOR2_X1 U15980 ( .A(_03299__PTR1), .B(_03427__PTR0), .Z(_03429__PTR1) );
  XOR2_X1 U15981 ( .A(_03428__PTR2), .B(_03427__PTR1), .Z(_03429__PTR2) );
  XOR2_X1 U15982 ( .A(_03428__PTR3), .B(_03427__PTR2), .Z(_03429__PTR3) );
  XOR2_X1 U15983 ( .A(_03428__PTR4), .B(_03427__PTR3), .Z(_03429__PTR4) );
  XOR2_X1 U15984 ( .A(_03428__PTR5), .B(_03427__PTR4), .Z(_03429__PTR5) );
  XOR2_X1 U15985 ( .A(_03428__PTR6), .B(_03427__PTR5), .Z(_03429__PTR6) );
  XOR2_X1 U15986 ( .A(_03428__PTR7), .B(_03427__PTR6), .Z(_03429__PTR7) );
  XOR2_X1 U15987 ( .A(_03428__PTR8), .B(_03427__PTR7), .Z(_03429__PTR8) );
  XOR2_X1 U15988 ( .A(_03428__PTR9), .B(_03427__PTR8), .Z(_03429__PTR9) );
  XOR2_X1 U15989 ( .A(_03428__PTR10), .B(_03427__PTR9), .Z(_03429__PTR10) );
  XOR2_X1 U15990 ( .A(_03428__PTR11), .B(_03427__PTR10), .Z(_03429__PTR11) );
  XOR2_X1 U15991 ( .A(_03428__PTR12), .B(_03427__PTR11), .Z(_03429__PTR12) );
  XOR2_X1 U15992 ( .A(_03428__PTR13), .B(_03427__PTR12), .Z(_03429__PTR13) );
  XOR2_X1 U15993 ( .A(_03428__PTR14), .B(_03427__PTR13), .Z(_03429__PTR14) );
  XOR2_X1 U15994 ( .A(_03428__PTR15), .B(_03427__PTR14), .Z(_03429__PTR15) );
  XOR2_X1 U15995 ( .A(_03428__PTR16), .B(_03427__PTR15), .Z(_03429__PTR16) );
  XOR2_X1 U15996 ( .A(_03428__PTR17), .B(_03427__PTR16), .Z(_03429__PTR17) );
  XOR2_X1 U15997 ( .A(_03428__PTR18), .B(_03427__PTR17), .Z(_03429__PTR18) );
  XOR2_X1 U15998 ( .A(_03428__PTR19), .B(_03427__PTR18), .Z(_03429__PTR19) );
  XOR2_X1 U15999 ( .A(_03428__PTR20), .B(_03427__PTR19), .Z(_03429__PTR20) );
  XOR2_X1 U16000 ( .A(_03428__PTR21), .B(_03427__PTR20), .Z(_03429__PTR21) );
  XOR2_X1 U16001 ( .A(_03428__PTR22), .B(_03427__PTR21), .Z(_03429__PTR22) );
  XOR2_X1 U16002 ( .A(_03428__PTR23), .B(_03427__PTR22), .Z(_03429__PTR23) );
  XOR2_X1 U16003 ( .A(_03428__PTR24), .B(_03427__PTR23), .Z(_03429__PTR24) );
  XOR2_X1 U16004 ( .A(_03428__PTR25), .B(_03427__PTR24), .Z(_03429__PTR25) );
  XOR2_X1 U16005 ( .A(_03428__PTR26), .B(_03427__PTR25), .Z(_03429__PTR26) );
  XOR2_X1 U16006 ( .A(_03428__PTR27), .B(_03427__PTR26), .Z(_03429__PTR27) );
  XOR2_X1 U16007 ( .A(_03428__PTR28), .B(_03427__PTR27), .Z(_03429__PTR28) );
  XOR2_X1 U16008 ( .A(_03428__PTR29), .B(_03427__PTR28), .Z(_03429__PTR29) );
  XOR2_X1 U16009 ( .A(_03428__PTR30), .B(_03427__PTR29), .Z(_03429__PTR30) );
  XOR2_X1 U16010 ( .A(_03428__PTR32), .B(_03427__PTR30), .Z(_03429__PTR31) );
  XOR2_X1 U16011 ( .A(_02662__PTR1), .B(_02466__PTR1), .Z(_03299__PTR1) );
  XOR2_X1 U16012 ( .A(_02662__PTR2), .B(_02466__PTR2), .Z(_03428__PTR2) );
  XOR2_X1 U16013 ( .A(_02662__PTR3), .B(_02466__PTR3), .Z(_03428__PTR3) );
  XOR2_X1 U16014 ( .A(_02662__PTR4), .B(_03426__PTR4), .Z(_03428__PTR4) );
  XOR2_X1 U16015 ( .A(_02662__PTR5), .B(_03426__PTR5), .Z(_03428__PTR5) );
  XOR2_X1 U16016 ( .A(_02662__PTR6), .B(_03426__PTR6), .Z(_03428__PTR6) );
  XOR2_X1 U16017 ( .A(_02662__PTR7), .B(_03426__PTR7), .Z(_03428__PTR7) );
  XOR2_X1 U16018 ( .A(_02662__PTR8), .B(_03424__PTR8), .Z(_03428__PTR8) );
  XOR2_X1 U16019 ( .A(_02662__PTR9), .B(_03424__PTR8), .Z(_03428__PTR9) );
  XOR2_X1 U16020 ( .A(_02662__PTR10), .B(_03424__PTR8), .Z(_03428__PTR10) );
  XOR2_X1 U16021 ( .A(_02662__PTR11), .B(_03424__PTR8), .Z(_03428__PTR11) );
  XOR2_X1 U16022 ( .A(_02662__PTR12), .B(_03424__PTR8), .Z(_03428__PTR12) );
  XOR2_X1 U16023 ( .A(_02662__PTR13), .B(_03424__PTR8), .Z(_03428__PTR13) );
  XOR2_X1 U16024 ( .A(_02662__PTR14), .B(_03424__PTR8), .Z(_03428__PTR14) );
  XOR2_X1 U16025 ( .A(_02662__PTR15), .B(_03424__PTR8), .Z(_03428__PTR15) );
  XOR2_X1 U16026 ( .A(_02662__PTR16), .B(_03424__PTR8), .Z(_03428__PTR16) );
  XOR2_X1 U16027 ( .A(_02662__PTR17), .B(_03424__PTR8), .Z(_03428__PTR17) );
  XOR2_X1 U16028 ( .A(_02662__PTR18), .B(_03424__PTR8), .Z(_03428__PTR18) );
  XOR2_X1 U16029 ( .A(_02662__PTR19), .B(_03424__PTR8), .Z(_03428__PTR19) );
  XOR2_X1 U16030 ( .A(_02662__PTR20), .B(_03424__PTR8), .Z(_03428__PTR20) );
  XOR2_X1 U16031 ( .A(_02662__PTR21), .B(_03424__PTR8), .Z(_03428__PTR21) );
  XOR2_X1 U16032 ( .A(_02662__PTR22), .B(_03424__PTR8), .Z(_03428__PTR22) );
  XOR2_X1 U16033 ( .A(_02662__PTR23), .B(_03424__PTR8), .Z(_03428__PTR23) );
  XOR2_X1 U16034 ( .A(_02662__PTR24), .B(_03424__PTR8), .Z(_03428__PTR24) );
  XOR2_X1 U16035 ( .A(_02662__PTR25), .B(_03424__PTR8), .Z(_03428__PTR25) );
  XOR2_X1 U16036 ( .A(_02662__PTR26), .B(_03424__PTR8), .Z(_03428__PTR26) );
  XOR2_X1 U16037 ( .A(_02662__PTR27), .B(_03424__PTR8), .Z(_03428__PTR27) );
  XOR2_X1 U16038 ( .A(_02662__PTR28), .B(_03424__PTR8), .Z(_03428__PTR28) );
  XOR2_X1 U16039 ( .A(_02662__PTR29), .B(_03424__PTR8), .Z(_03428__PTR29) );
  XOR2_X1 U16040 ( .A(_02662__PTR30), .B(_03424__PTR8), .Z(_03428__PTR30) );
  XOR2_X1 U16041 ( .A(_02662__PTR31), .B(_03424__PTR8), .Z(_03428__PTR32) );
  AND2_X1 U16042 ( .A1(_02662__PTR0), .A2(_02466__PTR0), .ZN(_03298__PTR0) );
  AND2_X1 U16043 ( .A1(_02662__PTR2), .A2(_02466__PTR2), .ZN(_03430__PTR2) );
  AND2_X1 U16044 ( .A1(_02662__PTR3), .A2(_02466__PTR3), .ZN(_03430__PTR3) );
  AND2_X1 U16045 ( .A1(_02662__PTR4), .A2(_03426__PTR4), .ZN(_03430__PTR4) );
  AND2_X1 U16046 ( .A1(_02662__PTR5), .A2(_03426__PTR5), .ZN(_03430__PTR5) );
  AND2_X1 U16047 ( .A1(_02662__PTR6), .A2(_03426__PTR6), .ZN(_03430__PTR6) );
  AND2_X1 U16048 ( .A1(_02662__PTR7), .A2(_03426__PTR7), .ZN(_03430__PTR7) );
  AND2_X1 U16049 ( .A1(_02662__PTR8), .A2(_03424__PTR8), .ZN(_03430__PTR8) );
  AND2_X1 U16050 ( .A1(_02662__PTR9), .A2(_03424__PTR8), .ZN(_03430__PTR9) );
  AND2_X1 U16051 ( .A1(_02662__PTR10), .A2(_03424__PTR8), .ZN(_03430__PTR10) );
  AND2_X1 U16052 ( .A1(_02662__PTR11), .A2(_03424__PTR8), .ZN(_03430__PTR11) );
  AND2_X1 U16053 ( .A1(_02662__PTR12), .A2(_03424__PTR8), .ZN(_03430__PTR12) );
  AND2_X1 U16054 ( .A1(_02662__PTR13), .A2(_03424__PTR8), .ZN(_03430__PTR13) );
  AND2_X1 U16055 ( .A1(_02662__PTR14), .A2(_03424__PTR8), .ZN(_03430__PTR14) );
  AND2_X1 U16056 ( .A1(_02662__PTR15), .A2(_03424__PTR8), .ZN(_03430__PTR15) );
  AND2_X1 U16057 ( .A1(_02662__PTR16), .A2(_03424__PTR8), .ZN(_03430__PTR16) );
  AND2_X1 U16058 ( .A1(_02662__PTR17), .A2(_03424__PTR8), .ZN(_03430__PTR17) );
  AND2_X1 U16059 ( .A1(_02662__PTR18), .A2(_03424__PTR8), .ZN(_03430__PTR18) );
  AND2_X1 U16060 ( .A1(_02662__PTR19), .A2(_03424__PTR8), .ZN(_03430__PTR19) );
  AND2_X1 U16061 ( .A1(_02662__PTR20), .A2(_03424__PTR8), .ZN(_03430__PTR20) );
  AND2_X1 U16062 ( .A1(_02662__PTR21), .A2(_03424__PTR8), .ZN(_03430__PTR21) );
  AND2_X1 U16063 ( .A1(_02662__PTR22), .A2(_03424__PTR8), .ZN(_03430__PTR22) );
  AND2_X1 U16064 ( .A1(_02662__PTR23), .A2(_03424__PTR8), .ZN(_03430__PTR23) );
  AND2_X1 U16065 ( .A1(_02662__PTR24), .A2(_03424__PTR8), .ZN(_03430__PTR24) );
  AND2_X1 U16066 ( .A1(_02662__PTR25), .A2(_03424__PTR8), .ZN(_03430__PTR25) );
  AND2_X1 U16067 ( .A1(_02662__PTR26), .A2(_03424__PTR8), .ZN(_03430__PTR26) );
  AND2_X1 U16068 ( .A1(_02662__PTR27), .A2(_03424__PTR8), .ZN(_03430__PTR27) );
  AND2_X1 U16069 ( .A1(_02662__PTR28), .A2(_03424__PTR8), .ZN(_03430__PTR28) );
  AND2_X1 U16070 ( .A1(_02662__PTR29), .A2(_03424__PTR8), .ZN(_03430__PTR29) );
  AND2_X1 U16071 ( .A1(_02662__PTR30), .A2(_03424__PTR8), .ZN(_03430__PTR30) );
  XOR2_X1 U16072 ( .A(_02466__PTR5), .B(_03214__PTR4), .Z(_03215__PTR5) );
  XOR2_X1 U16073 ( .A(P3_P1_InstQueueRd_Addr_PTR2), .B(_03240__PTR1), .Z(_02465__PTR5) );
  XOR2_X1 U16074 ( .A(P3_P1_InstQueueRd_Addr_PTR3), .B(_03240__PTR2), .Z(_02465__PTR6) );
  XOR2_X1 U16075 ( .A(P3_P1_InstQueueRd_Addr_PTR4), .B(_03240__PTR3), .Z(_03290__PTR4) );
  XOR2_X1 U16076 ( .A(P3_P1_PhyAddrPointer_PTR2), .B(P3_P1_PhyAddrPointer_PTR1), .Z(_02473__PTR130) );
  XOR2_X1 U16077 ( .A(P3_P1_PhyAddrPointer_PTR3), .B(_03287__PTR1), .Z(_02473__PTR131) );
  XOR2_X1 U16078 ( .A(P3_P1_PhyAddrPointer_PTR4), .B(_03287__PTR2), .Z(_02473__PTR132) );
  XOR2_X1 U16079 ( .A(P3_P1_PhyAddrPointer_PTR5), .B(_03287__PTR3), .Z(_02473__PTR133) );
  XOR2_X1 U16080 ( .A(P3_P1_PhyAddrPointer_PTR6), .B(_03287__PTR4), .Z(_02473__PTR134) );
  XOR2_X1 U16081 ( .A(P3_P1_PhyAddrPointer_PTR7), .B(_03287__PTR5), .Z(_02473__PTR135) );
  XOR2_X1 U16082 ( .A(P3_P1_PhyAddrPointer_PTR8), .B(_03287__PTR6), .Z(_02473__PTR136) );
  XOR2_X1 U16083 ( .A(P3_P1_PhyAddrPointer_PTR9), .B(_03287__PTR7), .Z(_02473__PTR137) );
  XOR2_X1 U16084 ( .A(P3_P1_PhyAddrPointer_PTR10), .B(_03287__PTR8), .Z(_02473__PTR138) );
  XOR2_X1 U16085 ( .A(P3_P1_PhyAddrPointer_PTR11), .B(_03287__PTR9), .Z(_02473__PTR139) );
  XOR2_X1 U16086 ( .A(P3_P1_PhyAddrPointer_PTR12), .B(_03287__PTR10), .Z(_02473__PTR140) );
  XOR2_X1 U16087 ( .A(P3_P1_PhyAddrPointer_PTR13), .B(_03287__PTR11), .Z(_02473__PTR141) );
  XOR2_X1 U16088 ( .A(P3_P1_PhyAddrPointer_PTR14), .B(_03287__PTR12), .Z(_02473__PTR142) );
  XOR2_X1 U16089 ( .A(P3_P1_PhyAddrPointer_PTR15), .B(_03287__PTR13), .Z(_02473__PTR143) );
  XOR2_X1 U16090 ( .A(P3_P1_PhyAddrPointer_PTR16), .B(_03287__PTR14), .Z(_02473__PTR144) );
  XOR2_X1 U16091 ( .A(P3_P1_PhyAddrPointer_PTR17), .B(_03287__PTR15), .Z(_02473__PTR145) );
  XOR2_X1 U16092 ( .A(P3_P1_PhyAddrPointer_PTR18), .B(_03287__PTR16), .Z(_02473__PTR146) );
  XOR2_X1 U16093 ( .A(P3_P1_PhyAddrPointer_PTR19), .B(_03287__PTR17), .Z(_02473__PTR147) );
  XOR2_X1 U16094 ( .A(P3_P1_PhyAddrPointer_PTR20), .B(_03287__PTR18), .Z(_02473__PTR148) );
  XOR2_X1 U16095 ( .A(P3_P1_PhyAddrPointer_PTR21), .B(_03287__PTR19), .Z(_02473__PTR149) );
  XOR2_X1 U16096 ( .A(P3_P1_PhyAddrPointer_PTR22), .B(_03287__PTR20), .Z(_02473__PTR150) );
  XOR2_X1 U16097 ( .A(P3_P1_PhyAddrPointer_PTR23), .B(_03287__PTR21), .Z(_02473__PTR151) );
  XOR2_X1 U16098 ( .A(P3_P1_PhyAddrPointer_PTR24), .B(_03287__PTR22), .Z(_02473__PTR152) );
  XOR2_X1 U16099 ( .A(P3_P1_PhyAddrPointer_PTR25), .B(_03287__PTR23), .Z(_02473__PTR153) );
  XOR2_X1 U16100 ( .A(P3_P1_PhyAddrPointer_PTR26), .B(_03287__PTR24), .Z(_02473__PTR154) );
  XOR2_X1 U16101 ( .A(P3_P1_PhyAddrPointer_PTR27), .B(_03287__PTR25), .Z(_02473__PTR155) );
  XOR2_X1 U16102 ( .A(P3_P1_PhyAddrPointer_PTR28), .B(_03287__PTR26), .Z(_02473__PTR156) );
  XOR2_X1 U16103 ( .A(P3_P1_PhyAddrPointer_PTR29), .B(_03287__PTR27), .Z(_02473__PTR157) );
  XOR2_X1 U16104 ( .A(P3_P1_PhyAddrPointer_PTR30), .B(_03287__PTR28), .Z(_02473__PTR158) );
  XOR2_X1 U16105 ( .A(P3_P1_PhyAddrPointer_PTR31), .B(_03287__PTR29), .Z(_02473__PTR159) );
  XOR2_X1 U16106 ( .A(P3_P1_PhyAddrPointer_PTR1), .B(_03205__PTR0), .Z(_03436__PTR1) );
  XOR2_X1 U16107 ( .A(_03205__PTR2), .B(_03435__PTR1), .Z(_03436__PTR2) );
  XOR2_X1 U16108 ( .A(_03205__PTR3), .B(_03435__PTR2), .Z(_03436__PTR3) );
  XOR2_X1 U16109 ( .A(_03205__PTR4), .B(_03435__PTR3), .Z(_03436__PTR4) );
  XOR2_X1 U16110 ( .A(_03205__PTR5), .B(_03435__PTR4), .Z(_03436__PTR5) );
  XOR2_X1 U16111 ( .A(_03205__PTR6), .B(_03435__PTR5), .Z(_03436__PTR6) );
  XOR2_X1 U16112 ( .A(_03205__PTR7), .B(_03435__PTR6), .Z(_03436__PTR7) );
  XOR2_X1 U16113 ( .A(_03205__PTR8), .B(_03435__PTR7), .Z(_03436__PTR8) );
  XOR2_X1 U16114 ( .A(_03205__PTR9), .B(_03435__PTR8), .Z(_03436__PTR9) );
  XOR2_X1 U16115 ( .A(_03205__PTR10), .B(_03435__PTR9), .Z(_03436__PTR10) );
  XOR2_X1 U16116 ( .A(_03205__PTR11), .B(_03435__PTR10), .Z(_03436__PTR11) );
  XOR2_X1 U16117 ( .A(_03205__PTR12), .B(_03435__PTR11), .Z(_03436__PTR12) );
  XOR2_X1 U16118 ( .A(_03205__PTR13), .B(_03435__PTR12), .Z(_03436__PTR13) );
  XOR2_X1 U16119 ( .A(_03205__PTR14), .B(_03435__PTR13), .Z(_03436__PTR14) );
  XOR2_X1 U16120 ( .A(_03205__PTR15), .B(_03435__PTR14), .Z(_03436__PTR15) );
  XOR2_X1 U16121 ( .A(_03205__PTR16), .B(_03435__PTR15), .Z(_03436__PTR16) );
  XOR2_X1 U16122 ( .A(_03205__PTR17), .B(_03435__PTR16), .Z(_03436__PTR17) );
  XOR2_X1 U16123 ( .A(_03205__PTR18), .B(_03435__PTR17), .Z(_03436__PTR18) );
  XOR2_X1 U16124 ( .A(_03205__PTR19), .B(_03435__PTR18), .Z(_03436__PTR19) );
  XOR2_X1 U16125 ( .A(_03205__PTR20), .B(_03435__PTR19), .Z(_03436__PTR20) );
  XOR2_X1 U16126 ( .A(_03205__PTR21), .B(_03435__PTR20), .Z(_03436__PTR21) );
  XOR2_X1 U16127 ( .A(_03205__PTR22), .B(_03435__PTR21), .Z(_03436__PTR22) );
  XOR2_X1 U16128 ( .A(_03205__PTR23), .B(_03435__PTR22), .Z(_03436__PTR23) );
  XOR2_X1 U16129 ( .A(_03205__PTR24), .B(_03435__PTR23), .Z(_03436__PTR24) );
  XOR2_X1 U16130 ( .A(_03205__PTR25), .B(_03435__PTR24), .Z(_03436__PTR25) );
  XOR2_X1 U16131 ( .A(_03205__PTR26), .B(_03435__PTR25), .Z(_03436__PTR26) );
  XOR2_X1 U16132 ( .A(_03205__PTR27), .B(_03435__PTR26), .Z(_03436__PTR27) );
  XOR2_X1 U16133 ( .A(_03205__PTR28), .B(_03435__PTR27), .Z(_03436__PTR28) );
  XOR2_X1 U16134 ( .A(_03205__PTR29), .B(_03435__PTR28), .Z(_03436__PTR29) );
  XOR2_X1 U16135 ( .A(_03205__PTR30), .B(_03435__PTR29), .Z(_03436__PTR30) );
  XOR2_X1 U16136 ( .A(_03203__PTR31), .B(_03435__PTR30), .Z(_03436__PTR31) );
  XOR2_X1 U16137 ( .A(P3_P1_PhyAddrPointer_PTR3), .B(P3_P1_PhyAddrPointer_PTR2), .Z(_03286__PTR1) );
  XOR2_X1 U16138 ( .A(P3_P1_PhyAddrPointer_PTR4), .B(_03284__PTR1), .Z(_03286__PTR2) );
  XOR2_X1 U16139 ( .A(P3_P1_PhyAddrPointer_PTR5), .B(_03284__PTR2), .Z(_03286__PTR3) );
  XOR2_X1 U16140 ( .A(P3_P1_PhyAddrPointer_PTR6), .B(_03284__PTR3), .Z(_03286__PTR4) );
  XOR2_X1 U16141 ( .A(P3_P1_PhyAddrPointer_PTR7), .B(_03284__PTR4), .Z(_03286__PTR5) );
  XOR2_X1 U16142 ( .A(P3_P1_PhyAddrPointer_PTR8), .B(_03284__PTR5), .Z(_03286__PTR6) );
  XOR2_X1 U16143 ( .A(P3_P1_PhyAddrPointer_PTR9), .B(_03284__PTR6), .Z(_03286__PTR7) );
  XOR2_X1 U16144 ( .A(P3_P1_PhyAddrPointer_PTR10), .B(_03284__PTR7), .Z(_03286__PTR8) );
  XOR2_X1 U16145 ( .A(P3_P1_PhyAddrPointer_PTR11), .B(_03284__PTR8), .Z(_03286__PTR9) );
  XOR2_X1 U16146 ( .A(P3_P1_PhyAddrPointer_PTR12), .B(_03284__PTR9), .Z(_03286__PTR10) );
  XOR2_X1 U16147 ( .A(P3_P1_PhyAddrPointer_PTR13), .B(_03284__PTR10), .Z(_03286__PTR11) );
  XOR2_X1 U16148 ( .A(P3_P1_PhyAddrPointer_PTR14), .B(_03284__PTR11), .Z(_03286__PTR12) );
  XOR2_X1 U16149 ( .A(P3_P1_PhyAddrPointer_PTR15), .B(_03284__PTR12), .Z(_03286__PTR13) );
  XOR2_X1 U16150 ( .A(P3_P1_PhyAddrPointer_PTR16), .B(_03284__PTR13), .Z(_03286__PTR14) );
  XOR2_X1 U16151 ( .A(P3_P1_PhyAddrPointer_PTR17), .B(_03284__PTR14), .Z(_03286__PTR15) );
  XOR2_X1 U16152 ( .A(P3_P1_PhyAddrPointer_PTR18), .B(_03284__PTR15), .Z(_03286__PTR16) );
  XOR2_X1 U16153 ( .A(P3_P1_PhyAddrPointer_PTR19), .B(_03284__PTR16), .Z(_03286__PTR17) );
  XOR2_X1 U16154 ( .A(P3_P1_PhyAddrPointer_PTR20), .B(_03284__PTR17), .Z(_03286__PTR18) );
  XOR2_X1 U16155 ( .A(P3_P1_PhyAddrPointer_PTR21), .B(_03284__PTR18), .Z(_03286__PTR19) );
  XOR2_X1 U16156 ( .A(P3_P1_PhyAddrPointer_PTR22), .B(_03284__PTR19), .Z(_03286__PTR20) );
  XOR2_X1 U16157 ( .A(P3_P1_PhyAddrPointer_PTR23), .B(_03284__PTR20), .Z(_03286__PTR21) );
  XOR2_X1 U16158 ( .A(P3_P1_PhyAddrPointer_PTR24), .B(_03284__PTR21), .Z(_03286__PTR22) );
  XOR2_X1 U16159 ( .A(P3_P1_PhyAddrPointer_PTR25), .B(_03284__PTR22), .Z(_03286__PTR23) );
  XOR2_X1 U16160 ( .A(P3_P1_PhyAddrPointer_PTR26), .B(_03284__PTR23), .Z(_03286__PTR24) );
  XOR2_X1 U16161 ( .A(P3_P1_PhyAddrPointer_PTR27), .B(_03284__PTR24), .Z(_03286__PTR25) );
  XOR2_X1 U16162 ( .A(P3_P1_PhyAddrPointer_PTR28), .B(_03284__PTR25), .Z(_03286__PTR26) );
  XOR2_X1 U16163 ( .A(P3_P1_PhyAddrPointer_PTR29), .B(_03284__PTR26), .Z(_03286__PTR27) );
  XOR2_X1 U16164 ( .A(P3_P1_PhyAddrPointer_PTR30), .B(_03284__PTR27), .Z(_03286__PTR28) );
  XOR2_X1 U16165 ( .A(P3_P1_PhyAddrPointer_PTR31), .B(_03284__PTR28), .Z(_03286__PTR29) );
  XOR2_X1 U16166 ( .A(P3_P1_InstQueueWr_Addr_PTR1), .B(P3_P1_InstQueueWr_Addr_PTR0), .Z(_02418__PTR1) );
  XOR2_X1 U16167 ( .A(P3_P1_InstQueueWr_Addr_PTR2), .B(_03269__PTR1), .Z(_02418__PTR2) );
  XOR2_X1 U16168 ( .A(P3_P1_InstQueueWr_Addr_PTR3), .B(_03269__PTR2), .Z(_02418__PTR3) );
  XOR2_X1 U16169 ( .A(_02418__PTR1), .B(_02418__PTR0), .Z(_02420__PTR1) );
  XOR2_X1 U16170 ( .A(_02418__PTR2), .B(_03270__PTR1), .Z(_02420__PTR2) );
  XOR2_X1 U16171 ( .A(_02418__PTR3), .B(_03270__PTR2), .Z(_02420__PTR3) );
  XOR2_X1 U16172 ( .A(_02420__PTR1), .B(P3_P1_InstQueueWr_Addr_PTR0), .Z(_02422__PTR1) );
  XOR2_X1 U16173 ( .A(_02420__PTR2), .B(_03275__PTR1), .Z(_02422__PTR2) );
  XOR2_X1 U16174 ( .A(_02420__PTR3), .B(_03275__PTR2), .Z(_02422__PTR3) );
  XOR2_X1 U16175 ( .A(_02422__PTR1), .B(_02418__PTR0), .Z(_03281__PTR1) );
  XOR2_X1 U16176 ( .A(_02422__PTR2), .B(_03280__PTR1), .Z(_03281__PTR2) );
  XOR2_X1 U16177 ( .A(_02422__PTR3), .B(_03280__PTR2), .Z(_03281__PTR3) );
  XOR2_X1 U16178 ( .A(buf2_PTR25), .B(_03277__PTR0), .Z(_03279__PTR1) );
  XOR2_X1 U16179 ( .A(buf2_PTR26), .B(_03277__PTR1), .Z(_03279__PTR2) );
  XOR2_X1 U16180 ( .A(buf2_PTR27), .B(_03277__PTR2), .Z(_03279__PTR3) );
  XOR2_X1 U16181 ( .A(buf2_PTR28), .B(_03277__PTR3), .Z(_03279__PTR4) );
  XOR2_X1 U16182 ( .A(buf2_PTR29), .B(_03277__PTR4), .Z(_03279__PTR5) );
  XOR2_X1 U16183 ( .A(buf2_PTR30), .B(_03277__PTR5), .Z(_03279__PTR6) );
  XOR2_X1 U16184 ( .A(buf2_PTR31), .B(_03277__PTR6), .Z(_03279__PTR7) );
  XOR2_X1 U16185 ( .A(_03276_), .B(buf2_PTR24), .Z(_03278__PTR0) );
  AND2_X1 U16186 ( .A1(_03276_), .A2(buf2_PTR24), .ZN(_03277__PTR0) );
  XOR2_X1 U16187 ( .A(buf2_PTR17), .B(_03272__PTR0), .Z(_03274__PTR1) );
  XOR2_X1 U16188 ( .A(buf2_PTR18), .B(_03272__PTR1), .Z(_03274__PTR2) );
  XOR2_X1 U16189 ( .A(buf2_PTR19), .B(_03272__PTR2), .Z(_03274__PTR3) );
  XOR2_X1 U16190 ( .A(buf2_PTR20), .B(_03272__PTR3), .Z(_03274__PTR4) );
  XOR2_X1 U16191 ( .A(buf2_PTR21), .B(_03272__PTR4), .Z(_03274__PTR5) );
  XOR2_X1 U16192 ( .A(buf2_PTR22), .B(_03272__PTR5), .Z(_03274__PTR6) );
  XOR2_X1 U16193 ( .A(buf2_PTR23), .B(_03272__PTR6), .Z(_03274__PTR7) );
  XOR2_X1 U16194 ( .A(_03271_), .B(buf2_PTR16), .Z(_03273__PTR0) );
  AND2_X1 U16195 ( .A1(_03271_), .A2(buf2_PTR16), .ZN(_03272__PTR0) );
  XOR2_X1 U16196 ( .A(P3_rEIP_PTR2), .B(_03268__PTR0), .Z(_02461__PTR193) );
  XOR2_X1 U16197 ( .A(P3_rEIP_PTR3), .B(_03268__PTR1), .Z(_02461__PTR194) );
  XOR2_X1 U16198 ( .A(P3_rEIP_PTR4), .B(_03268__PTR2), .Z(_02461__PTR195) );
  XOR2_X1 U16199 ( .A(P3_rEIP_PTR5), .B(_03268__PTR3), .Z(_02461__PTR196) );
  XOR2_X1 U16200 ( .A(P3_rEIP_PTR6), .B(_03268__PTR4), .Z(_02461__PTR197) );
  XOR2_X1 U16201 ( .A(P3_rEIP_PTR7), .B(_03268__PTR5), .Z(_02461__PTR198) );
  XOR2_X1 U16202 ( .A(P3_rEIP_PTR8), .B(_03268__PTR6), .Z(_02461__PTR199) );
  XOR2_X1 U16203 ( .A(P3_rEIP_PTR9), .B(_03268__PTR7), .Z(_02461__PTR200) );
  XOR2_X1 U16204 ( .A(P3_rEIP_PTR10), .B(_03268__PTR8), .Z(_02461__PTR201) );
  XOR2_X1 U16205 ( .A(P3_rEIP_PTR11), .B(_03268__PTR9), .Z(_02461__PTR202) );
  XOR2_X1 U16206 ( .A(P3_rEIP_PTR12), .B(_03268__PTR10), .Z(_02461__PTR203) );
  XOR2_X1 U16207 ( .A(P3_rEIP_PTR13), .B(_03268__PTR11), .Z(_02461__PTR204) );
  XOR2_X1 U16208 ( .A(P3_rEIP_PTR14), .B(_03268__PTR12), .Z(_02461__PTR205) );
  XOR2_X1 U16209 ( .A(P3_rEIP_PTR15), .B(_03268__PTR13), .Z(_02461__PTR206) );
  XOR2_X1 U16210 ( .A(P3_rEIP_PTR16), .B(_03268__PTR14), .Z(_02461__PTR207) );
  XOR2_X1 U16211 ( .A(P3_rEIP_PTR17), .B(_03268__PTR15), .Z(_02461__PTR208) );
  XOR2_X1 U16212 ( .A(P3_rEIP_PTR18), .B(_03268__PTR16), .Z(_02461__PTR209) );
  XOR2_X1 U16213 ( .A(P3_rEIP_PTR19), .B(_03268__PTR17), .Z(_02461__PTR210) );
  XOR2_X1 U16214 ( .A(P3_rEIP_PTR20), .B(_03268__PTR18), .Z(_02461__PTR211) );
  XOR2_X1 U16215 ( .A(P3_rEIP_PTR21), .B(_03268__PTR19), .Z(_02461__PTR212) );
  XOR2_X1 U16216 ( .A(P3_rEIP_PTR22), .B(_03268__PTR20), .Z(_02461__PTR213) );
  XOR2_X1 U16217 ( .A(P3_rEIP_PTR23), .B(_03268__PTR21), .Z(_02461__PTR214) );
  XOR2_X1 U16218 ( .A(P3_rEIP_PTR24), .B(_03268__PTR22), .Z(_02461__PTR215) );
  XOR2_X1 U16219 ( .A(P3_rEIP_PTR25), .B(_03268__PTR23), .Z(_02461__PTR216) );
  XOR2_X1 U16220 ( .A(P3_rEIP_PTR26), .B(_03268__PTR24), .Z(_02461__PTR217) );
  XOR2_X1 U16221 ( .A(P3_rEIP_PTR27), .B(_03268__PTR25), .Z(_02461__PTR218) );
  XOR2_X1 U16222 ( .A(P3_rEIP_PTR28), .B(_03268__PTR26), .Z(_02461__PTR219) );
  XOR2_X1 U16223 ( .A(P3_rEIP_PTR29), .B(_03268__PTR27), .Z(_02461__PTR220) );
  XOR2_X1 U16224 ( .A(P3_rEIP_PTR30), .B(_03268__PTR28), .Z(_02461__PTR221) );
  XOR2_X1 U16225 ( .A(_03267_), .B(P3_rEIP_PTR1), .Z(_02461__PTR192) );
  AND2_X1 U16226 ( .A1(_03267_), .A2(P3_rEIP_PTR1), .ZN(_03268__PTR0) );
  XOR2_X1 U16227 ( .A(P3_rEIP_PTR3), .B(_03283__PTR0), .Z(_02461__PTR65) );
  XOR2_X1 U16228 ( .A(P3_rEIP_PTR4), .B(_03283__PTR1), .Z(_02461__PTR66) );
  XOR2_X1 U16229 ( .A(P3_rEIP_PTR5), .B(_03283__PTR2), .Z(_02461__PTR67) );
  XOR2_X1 U16230 ( .A(P3_rEIP_PTR6), .B(_03283__PTR3), .Z(_02461__PTR68) );
  XOR2_X1 U16231 ( .A(P3_rEIP_PTR7), .B(_03283__PTR4), .Z(_02461__PTR69) );
  XOR2_X1 U16232 ( .A(P3_rEIP_PTR8), .B(_03283__PTR5), .Z(_02461__PTR70) );
  XOR2_X1 U16233 ( .A(P3_rEIP_PTR9), .B(_03283__PTR6), .Z(_02461__PTR71) );
  XOR2_X1 U16234 ( .A(P3_rEIP_PTR10), .B(_03283__PTR7), .Z(_02461__PTR72) );
  XOR2_X1 U16235 ( .A(P3_rEIP_PTR11), .B(_03283__PTR8), .Z(_02461__PTR73) );
  XOR2_X1 U16236 ( .A(P3_rEIP_PTR12), .B(_03283__PTR9), .Z(_02461__PTR74) );
  XOR2_X1 U16237 ( .A(P3_rEIP_PTR13), .B(_03283__PTR10), .Z(_02461__PTR75) );
  XOR2_X1 U16238 ( .A(P3_rEIP_PTR14), .B(_03283__PTR11), .Z(_02461__PTR76) );
  XOR2_X1 U16239 ( .A(P3_rEIP_PTR15), .B(_03283__PTR12), .Z(_02461__PTR77) );
  XOR2_X1 U16240 ( .A(P3_rEIP_PTR16), .B(_03283__PTR13), .Z(_02461__PTR78) );
  XOR2_X1 U16241 ( .A(P3_rEIP_PTR17), .B(_03283__PTR14), .Z(_02461__PTR79) );
  XOR2_X1 U16242 ( .A(P3_rEIP_PTR18), .B(_03283__PTR15), .Z(_02461__PTR80) );
  XOR2_X1 U16243 ( .A(P3_rEIP_PTR19), .B(_03283__PTR16), .Z(_02461__PTR81) );
  XOR2_X1 U16244 ( .A(P3_rEIP_PTR20), .B(_03283__PTR17), .Z(_02461__PTR82) );
  XOR2_X1 U16245 ( .A(P3_rEIP_PTR21), .B(_03283__PTR18), .Z(_02461__PTR83) );
  XOR2_X1 U16246 ( .A(P3_rEIP_PTR22), .B(_03283__PTR19), .Z(_02461__PTR84) );
  XOR2_X1 U16247 ( .A(P3_rEIP_PTR23), .B(_03283__PTR20), .Z(_02461__PTR85) );
  XOR2_X1 U16248 ( .A(P3_rEIP_PTR24), .B(_03283__PTR21), .Z(_02461__PTR86) );
  XOR2_X1 U16249 ( .A(P3_rEIP_PTR25), .B(_03283__PTR22), .Z(_02461__PTR87) );
  XOR2_X1 U16250 ( .A(P3_rEIP_PTR26), .B(_03283__PTR23), .Z(_02461__PTR88) );
  XOR2_X1 U16251 ( .A(P3_rEIP_PTR27), .B(_03283__PTR24), .Z(_02461__PTR89) );
  XOR2_X1 U16252 ( .A(P3_rEIP_PTR28), .B(_03283__PTR25), .Z(_02461__PTR90) );
  XOR2_X1 U16253 ( .A(P3_rEIP_PTR29), .B(_03283__PTR26), .Z(_02461__PTR91) );
  XOR2_X1 U16254 ( .A(P3_rEIP_PTR30), .B(_03283__PTR27), .Z(_02461__PTR92) );
  XOR2_X1 U16255 ( .A(P3_rEIP_PTR31), .B(_03283__PTR28), .Z(_02461__PTR93) );
  XOR2_X1 U16256 ( .A(_03282_), .B(P3_rEIP_PTR2), .Z(_02461__PTR64) );
  AND2_X1 U16257 ( .A1(_03282_), .A2(P3_rEIP_PTR2), .ZN(_03283__PTR0) );
  AND2_X1 U16258 ( .A1(_05730__PTR3), .A2(P3_Datao_PTR2), .ZN(_05634_) );
  AND2_X1 U16259 ( .A1(_05730__PTR5), .A2(P3_Datao_PTR4), .ZN(_05635_) );
  AND2_X1 U16260 ( .A1(_05730__PTR7), .A2(P3_Datao_PTR6), .ZN(_05636_) );
  AND2_X1 U16261 ( .A1(_05730__PTR9), .A2(P3_Datao_PTR8), .ZN(_05637_) );
  AND2_X1 U16262 ( .A1(_05730__PTR11), .A2(P3_Datao_PTR10), .ZN(_05638_) );
  AND2_X1 U16263 ( .A1(_05730__PTR13), .A2(P3_Datao_PTR12), .ZN(_05639_) );
  AND2_X1 U16264 ( .A1(_05730__PTR15), .A2(P3_Datao_PTR14), .ZN(_05640_) );
  AND2_X1 U16265 ( .A1(_05730__PTR17), .A2(P3_Datao_PTR16), .ZN(_05641_) );
  AND2_X1 U16266 ( .A1(_05730__PTR19), .A2(P3_Datao_PTR18), .ZN(_05642_) );
  AND2_X1 U16267 ( .A1(_05730__PTR21), .A2(P3_Datao_PTR20), .ZN(_05643_) );
  AND2_X1 U16268 ( .A1(_05730__PTR23), .A2(P3_Datao_PTR22), .ZN(_05644_) );
  AND2_X1 U16269 ( .A1(_05730__PTR25), .A2(P3_Datao_PTR24), .ZN(_05645_) );
  AND2_X1 U16270 ( .A1(_05730__PTR27), .A2(P3_Datao_PTR26), .ZN(_05646_) );
  AND2_X1 U16271 ( .A1(_05730__PTR29), .A2(P3_Datao_PTR28), .ZN(_05647_) );
  AND2_X1 U16272 ( .A1(_05664_), .A2(_05689_), .ZN(_05649_) );
  AND2_X1 U16273 ( .A1(_05666_), .A2(_05691_), .ZN(_05650_) );
  AND2_X1 U16274 ( .A1(_05668_), .A2(_05693_), .ZN(_05651_) );
  AND2_X1 U16275 ( .A1(_05670_), .A2(_05695_), .ZN(_05652_) );
  AND2_X1 U16276 ( .A1(_05672_), .A2(_05697_), .ZN(_05653_) );
  AND2_X1 U16277 ( .A1(_05674_), .A2(_05699_), .ZN(_05654_) );
  AND2_X1 U16278 ( .A1(_05676_), .A2(_05701_), .ZN(_05655_) );
  AND2_X1 U16279 ( .A1(_05677_), .A2(_05729__PTR3), .ZN(_05656_) );
  AND2_X1 U16280 ( .A1(_05679_), .A2(_05703_), .ZN(_05657_) );
  AND2_X1 U16281 ( .A1(_05681_), .A2(_05705_), .ZN(_05658_) );
  AND2_X1 U16282 ( .A1(_05683_), .A2(_05707_), .ZN(_05659_) );
  AND2_X1 U16283 ( .A1(_05684_), .A2(_05729__PTR7), .ZN(_05660_) );
  AND2_X1 U16284 ( .A1(_05686_), .A2(_05709_), .ZN(_05661_) );
  AND2_X1 U16285 ( .A1(_05687_), .A2(_05729__PTR15), .ZN(_05662_) );
  AND2_X1 U16286 ( .A1(_05730__PTR3), .A2(_05730__PTR2), .ZN(_05648_) );
  AND2_X1 U16287 ( .A1(_05730__PTR5), .A2(_05730__PTR4), .ZN(_05663_) );
  AND2_X1 U16288 ( .A1(_05730__PTR7), .A2(_05730__PTR6), .ZN(_05664_) );
  AND2_X1 U16289 ( .A1(_05730__PTR9), .A2(_05730__PTR8), .ZN(_05665_) );
  AND2_X1 U16290 ( .A1(_05730__PTR11), .A2(_05730__PTR10), .ZN(_05666_) );
  AND2_X1 U16291 ( .A1(_05730__PTR13), .A2(_05730__PTR12), .ZN(_05667_) );
  AND2_X1 U16292 ( .A1(_05730__PTR15), .A2(_05730__PTR14), .ZN(_05668_) );
  AND2_X1 U16293 ( .A1(_05730__PTR17), .A2(_05730__PTR16), .ZN(_05669_) );
  AND2_X1 U16294 ( .A1(_05730__PTR19), .A2(_05730__PTR18), .ZN(_05670_) );
  AND2_X1 U16295 ( .A1(_05730__PTR21), .A2(_05730__PTR20), .ZN(_05671_) );
  AND2_X1 U16296 ( .A1(_05730__PTR23), .A2(_05730__PTR22), .ZN(_05672_) );
  AND2_X1 U16297 ( .A1(_05730__PTR25), .A2(_05730__PTR24), .ZN(_05673_) );
  AND2_X1 U16298 ( .A1(_05730__PTR27), .A2(_05730__PTR26), .ZN(_05674_) );
  AND2_X1 U16299 ( .A1(_05730__PTR29), .A2(_05730__PTR28), .ZN(_05675_) );
  AND2_X1 U16300 ( .A1(_05728__PTR31), .A2(P3_Datao_PTR30), .ZN(_05676_) );
  AND2_X1 U16301 ( .A1(_05664_), .A2(_05663_), .ZN(_05677_) );
  AND2_X1 U16302 ( .A1(_05666_), .A2(_05665_), .ZN(_05678_) );
  AND2_X1 U16303 ( .A1(_05668_), .A2(_05667_), .ZN(_05679_) );
  AND2_X1 U16304 ( .A1(_05670_), .A2(_05669_), .ZN(_05680_) );
  AND2_X1 U16305 ( .A1(_05672_), .A2(_05671_), .ZN(_05681_) );
  AND2_X1 U16306 ( .A1(_05674_), .A2(_05673_), .ZN(_05682_) );
  AND2_X1 U16307 ( .A1(_05676_), .A2(_05675_), .ZN(_05683_) );
  AND2_X1 U16308 ( .A1(_05679_), .A2(_05678_), .ZN(_05684_) );
  AND2_X1 U16309 ( .A1(_05681_), .A2(_05680_), .ZN(_05685_) );
  AND2_X1 U16310 ( .A1(_05683_), .A2(_05682_), .ZN(_05686_) );
  AND2_X1 U16311 ( .A1(_05686_), .A2(_05685_), .ZN(_05687_) );
  OR2_X1 U16312 ( .A1(P3_Datao_PTR3), .A2(_05634_), .ZN(_05688_) );
  OR2_X1 U16313 ( .A1(P3_Datao_PTR5), .A2(_05635_), .ZN(_05689_) );
  OR2_X1 U16314 ( .A1(P3_Datao_PTR7), .A2(_05636_), .ZN(_05690_) );
  OR2_X1 U16315 ( .A1(P3_Datao_PTR9), .A2(_05637_), .ZN(_05691_) );
  OR2_X1 U16316 ( .A1(P3_Datao_PTR11), .A2(_05638_), .ZN(_05692_) );
  OR2_X1 U16317 ( .A1(P3_Datao_PTR13), .A2(_05639_), .ZN(_05693_) );
  OR2_X1 U16318 ( .A1(P3_Datao_PTR15), .A2(_05640_), .ZN(_05694_) );
  OR2_X1 U16319 ( .A1(P3_Datao_PTR17), .A2(_05641_), .ZN(_05695_) );
  OR2_X1 U16320 ( .A1(P3_Datao_PTR19), .A2(_05642_), .ZN(_05696_) );
  OR2_X1 U16321 ( .A1(P3_Datao_PTR21), .A2(_05643_), .ZN(_05697_) );
  OR2_X1 U16322 ( .A1(P3_Datao_PTR23), .A2(_05644_), .ZN(_05698_) );
  OR2_X1 U16323 ( .A1(P3_Datao_PTR25), .A2(_05645_), .ZN(_05699_) );
  OR2_X1 U16324 ( .A1(P3_Datao_PTR27), .A2(_05646_), .ZN(_05700_) );
  OR2_X1 U16325 ( .A1(P3_Datao_PTR29), .A2(_05647_), .ZN(_05701_) );
  OR2_X1 U16326 ( .A1(_05688_), .A2(_05648_), .ZN(_05729__PTR3) );
  OR2_X1 U16327 ( .A1(_05690_), .A2(_05649_), .ZN(_05702_) );
  OR2_X1 U16328 ( .A1(_05692_), .A2(_05650_), .ZN(_05703_) );
  OR2_X1 U16329 ( .A1(_05694_), .A2(_05651_), .ZN(_05704_) );
  OR2_X1 U16330 ( .A1(_05696_), .A2(_05652_), .ZN(_05705_) );
  OR2_X1 U16331 ( .A1(_05698_), .A2(_05653_), .ZN(_05706_) );
  OR2_X1 U16332 ( .A1(_05700_), .A2(_05654_), .ZN(_05707_) );
  OR2_X1 U16333 ( .A1(_05702_), .A2(_05656_), .ZN(_05729__PTR7) );
  OR2_X1 U16334 ( .A1(_05704_), .A2(_05657_), .ZN(_05708_) );
  OR2_X1 U16335 ( .A1(_05706_), .A2(_05658_), .ZN(_05709_) );
  OR2_X1 U16336 ( .A1(_05655_), .A2(_05659_), .ZN(_05710_) );
  OR2_X1 U16337 ( .A1(_05708_), .A2(_05660_), .ZN(_05729__PTR15) );
  OR2_X1 U16338 ( .A1(_05710_), .A2(_05661_), .ZN(_05711_) );
  OR2_X1 U16339 ( .A1(_05711_), .A2(_05662_), .ZN(_05729__PTR31) );
  AND2_X1 U16340 ( .A1(_05726__PTR3), .A2(P2_Datao_PTR2), .ZN(_05556_) );
  AND2_X1 U16341 ( .A1(_05726__PTR5), .A2(P2_Datao_PTR4), .ZN(_05557_) );
  AND2_X1 U16342 ( .A1(_05726__PTR7), .A2(P2_Datao_PTR6), .ZN(_05558_) );
  AND2_X1 U16343 ( .A1(_05726__PTR9), .A2(P2_Datao_PTR8), .ZN(_05559_) );
  AND2_X1 U16344 ( .A1(_05726__PTR11), .A2(P2_Datao_PTR10), .ZN(_05560_) );
  AND2_X1 U16345 ( .A1(_05726__PTR13), .A2(P2_Datao_PTR12), .ZN(_05561_) );
  AND2_X1 U16346 ( .A1(_05726__PTR15), .A2(P2_Datao_PTR14), .ZN(_05562_) );
  AND2_X1 U16347 ( .A1(_05726__PTR17), .A2(P2_Datao_PTR16), .ZN(_05563_) );
  AND2_X1 U16348 ( .A1(_05726__PTR19), .A2(P2_Datao_PTR18), .ZN(_05564_) );
  AND2_X1 U16349 ( .A1(_05726__PTR21), .A2(P2_Datao_PTR20), .ZN(_05565_) );
  AND2_X1 U16350 ( .A1(_05726__PTR23), .A2(P2_Datao_PTR22), .ZN(_05566_) );
  AND2_X1 U16351 ( .A1(_05726__PTR25), .A2(P2_Datao_PTR24), .ZN(_05567_) );
  AND2_X1 U16352 ( .A1(_05726__PTR27), .A2(P2_Datao_PTR26), .ZN(_05568_) );
  AND2_X1 U16353 ( .A1(_05726__PTR29), .A2(P2_Datao_PTR28), .ZN(_05569_) );
  AND2_X1 U16354 ( .A1(_05586_), .A2(_05611_), .ZN(_05571_) );
  AND2_X1 U16355 ( .A1(_05588_), .A2(_05613_), .ZN(_05572_) );
  AND2_X1 U16356 ( .A1(_05590_), .A2(_05615_), .ZN(_05573_) );
  AND2_X1 U16357 ( .A1(_05592_), .A2(_05617_), .ZN(_05574_) );
  AND2_X1 U16358 ( .A1(_05594_), .A2(_05619_), .ZN(_05575_) );
  AND2_X1 U16359 ( .A1(_05596_), .A2(_05621_), .ZN(_05576_) );
  AND2_X1 U16360 ( .A1(_05598_), .A2(_05623_), .ZN(_05577_) );
  AND2_X1 U16361 ( .A1(_05599_), .A2(_05725__PTR3), .ZN(_05578_) );
  AND2_X1 U16362 ( .A1(_05601_), .A2(_05625_), .ZN(_05579_) );
  AND2_X1 U16363 ( .A1(_05603_), .A2(_05627_), .ZN(_05580_) );
  AND2_X1 U16364 ( .A1(_05605_), .A2(_05629_), .ZN(_05581_) );
  AND2_X1 U16365 ( .A1(_05606_), .A2(_05725__PTR7), .ZN(_05582_) );
  AND2_X1 U16366 ( .A1(_05608_), .A2(_05631_), .ZN(_05583_) );
  AND2_X1 U16367 ( .A1(_05609_), .A2(_05725__PTR15), .ZN(_05584_) );
  AND2_X1 U16368 ( .A1(_05726__PTR3), .A2(_05726__PTR2), .ZN(_05570_) );
  AND2_X1 U16369 ( .A1(_05726__PTR5), .A2(_05726__PTR4), .ZN(_05585_) );
  AND2_X1 U16370 ( .A1(_05726__PTR7), .A2(_05726__PTR6), .ZN(_05586_) );
  AND2_X1 U16371 ( .A1(_05726__PTR9), .A2(_05726__PTR8), .ZN(_05587_) );
  AND2_X1 U16372 ( .A1(_05726__PTR11), .A2(_05726__PTR10), .ZN(_05588_) );
  AND2_X1 U16373 ( .A1(_05726__PTR13), .A2(_05726__PTR12), .ZN(_05589_) );
  AND2_X1 U16374 ( .A1(_05726__PTR15), .A2(_05726__PTR14), .ZN(_05590_) );
  AND2_X1 U16375 ( .A1(_05726__PTR17), .A2(_05726__PTR16), .ZN(_05591_) );
  AND2_X1 U16376 ( .A1(_05726__PTR19), .A2(_05726__PTR18), .ZN(_05592_) );
  AND2_X1 U16377 ( .A1(_05726__PTR21), .A2(_05726__PTR20), .ZN(_05593_) );
  AND2_X1 U16378 ( .A1(_05726__PTR23), .A2(_05726__PTR22), .ZN(_05594_) );
  AND2_X1 U16379 ( .A1(_05726__PTR25), .A2(_05726__PTR24), .ZN(_05595_) );
  AND2_X1 U16380 ( .A1(_05726__PTR27), .A2(_05726__PTR26), .ZN(_05596_) );
  AND2_X1 U16381 ( .A1(_05726__PTR29), .A2(_05726__PTR28), .ZN(_05597_) );
  AND2_X1 U16382 ( .A1(_05724__PTR31), .A2(P2_Datao_PTR30), .ZN(_05598_) );
  AND2_X1 U16383 ( .A1(_05586_), .A2(_05585_), .ZN(_05599_) );
  AND2_X1 U16384 ( .A1(_05588_), .A2(_05587_), .ZN(_05600_) );
  AND2_X1 U16385 ( .A1(_05590_), .A2(_05589_), .ZN(_05601_) );
  AND2_X1 U16386 ( .A1(_05592_), .A2(_05591_), .ZN(_05602_) );
  AND2_X1 U16387 ( .A1(_05594_), .A2(_05593_), .ZN(_05603_) );
  AND2_X1 U16388 ( .A1(_05596_), .A2(_05595_), .ZN(_05604_) );
  AND2_X1 U16389 ( .A1(_05598_), .A2(_05597_), .ZN(_05605_) );
  AND2_X1 U16390 ( .A1(_05601_), .A2(_05600_), .ZN(_05606_) );
  AND2_X1 U16391 ( .A1(_05603_), .A2(_05602_), .ZN(_05607_) );
  AND2_X1 U16392 ( .A1(_05605_), .A2(_05604_), .ZN(_05608_) );
  AND2_X1 U16393 ( .A1(_05608_), .A2(_05607_), .ZN(_05609_) );
  OR2_X1 U16394 ( .A1(P2_Datao_PTR3), .A2(_05556_), .ZN(_05610_) );
  OR2_X1 U16395 ( .A1(P2_Datao_PTR5), .A2(_05557_), .ZN(_05611_) );
  OR2_X1 U16396 ( .A1(P2_Datao_PTR7), .A2(_05558_), .ZN(_05612_) );
  OR2_X1 U16397 ( .A1(P2_Datao_PTR9), .A2(_05559_), .ZN(_05613_) );
  OR2_X1 U16398 ( .A1(P2_Datao_PTR11), .A2(_05560_), .ZN(_05614_) );
  OR2_X1 U16399 ( .A1(P2_Datao_PTR13), .A2(_05561_), .ZN(_05615_) );
  OR2_X1 U16400 ( .A1(P2_Datao_PTR15), .A2(_05562_), .ZN(_05616_) );
  OR2_X1 U16401 ( .A1(P2_Datao_PTR17), .A2(_05563_), .ZN(_05617_) );
  OR2_X1 U16402 ( .A1(P2_Datao_PTR19), .A2(_05564_), .ZN(_05618_) );
  OR2_X1 U16403 ( .A1(P2_Datao_PTR21), .A2(_05565_), .ZN(_05619_) );
  OR2_X1 U16404 ( .A1(P2_Datao_PTR23), .A2(_05566_), .ZN(_05620_) );
  OR2_X1 U16405 ( .A1(P2_Datao_PTR25), .A2(_05567_), .ZN(_05621_) );
  OR2_X1 U16406 ( .A1(P2_Datao_PTR27), .A2(_05568_), .ZN(_05622_) );
  OR2_X1 U16407 ( .A1(P2_Datao_PTR29), .A2(_05569_), .ZN(_05623_) );
  OR2_X1 U16408 ( .A1(_05610_), .A2(_05570_), .ZN(_05725__PTR3) );
  OR2_X1 U16409 ( .A1(_05612_), .A2(_05571_), .ZN(_05624_) );
  OR2_X1 U16410 ( .A1(_05614_), .A2(_05572_), .ZN(_05625_) );
  OR2_X1 U16411 ( .A1(_05616_), .A2(_05573_), .ZN(_05626_) );
  OR2_X1 U16412 ( .A1(_05618_), .A2(_05574_), .ZN(_05627_) );
  OR2_X1 U16413 ( .A1(_05620_), .A2(_05575_), .ZN(_05628_) );
  OR2_X1 U16414 ( .A1(_05622_), .A2(_05576_), .ZN(_05629_) );
  OR2_X1 U16415 ( .A1(_05624_), .A2(_05578_), .ZN(_05725__PTR7) );
  OR2_X1 U16416 ( .A1(_05626_), .A2(_05579_), .ZN(_05630_) );
  OR2_X1 U16417 ( .A1(_05628_), .A2(_05580_), .ZN(_05631_) );
  OR2_X1 U16418 ( .A1(_05577_), .A2(_05581_), .ZN(_05632_) );
  OR2_X1 U16419 ( .A1(_05630_), .A2(_05582_), .ZN(_05725__PTR15) );
  OR2_X1 U16420 ( .A1(_05632_), .A2(_05583_), .ZN(_05633_) );
  OR2_X1 U16421 ( .A1(_05633_), .A2(_05584_), .ZN(_05725__PTR31) );
  AND2_X1 U16422 ( .A1(_05722__PTR3), .A2(P1_Datao_PTR2), .ZN(_05478_) );
  AND2_X1 U16423 ( .A1(_05722__PTR5), .A2(P1_Datao_PTR4), .ZN(_05479_) );
  AND2_X1 U16424 ( .A1(_05722__PTR7), .A2(P1_Datao_PTR6), .ZN(_05480_) );
  AND2_X1 U16425 ( .A1(_05722__PTR9), .A2(P1_Datao_PTR8), .ZN(_05481_) );
  AND2_X1 U16426 ( .A1(_05722__PTR11), .A2(P1_Datao_PTR10), .ZN(_05482_) );
  AND2_X1 U16427 ( .A1(_05722__PTR13), .A2(P1_Datao_PTR12), .ZN(_05483_) );
  AND2_X1 U16428 ( .A1(_05722__PTR15), .A2(P1_Datao_PTR14), .ZN(_05484_) );
  AND2_X1 U16429 ( .A1(_05722__PTR17), .A2(P1_Datao_PTR16), .ZN(_05485_) );
  AND2_X1 U16430 ( .A1(_05722__PTR19), .A2(P1_Datao_PTR18), .ZN(_05486_) );
  AND2_X1 U16431 ( .A1(_05722__PTR21), .A2(P1_Datao_PTR20), .ZN(_05487_) );
  AND2_X1 U16432 ( .A1(_05722__PTR23), .A2(P1_Datao_PTR22), .ZN(_05488_) );
  AND2_X1 U16433 ( .A1(_05722__PTR25), .A2(P1_Datao_PTR24), .ZN(_05489_) );
  AND2_X1 U16434 ( .A1(_05722__PTR27), .A2(P1_Datao_PTR26), .ZN(_05490_) );
  AND2_X1 U16435 ( .A1(_05722__PTR29), .A2(P1_Datao_PTR28), .ZN(_05491_) );
  AND2_X1 U16436 ( .A1(_05508_), .A2(_05533_), .ZN(_05493_) );
  AND2_X1 U16437 ( .A1(_05510_), .A2(_05535_), .ZN(_05494_) );
  AND2_X1 U16438 ( .A1(_05512_), .A2(_05537_), .ZN(_05495_) );
  AND2_X1 U16439 ( .A1(_05514_), .A2(_05539_), .ZN(_05496_) );
  AND2_X1 U16440 ( .A1(_05516_), .A2(_05541_), .ZN(_05497_) );
  AND2_X1 U16441 ( .A1(_05518_), .A2(_05543_), .ZN(_05498_) );
  AND2_X1 U16442 ( .A1(_05520_), .A2(_05545_), .ZN(_05499_) );
  AND2_X1 U16443 ( .A1(_05521_), .A2(_05721__PTR3), .ZN(_05500_) );
  AND2_X1 U16444 ( .A1(_05523_), .A2(_05547_), .ZN(_05501_) );
  AND2_X1 U16445 ( .A1(_05525_), .A2(_05549_), .ZN(_05502_) );
  AND2_X1 U16446 ( .A1(_05527_), .A2(_05551_), .ZN(_05503_) );
  AND2_X1 U16447 ( .A1(_05528_), .A2(_05721__PTR7), .ZN(_05504_) );
  AND2_X1 U16448 ( .A1(_05530_), .A2(_05553_), .ZN(_05505_) );
  AND2_X1 U16449 ( .A1(_05531_), .A2(_05721__PTR15), .ZN(_05506_) );
  AND2_X1 U16450 ( .A1(_05722__PTR3), .A2(_05722__PTR2), .ZN(_05492_) );
  AND2_X1 U16451 ( .A1(_05722__PTR5), .A2(_05722__PTR4), .ZN(_05507_) );
  AND2_X1 U16452 ( .A1(_05722__PTR7), .A2(_05722__PTR6), .ZN(_05508_) );
  AND2_X1 U16453 ( .A1(_05722__PTR9), .A2(_05722__PTR8), .ZN(_05509_) );
  AND2_X1 U16454 ( .A1(_05722__PTR11), .A2(_05722__PTR10), .ZN(_05510_) );
  AND2_X1 U16455 ( .A1(_05722__PTR13), .A2(_05722__PTR12), .ZN(_05511_) );
  AND2_X1 U16456 ( .A1(_05722__PTR15), .A2(_05722__PTR14), .ZN(_05512_) );
  AND2_X1 U16457 ( .A1(_05722__PTR17), .A2(_05722__PTR16), .ZN(_05513_) );
  AND2_X1 U16458 ( .A1(_05722__PTR19), .A2(_05722__PTR18), .ZN(_05514_) );
  AND2_X1 U16459 ( .A1(_05722__PTR21), .A2(_05722__PTR20), .ZN(_05515_) );
  AND2_X1 U16460 ( .A1(_05722__PTR23), .A2(_05722__PTR22), .ZN(_05516_) );
  AND2_X1 U16461 ( .A1(_05722__PTR25), .A2(_05722__PTR24), .ZN(_05517_) );
  AND2_X1 U16462 ( .A1(_05722__PTR27), .A2(_05722__PTR26), .ZN(_05518_) );
  AND2_X1 U16463 ( .A1(_05722__PTR29), .A2(_05722__PTR28), .ZN(_05519_) );
  AND2_X1 U16464 ( .A1(_05720__PTR31), .A2(P1_Datao_PTR30), .ZN(_05520_) );
  AND2_X1 U16465 ( .A1(_05508_), .A2(_05507_), .ZN(_05521_) );
  AND2_X1 U16466 ( .A1(_05510_), .A2(_05509_), .ZN(_05522_) );
  AND2_X1 U16467 ( .A1(_05512_), .A2(_05511_), .ZN(_05523_) );
  AND2_X1 U16468 ( .A1(_05514_), .A2(_05513_), .ZN(_05524_) );
  AND2_X1 U16469 ( .A1(_05516_), .A2(_05515_), .ZN(_05525_) );
  AND2_X1 U16470 ( .A1(_05518_), .A2(_05517_), .ZN(_05526_) );
  AND2_X1 U16471 ( .A1(_05520_), .A2(_05519_), .ZN(_05527_) );
  AND2_X1 U16472 ( .A1(_05523_), .A2(_05522_), .ZN(_05528_) );
  AND2_X1 U16473 ( .A1(_05525_), .A2(_05524_), .ZN(_05529_) );
  AND2_X1 U16474 ( .A1(_05527_), .A2(_05526_), .ZN(_05530_) );
  AND2_X1 U16475 ( .A1(_05530_), .A2(_05529_), .ZN(_05531_) );
  OR2_X1 U16476 ( .A1(P1_Datao_PTR3), .A2(_05478_), .ZN(_05532_) );
  OR2_X1 U16477 ( .A1(P1_Datao_PTR5), .A2(_05479_), .ZN(_05533_) );
  OR2_X1 U16478 ( .A1(P1_Datao_PTR7), .A2(_05480_), .ZN(_05534_) );
  OR2_X1 U16479 ( .A1(P1_Datao_PTR9), .A2(_05481_), .ZN(_05535_) );
  OR2_X1 U16480 ( .A1(P1_Datao_PTR11), .A2(_05482_), .ZN(_05536_) );
  OR2_X1 U16481 ( .A1(P1_Datao_PTR13), .A2(_05483_), .ZN(_05537_) );
  OR2_X1 U16482 ( .A1(P1_Datao_PTR15), .A2(_05484_), .ZN(_05538_) );
  OR2_X1 U16483 ( .A1(P1_Datao_PTR17), .A2(_05485_), .ZN(_05539_) );
  OR2_X1 U16484 ( .A1(P1_Datao_PTR19), .A2(_05486_), .ZN(_05540_) );
  OR2_X1 U16485 ( .A1(P1_Datao_PTR21), .A2(_05487_), .ZN(_05541_) );
  OR2_X1 U16486 ( .A1(P1_Datao_PTR23), .A2(_05488_), .ZN(_05542_) );
  OR2_X1 U16487 ( .A1(P1_Datao_PTR25), .A2(_05489_), .ZN(_05543_) );
  OR2_X1 U16488 ( .A1(P1_Datao_PTR27), .A2(_05490_), .ZN(_05544_) );
  OR2_X1 U16489 ( .A1(P1_Datao_PTR29), .A2(_05491_), .ZN(_05545_) );
  OR2_X1 U16490 ( .A1(_05532_), .A2(_05492_), .ZN(_05721__PTR3) );
  OR2_X1 U16491 ( .A1(_05534_), .A2(_05493_), .ZN(_05546_) );
  OR2_X1 U16492 ( .A1(_05536_), .A2(_05494_), .ZN(_05547_) );
  OR2_X1 U16493 ( .A1(_05538_), .A2(_05495_), .ZN(_05548_) );
  OR2_X1 U16494 ( .A1(_05540_), .A2(_05496_), .ZN(_05549_) );
  OR2_X1 U16495 ( .A1(_05542_), .A2(_05497_), .ZN(_05550_) );
  OR2_X1 U16496 ( .A1(_05544_), .A2(_05498_), .ZN(_05551_) );
  OR2_X1 U16497 ( .A1(_05546_), .A2(_05500_), .ZN(_05721__PTR7) );
  OR2_X1 U16498 ( .A1(_05548_), .A2(_05501_), .ZN(_05552_) );
  OR2_X1 U16499 ( .A1(_05550_), .A2(_05502_), .ZN(_05553_) );
  OR2_X1 U16500 ( .A1(_05499_), .A2(_05503_), .ZN(_05554_) );
  OR2_X1 U16501 ( .A1(_05552_), .A2(_05504_), .ZN(_05721__PTR15) );
  OR2_X1 U16502 ( .A1(_05554_), .A2(_05505_), .ZN(_05555_) );
  OR2_X1 U16503 ( .A1(_05555_), .A2(_05506_), .ZN(_05721__PTR31) );
  AND2_X1 U16504 ( .A1(_05712__PTR3), .A2(P2_Address_PTR2), .ZN(_05407_) );
  AND2_X1 U16505 ( .A1(_05712__PTR5), .A2(P2_Address_PTR4), .ZN(_05408_) );
  AND2_X1 U16506 ( .A1(_05712__PTR7), .A2(P2_Address_PTR6), .ZN(_05409_) );
  AND2_X1 U16507 ( .A1(_05712__PTR9), .A2(P2_Address_PTR8), .ZN(_05410_) );
  AND2_X1 U16508 ( .A1(_05712__PTR11), .A2(P2_Address_PTR10), .ZN(_05411_) );
  AND2_X1 U16509 ( .A1(_05712__PTR13), .A2(P2_Address_PTR12), .ZN(_05412_) );
  AND2_X1 U16510 ( .A1(_05712__PTR15), .A2(P2_Address_PTR14), .ZN(_05413_) );
  AND2_X1 U16511 ( .A1(_05712__PTR17), .A2(P2_Address_PTR16), .ZN(_05414_) );
  AND2_X1 U16512 ( .A1(_05712__PTR19), .A2(P2_Address_PTR18), .ZN(_05415_) );
  AND2_X1 U16513 ( .A1(_05712__PTR21), .A2(P2_Address_PTR20), .ZN(_05416_) );
  AND2_X1 U16514 ( .A1(_05712__PTR23), .A2(P2_Address_PTR22), .ZN(_05417_) );
  AND2_X1 U16515 ( .A1(_05712__PTR25), .A2(P2_Address_PTR24), .ZN(_05418_) );
  AND2_X1 U16516 ( .A1(_05712__PTR27), .A2(P2_Address_PTR26), .ZN(_05419_) );
  AND2_X1 U16517 ( .A1(P2_Address_PTR29), .A2(P2_Address_PTR28), .ZN(_05420_) );
  AND2_X1 U16518 ( .A1(_05386_), .A2(_05435_), .ZN(_05421_) );
  AND2_X1 U16519 ( .A1(_05388_), .A2(_05437_), .ZN(_05422_) );
  AND2_X1 U16520 ( .A1(_05390_), .A2(_05439_), .ZN(_05423_) );
  AND2_X1 U16521 ( .A1(_05392_), .A2(_05441_), .ZN(_05424_) );
  AND2_X1 U16522 ( .A1(_05394_), .A2(_05443_), .ZN(_05425_) );
  AND2_X1 U16523 ( .A1(_05396_), .A2(_05445_), .ZN(_05426_) );
  AND2_X1 U16524 ( .A1(_05398_), .A2(_05715__PTR3), .ZN(_05427_) );
  AND2_X1 U16525 ( .A1(_05400_), .A2(_05448_), .ZN(_05428_) );
  AND2_X1 U16526 ( .A1(_05402_), .A2(_05450_), .ZN(_05429_) );
  AND2_X1 U16527 ( .A1(_05404_), .A2(_05715__PTR7), .ZN(_05430_) );
  AND2_X1 U16528 ( .A1(_05405_), .A2(_05715__PTR15), .ZN(_05431_) );
  AND2_X1 U16529 ( .A1(_05403_), .A2(_05715__PTR23), .ZN(_05432_) );
  AND2_X1 U16530 ( .A1(_05397_), .A2(_05715__PTR27), .ZN(_05433_) );
  OR2_X1 U16531 ( .A1(P2_Address_PTR3), .A2(_05407_), .ZN(_05434_) );
  OR2_X1 U16532 ( .A1(P2_Address_PTR5), .A2(_05408_), .ZN(_05435_) );
  OR2_X1 U16533 ( .A1(P2_Address_PTR7), .A2(_05409_), .ZN(_05436_) );
  OR2_X1 U16534 ( .A1(P2_Address_PTR9), .A2(_05410_), .ZN(_05437_) );
  OR2_X1 U16535 ( .A1(P2_Address_PTR11), .A2(_05411_), .ZN(_05438_) );
  OR2_X1 U16536 ( .A1(P2_Address_PTR13), .A2(_05412_), .ZN(_05439_) );
  OR2_X1 U16537 ( .A1(P2_Address_PTR15), .A2(_05413_), .ZN(_05440_) );
  OR2_X1 U16538 ( .A1(P2_Address_PTR17), .A2(_05414_), .ZN(_05441_) );
  OR2_X1 U16539 ( .A1(P2_Address_PTR19), .A2(_05415_), .ZN(_05442_) );
  OR2_X1 U16540 ( .A1(P2_Address_PTR21), .A2(_05416_), .ZN(_05443_) );
  OR2_X1 U16541 ( .A1(P2_Address_PTR23), .A2(_05417_), .ZN(_05444_) );
  OR2_X1 U16542 ( .A1(P2_Address_PTR25), .A2(_05418_), .ZN(_05445_) );
  OR2_X1 U16543 ( .A1(P2_Address_PTR27), .A2(_05419_), .ZN(_05446_) );
  OR2_X1 U16544 ( .A1(_05434_), .A2(_05384_), .ZN(_05715__PTR3) );
  OR2_X1 U16545 ( .A1(_05436_), .A2(_05421_), .ZN(_05447_) );
  OR2_X1 U16546 ( .A1(_05438_), .A2(_05422_), .ZN(_05448_) );
  OR2_X1 U16547 ( .A1(_05440_), .A2(_05423_), .ZN(_05449_) );
  OR2_X1 U16548 ( .A1(_05442_), .A2(_05424_), .ZN(_05450_) );
  OR2_X1 U16549 ( .A1(_05444_), .A2(_05425_), .ZN(_05451_) );
  OR2_X1 U16550 ( .A1(_05446_), .A2(_05426_), .ZN(_05452_) );
  OR2_X1 U16551 ( .A1(_05447_), .A2(_05427_), .ZN(_05715__PTR7) );
  OR2_X1 U16552 ( .A1(_05449_), .A2(_05428_), .ZN(_05453_) );
  OR2_X1 U16553 ( .A1(_05451_), .A2(_05429_), .ZN(_05454_) );
  OR2_X1 U16554 ( .A1(_05453_), .A2(_05430_), .ZN(_05715__PTR15) );
  OR2_X1 U16555 ( .A1(_05454_), .A2(_05431_), .ZN(_05715__PTR23) );
  OR2_X1 U16556 ( .A1(_05452_), .A2(_05432_), .ZN(_05715__PTR27) );
  OR2_X1 U16557 ( .A1(_05420_), .A2(_05433_), .ZN(_05715__PTR29) );
  AND2_X1 U16558 ( .A1(_05712__PTR1), .A2(_05712__PTR0), .ZN(_05713__PTR1) );
  AND2_X1 U16559 ( .A1(_05384_), .A2(_05713__PTR1), .ZN(_05713__PTR3) );
  AND2_X1 U16560 ( .A1(_05398_), .A2(_05713__PTR3), .ZN(_05713__PTR7) );
  AND2_X1 U16561 ( .A1(_05404_), .A2(_05713__PTR7), .ZN(_05713__PTR15) );
  AND2_X1 U16562 ( .A1(_05712__PTR3), .A2(_05712__PTR2), .ZN(_05384_) );
  AND2_X1 U16563 ( .A1(_05712__PTR5), .A2(_05712__PTR4), .ZN(_05385_) );
  AND2_X1 U16564 ( .A1(_05712__PTR7), .A2(_05712__PTR6), .ZN(_05386_) );
  AND2_X1 U16565 ( .A1(_05712__PTR9), .A2(_05712__PTR8), .ZN(_05387_) );
  AND2_X1 U16566 ( .A1(_05712__PTR11), .A2(_05712__PTR10), .ZN(_05388_) );
  AND2_X1 U16567 ( .A1(_05712__PTR13), .A2(_05712__PTR12), .ZN(_05389_) );
  AND2_X1 U16568 ( .A1(_05712__PTR15), .A2(_05712__PTR14), .ZN(_05390_) );
  AND2_X1 U16569 ( .A1(_05712__PTR17), .A2(_05712__PTR16), .ZN(_05391_) );
  AND2_X1 U16570 ( .A1(_05712__PTR19), .A2(_05712__PTR18), .ZN(_05392_) );
  AND2_X1 U16571 ( .A1(_05712__PTR21), .A2(_05712__PTR20), .ZN(_05393_) );
  AND2_X1 U16572 ( .A1(_05712__PTR23), .A2(_05712__PTR22), .ZN(_05394_) );
  AND2_X1 U16573 ( .A1(_05712__PTR25), .A2(_05712__PTR24), .ZN(_05395_) );
  AND2_X1 U16574 ( .A1(_05712__PTR27), .A2(_05712__PTR26), .ZN(_05396_) );
  AND2_X1 U16575 ( .A1(P2_Address_PTR29), .A2(_05712__PTR28), .ZN(_05397_) );
  AND2_X1 U16576 ( .A1(_05386_), .A2(_05385_), .ZN(_05398_) );
  AND2_X1 U16577 ( .A1(_05388_), .A2(_05387_), .ZN(_05399_) );
  AND2_X1 U16578 ( .A1(_05390_), .A2(_05389_), .ZN(_05400_) );
  AND2_X1 U16579 ( .A1(_05392_), .A2(_05391_), .ZN(_05401_) );
  AND2_X1 U16580 ( .A1(_05394_), .A2(_05393_), .ZN(_05402_) );
  AND2_X1 U16581 ( .A1(_05396_), .A2(_05395_), .ZN(_05403_) );
  AND2_X1 U16582 ( .A1(_05400_), .A2(_05399_), .ZN(_05404_) );
  AND2_X1 U16583 ( .A1(_05402_), .A2(_05401_), .ZN(_05405_) );
  AND2_X1 U16584 ( .A1(_05405_), .A2(_05713__PTR15), .ZN(_05713__PTR23) );
  AND2_X1 U16585 ( .A1(_05403_), .A2(_05713__PTR23), .ZN(_05713__PTR27) );
  AND2_X1 U16586 ( .A1(_05397_), .A2(_05713__PTR27), .ZN(_05406_) );
  OR2_X1 U16587 ( .A1(_05712__PTR29), .A2(_05406_), .ZN(_05713__PTR29) );
  AND2_X1 U16588 ( .A1(_05717__PTR1), .A2(_05717__PTR0), .ZN(_05718__PTR1) );
  AND2_X1 U16589 ( .A1(_05455_), .A2(_05718__PTR1), .ZN(_05718__PTR3) );
  AND2_X1 U16590 ( .A1(_05469_), .A2(_05718__PTR3), .ZN(_05718__PTR7) );
  AND2_X1 U16591 ( .A1(_05475_), .A2(_05718__PTR7), .ZN(_05718__PTR15) );
  AND2_X1 U16592 ( .A1(_05717__PTR3), .A2(_05717__PTR2), .ZN(_05455_) );
  AND2_X1 U16593 ( .A1(_05717__PTR5), .A2(_05717__PTR4), .ZN(_05456_) );
  AND2_X1 U16594 ( .A1(_05717__PTR7), .A2(_05717__PTR6), .ZN(_05457_) );
  AND2_X1 U16595 ( .A1(_05717__PTR9), .A2(_05717__PTR8), .ZN(_05458_) );
  AND2_X1 U16596 ( .A1(_05717__PTR11), .A2(_05717__PTR10), .ZN(_05459_) );
  AND2_X1 U16597 ( .A1(_05717__PTR13), .A2(_05717__PTR12), .ZN(_05460_) );
  AND2_X1 U16598 ( .A1(_05717__PTR15), .A2(_05717__PTR14), .ZN(_05461_) );
  AND2_X1 U16599 ( .A1(_05717__PTR17), .A2(_05717__PTR16), .ZN(_05462_) );
  AND2_X1 U16600 ( .A1(_05717__PTR19), .A2(_05717__PTR18), .ZN(_05463_) );
  AND2_X1 U16601 ( .A1(_05717__PTR21), .A2(_05717__PTR20), .ZN(_05464_) );
  AND2_X1 U16602 ( .A1(_05717__PTR23), .A2(_05717__PTR22), .ZN(_05465_) );
  AND2_X1 U16603 ( .A1(_05717__PTR25), .A2(_05717__PTR24), .ZN(_05466_) );
  AND2_X1 U16604 ( .A1(_05717__PTR27), .A2(_05717__PTR26), .ZN(_05467_) );
  AND2_X1 U16605 ( .A1(P1_Address_PTR29), .A2(_05717__PTR28), .ZN(_05468_) );
  AND2_X1 U16606 ( .A1(_05457_), .A2(_05456_), .ZN(_05469_) );
  AND2_X1 U16607 ( .A1(_05459_), .A2(_05458_), .ZN(_05470_) );
  AND2_X1 U16608 ( .A1(_05461_), .A2(_05460_), .ZN(_05471_) );
  AND2_X1 U16609 ( .A1(_05463_), .A2(_05462_), .ZN(_05472_) );
  AND2_X1 U16610 ( .A1(_05465_), .A2(_05464_), .ZN(_05473_) );
  AND2_X1 U16611 ( .A1(_05467_), .A2(_05466_), .ZN(_05474_) );
  AND2_X1 U16612 ( .A1(_05471_), .A2(_05470_), .ZN(_05475_) );
  AND2_X1 U16613 ( .A1(_05473_), .A2(_05472_), .ZN(_05476_) );
  AND2_X1 U16614 ( .A1(_05476_), .A2(_05718__PTR15), .ZN(_05718__PTR23) );
  AND2_X1 U16615 ( .A1(_05474_), .A2(_05718__PTR23), .ZN(_05718__PTR27) );
  AND2_X1 U16616 ( .A1(_05468_), .A2(_05718__PTR27), .ZN(_05477_) );
  OR2_X1 U16617 ( .A1(_05717__PTR29), .A2(_05477_), .ZN(_05718__PTR29) );
  AND2_X1 U16618 ( .A1(_02812__PTR1), .A2(_02750__PTR1), .ZN(_02750__PTR3) );
  AND2_X1 U16619 ( .A1(P1_P1_InstQueueRd_Addr_PTR2), .A2(_02750__PTR1), .ZN(_02750__PTR2) );
  AND2_X1 U16620 ( .A1(_02751__PTR4), .A2(_02750__PTR3), .ZN(_02753_) );
  OR2_X1 U16621 ( .A1(P1_P1_InstQueueRd_Addr_PTR4), .A2(_02753_), .ZN(_02750__PTR4) );
  AND2_X1 U16622 ( .A1(_02943__PTR4), .A2(_02944__PTR3), .ZN(_02747__PTR5) );
  OR2_X1 U16623 ( .A1(_03715_), .A2(_03712_), .ZN(_02944__PTR3) );
  AND2_X1 U16624 ( .A1(_02746__PTR1), .A2(_02746__PTR0), .ZN(_02748__PTR1) );
  AND2_X1 U16625 ( .A1(_01932__PTR59), .A2(_02746__PTR2), .ZN(_03709_) );
  AND2_X1 U16626 ( .A1(_02747__PTR5), .A2(_02746__PTR4), .ZN(_03710_) );
  AND2_X1 U16627 ( .A1(_03712_), .A2(_02748__PTR1), .ZN(_03711_) );
  AND2_X1 U16628 ( .A1(_01932__PTR59), .A2(_01932__PTR58), .ZN(_03712_) );
  AND2_X1 U16629 ( .A1(_02747__PTR5), .A2(_02749__PTR4), .ZN(_03713_) );
  AND2_X1 U16630 ( .A1(_03713_), .A2(_02748__PTR3), .ZN(_03714_) );
  OR2_X1 U16631 ( .A1(_02746__PTR3), .A2(_03709_), .ZN(_03715_) );
  OR2_X1 U16632 ( .A1(_03715_), .A2(_03711_), .ZN(_02748__PTR3) );
  OR2_X1 U16633 ( .A1(_03710_), .A2(_03714_), .ZN(_01894__PTR28) );
  AND2_X1 U16634 ( .A1(_02829__PTR1), .A2(P1_P1_InstAddrPointer_PTR0), .ZN(_02830__PTR1) );
  AND2_X1 U16635 ( .A1(_02745__PTR3), .A2(P1_P1_InstAddrPointer_PTR2), .ZN(_03629_) );
  AND2_X1 U16636 ( .A1(_02745__PTR5), .A2(P1_P1_InstAddrPointer_PTR4), .ZN(_03630_) );
  AND2_X1 U16637 ( .A1(_02745__PTR7), .A2(P1_P1_InstAddrPointer_PTR6), .ZN(_03631_) );
  AND2_X1 U16638 ( .A1(_02745__PTR9), .A2(P1_P1_InstAddrPointer_PTR8), .ZN(_03632_) );
  AND2_X1 U16639 ( .A1(_02745__PTR11), .A2(P1_P1_InstAddrPointer_PTR10), .ZN(_03633_) );
  AND2_X1 U16640 ( .A1(_02745__PTR13), .A2(P1_P1_InstAddrPointer_PTR12), .ZN(_03634_) );
  AND2_X1 U16641 ( .A1(_02745__PTR15), .A2(P1_P1_InstAddrPointer_PTR14), .ZN(_03635_) );
  AND2_X1 U16642 ( .A1(_02745__PTR17), .A2(P1_P1_InstAddrPointer_PTR16), .ZN(_03636_) );
  AND2_X1 U16643 ( .A1(_02745__PTR19), .A2(P1_P1_InstAddrPointer_PTR18), .ZN(_03637_) );
  AND2_X1 U16644 ( .A1(_02745__PTR21), .A2(P1_P1_InstAddrPointer_PTR20), .ZN(_03638_) );
  AND2_X1 U16645 ( .A1(_02745__PTR23), .A2(P1_P1_InstAddrPointer_PTR22), .ZN(_03639_) );
  AND2_X1 U16646 ( .A1(_02745__PTR25), .A2(P1_P1_InstAddrPointer_PTR24), .ZN(_03640_) );
  AND2_X1 U16647 ( .A1(_02745__PTR27), .A2(P1_P1_InstAddrPointer_PTR26), .ZN(_03641_) );
  AND2_X1 U16648 ( .A1(_02745__PTR29), .A2(P1_P1_InstAddrPointer_PTR28), .ZN(_03642_) );
  AND2_X1 U16649 ( .A1(_02743__PTR31), .A2(P1_P1_InstAddrPointer_PTR30), .ZN(_03643_) );
  AND2_X1 U16650 ( .A1(_03660_), .A2(_03685_), .ZN(_03645_) );
  AND2_X1 U16651 ( .A1(_03662_), .A2(_03687_), .ZN(_03646_) );
  AND2_X1 U16652 ( .A1(_03664_), .A2(_03689_), .ZN(_03647_) );
  AND2_X1 U16653 ( .A1(_03666_), .A2(_03691_), .ZN(_03648_) );
  AND2_X1 U16654 ( .A1(_03668_), .A2(_03693_), .ZN(_03649_) );
  AND2_X1 U16655 ( .A1(_03670_), .A2(_03695_), .ZN(_03650_) );
  AND2_X1 U16656 ( .A1(_03672_), .A2(_03697_), .ZN(_03651_) );
  AND2_X1 U16657 ( .A1(_03673_), .A2(_02744__PTR3), .ZN(_03652_) );
  AND2_X1 U16658 ( .A1(_03675_), .A2(_03699_), .ZN(_03653_) );
  AND2_X1 U16659 ( .A1(_03677_), .A2(_03701_), .ZN(_03654_) );
  AND2_X1 U16660 ( .A1(_03679_), .A2(_03703_), .ZN(_03655_) );
  AND2_X1 U16661 ( .A1(_03680_), .A2(_02744__PTR7), .ZN(_03656_) );
  AND2_X1 U16662 ( .A1(_03682_), .A2(_03706_), .ZN(_03657_) );
  AND2_X1 U16663 ( .A1(_03683_), .A2(_02744__PTR15), .ZN(_03658_) );
  AND2_X1 U16664 ( .A1(_02745__PTR3), .A2(_02745__PTR2), .ZN(_03644_) );
  AND2_X1 U16665 ( .A1(_02745__PTR5), .A2(_02745__PTR4), .ZN(_03659_) );
  AND2_X1 U16666 ( .A1(_02745__PTR7), .A2(_02745__PTR6), .ZN(_03660_) );
  AND2_X1 U16667 ( .A1(_02745__PTR9), .A2(_02745__PTR8), .ZN(_03661_) );
  AND2_X1 U16668 ( .A1(_02745__PTR11), .A2(_02745__PTR10), .ZN(_03662_) );
  AND2_X1 U16669 ( .A1(_02745__PTR13), .A2(_02745__PTR12), .ZN(_03663_) );
  AND2_X1 U16670 ( .A1(_02745__PTR15), .A2(_02745__PTR14), .ZN(_03664_) );
  AND2_X1 U16671 ( .A1(_02745__PTR17), .A2(_02745__PTR16), .ZN(_03665_) );
  AND2_X1 U16672 ( .A1(_02745__PTR19), .A2(_02745__PTR18), .ZN(_03666_) );
  AND2_X1 U16673 ( .A1(_02745__PTR21), .A2(_02745__PTR20), .ZN(_03667_) );
  AND2_X1 U16674 ( .A1(_02745__PTR23), .A2(_02745__PTR22), .ZN(_03668_) );
  AND2_X1 U16675 ( .A1(_02745__PTR25), .A2(_02745__PTR24), .ZN(_03669_) );
  AND2_X1 U16676 ( .A1(_02745__PTR27), .A2(_02745__PTR26), .ZN(_03670_) );
  AND2_X1 U16677 ( .A1(_02745__PTR29), .A2(_02745__PTR28), .ZN(_03671_) );
  AND2_X1 U16678 ( .A1(_02743__PTR31), .A2(_02745__PTR30), .ZN(_03672_) );
  AND2_X1 U16679 ( .A1(_03660_), .A2(_03659_), .ZN(_03673_) );
  AND2_X1 U16680 ( .A1(_03662_), .A2(_03661_), .ZN(_03674_) );
  AND2_X1 U16681 ( .A1(_03664_), .A2(_03663_), .ZN(_03675_) );
  AND2_X1 U16682 ( .A1(_03666_), .A2(_03665_), .ZN(_03676_) );
  AND2_X1 U16683 ( .A1(_03668_), .A2(_03667_), .ZN(_03677_) );
  AND2_X1 U16684 ( .A1(_03670_), .A2(_03669_), .ZN(_03678_) );
  AND2_X1 U16685 ( .A1(_03672_), .A2(_03671_), .ZN(_03679_) );
  AND2_X1 U16686 ( .A1(_03675_), .A2(_03674_), .ZN(_03680_) );
  AND2_X1 U16687 ( .A1(_03677_), .A2(_03676_), .ZN(_03681_) );
  AND2_X1 U16688 ( .A1(_03679_), .A2(_03678_), .ZN(_03682_) );
  AND2_X1 U16689 ( .A1(_03682_), .A2(_03681_), .ZN(_03683_) );
  OR2_X1 U16690 ( .A1(P1_P1_InstAddrPointer_PTR3), .A2(_03629_), .ZN(_03684_) );
  OR2_X1 U16691 ( .A1(P1_P1_InstAddrPointer_PTR5), .A2(_03630_), .ZN(_03685_) );
  OR2_X1 U16692 ( .A1(P1_P1_InstAddrPointer_PTR7), .A2(_03631_), .ZN(_03686_) );
  OR2_X1 U16693 ( .A1(P1_P1_InstAddrPointer_PTR9), .A2(_03632_), .ZN(_03687_) );
  OR2_X1 U16694 ( .A1(P1_P1_InstAddrPointer_PTR11), .A2(_03633_), .ZN(_03688_) );
  OR2_X1 U16695 ( .A1(P1_P1_InstAddrPointer_PTR13), .A2(_03634_), .ZN(_03689_) );
  OR2_X1 U16696 ( .A1(P1_P1_InstAddrPointer_PTR15), .A2(_03635_), .ZN(_03690_) );
  OR2_X1 U16697 ( .A1(P1_P1_InstAddrPointer_PTR17), .A2(_03636_), .ZN(_03691_) );
  OR2_X1 U16698 ( .A1(P1_P1_InstAddrPointer_PTR19), .A2(_03637_), .ZN(_03692_) );
  OR2_X1 U16699 ( .A1(P1_P1_InstAddrPointer_PTR21), .A2(_03638_), .ZN(_03693_) );
  OR2_X1 U16700 ( .A1(P1_P1_InstAddrPointer_PTR23), .A2(_03639_), .ZN(_03694_) );
  OR2_X1 U16701 ( .A1(P1_P1_InstAddrPointer_PTR25), .A2(_03640_), .ZN(_03695_) );
  OR2_X1 U16702 ( .A1(P1_P1_InstAddrPointer_PTR27), .A2(_03641_), .ZN(_03696_) );
  OR2_X1 U16703 ( .A1(P1_P1_InstAddrPointer_PTR29), .A2(_03642_), .ZN(_03697_) );
  OR2_X1 U16704 ( .A1(_03684_), .A2(_03644_), .ZN(_02744__PTR3) );
  OR2_X1 U16705 ( .A1(_03686_), .A2(_03645_), .ZN(_03698_) );
  OR2_X1 U16706 ( .A1(_03688_), .A2(_03646_), .ZN(_03699_) );
  OR2_X1 U16707 ( .A1(_03690_), .A2(_03647_), .ZN(_03700_) );
  OR2_X1 U16708 ( .A1(_03692_), .A2(_03648_), .ZN(_03701_) );
  OR2_X1 U16709 ( .A1(_03694_), .A2(_03649_), .ZN(_03702_) );
  OR2_X1 U16710 ( .A1(_03696_), .A2(_03650_), .ZN(_03703_) );
  OR2_X1 U16711 ( .A1(_03643_), .A2(_03651_), .ZN(_03704_) );
  OR2_X1 U16712 ( .A1(_03698_), .A2(_03652_), .ZN(_02744__PTR7) );
  OR2_X1 U16713 ( .A1(_03700_), .A2(_03653_), .ZN(_03705_) );
  OR2_X1 U16714 ( .A1(_03702_), .A2(_03654_), .ZN(_03706_) );
  OR2_X1 U16715 ( .A1(_03704_), .A2(_03655_), .ZN(_03707_) );
  OR2_X1 U16716 ( .A1(_03705_), .A2(_03656_), .ZN(_02744__PTR15) );
  OR2_X1 U16717 ( .A1(_03707_), .A2(_03657_), .ZN(_03708_) );
  OR2_X1 U16718 ( .A1(_03708_), .A2(_03658_), .ZN(_02744__PTR31) );
  AND2_X1 U16719 ( .A1(_01932__PTR43), .A2(_01932__PTR42), .ZN(_04087_) );
  AND2_X1 U16720 ( .A1(_02941__PTR4), .A2(_02942__PTR3), .ZN(_02740__PTR5) );
  OR2_X1 U16721 ( .A1(_02741__PTR3), .A2(_04087_), .ZN(_02942__PTR3) );
  AND2_X1 U16722 ( .A1(_02740__PTR5), .A2(_02739__PTR4), .ZN(_03625_) );
  AND2_X1 U16723 ( .A1(_01932__PTR43), .A2(_02739__PTR2), .ZN(_03626_) );
  AND2_X1 U16724 ( .A1(_02740__PTR5), .A2(_02742__PTR4), .ZN(_03627_) );
  AND2_X1 U16725 ( .A1(_03627_), .A2(_02741__PTR3), .ZN(_03628_) );
  OR2_X1 U16726 ( .A1(_02739__PTR3), .A2(_03626_), .ZN(_02741__PTR3) );
  OR2_X1 U16727 ( .A1(_03625_), .A2(_03628_), .ZN(_02741__PTR5) );
  AND2_X1 U16728 ( .A1(_02737__PTR1), .A2(_02736__PTR0), .ZN(_03619_) );
  AND2_X1 U16729 ( .A1(_02737__PTR3), .A2(_02738__PTR2), .ZN(_03620_) );
  AND2_X1 U16730 ( .A1(_03622_), .A2(_02736__PTR1), .ZN(_03621_) );
  AND2_X1 U16731 ( .A1(_02737__PTR3), .A2(_02737__PTR2), .ZN(_03622_) );
  AND2_X1 U16732 ( .A1(_02737__PTR4), .A2(_02736__PTR3), .ZN(_03623_) );
  OR2_X1 U16733 ( .A1(_02738__PTR0), .A2(_02737__PTR0), .ZN(_02736__PTR0) );
  OR2_X1 U16734 ( .A1(_02738__PTR1), .A2(_03619_), .ZN(_02736__PTR1) );
  OR2_X1 U16735 ( .A1(_02738__PTR3), .A2(_03620_), .ZN(_03624_) );
  OR2_X1 U16736 ( .A1(_03624_), .A2(_03621_), .ZN(_02736__PTR3) );
  OR2_X1 U16737 ( .A1(_02738__PTR4), .A2(_03623_), .ZN(_02736__PTR4) );
  AND2_X1 U16738 ( .A1(P1_EBX_PTR1), .A2(P1_EBX_PTR0), .ZN(_02828__PTR1) );
  AND2_X1 U16739 ( .A1(_03955_), .A2(_02828__PTR1), .ZN(_02828__PTR3) );
  AND2_X1 U16740 ( .A1(_03969_), .A2(_02828__PTR3), .ZN(_02828__PTR7) );
  AND2_X1 U16741 ( .A1(_03975_), .A2(_02828__PTR7), .ZN(_02828__PTR15) );
  AND2_X1 U16742 ( .A1(P1_EBX_PTR3), .A2(P1_EBX_PTR2), .ZN(_03955_) );
  AND2_X1 U16743 ( .A1(P1_EBX_PTR5), .A2(P1_EBX_PTR4), .ZN(_03956_) );
  AND2_X1 U16744 ( .A1(P1_EBX_PTR7), .A2(P1_EBX_PTR6), .ZN(_03957_) );
  AND2_X1 U16745 ( .A1(P1_EBX_PTR9), .A2(P1_EBX_PTR8), .ZN(_03958_) );
  AND2_X1 U16746 ( .A1(P1_EBX_PTR11), .A2(P1_EBX_PTR10), .ZN(_03959_) );
  AND2_X1 U16747 ( .A1(P1_EBX_PTR13), .A2(P1_EBX_PTR12), .ZN(_03960_) );
  AND2_X1 U16748 ( .A1(P1_EBX_PTR15), .A2(P1_EBX_PTR14), .ZN(_03961_) );
  AND2_X1 U16749 ( .A1(P1_EBX_PTR17), .A2(P1_EBX_PTR16), .ZN(_03962_) );
  AND2_X1 U16750 ( .A1(P1_EBX_PTR19), .A2(P1_EBX_PTR18), .ZN(_03963_) );
  AND2_X1 U16751 ( .A1(P1_EBX_PTR21), .A2(P1_EBX_PTR20), .ZN(_03964_) );
  AND2_X1 U16752 ( .A1(P1_EBX_PTR23), .A2(P1_EBX_PTR22), .ZN(_03965_) );
  AND2_X1 U16753 ( .A1(P1_EBX_PTR25), .A2(P1_EBX_PTR24), .ZN(_03966_) );
  AND2_X1 U16754 ( .A1(P1_EBX_PTR27), .A2(P1_EBX_PTR26), .ZN(_03967_) );
  AND2_X1 U16755 ( .A1(P1_EBX_PTR29), .A2(P1_EBX_PTR28), .ZN(_03968_) );
  AND2_X1 U16756 ( .A1(_03957_), .A2(_03956_), .ZN(_03969_) );
  AND2_X1 U16757 ( .A1(_03959_), .A2(_03958_), .ZN(_03970_) );
  AND2_X1 U16758 ( .A1(_03961_), .A2(_03960_), .ZN(_03971_) );
  AND2_X1 U16759 ( .A1(_03963_), .A2(_03962_), .ZN(_03972_) );
  AND2_X1 U16760 ( .A1(_03965_), .A2(_03964_), .ZN(_03973_) );
  AND2_X1 U16761 ( .A1(_03967_), .A2(_03966_), .ZN(_03974_) );
  AND2_X1 U16762 ( .A1(_03971_), .A2(_03970_), .ZN(_03975_) );
  AND2_X1 U16763 ( .A1(_03973_), .A2(_03972_), .ZN(_03976_) );
  AND2_X1 U16764 ( .A1(_03976_), .A2(_02828__PTR15), .ZN(_02828__PTR23) );
  AND2_X1 U16765 ( .A1(_03970_), .A2(_02828__PTR7), .ZN(_02828__PTR11) );
  AND2_X1 U16766 ( .A1(_03972_), .A2(_02828__PTR15), .ZN(_02828__PTR19) );
  AND2_X1 U16767 ( .A1(_03974_), .A2(_02828__PTR23), .ZN(_02828__PTR27) );
  AND2_X1 U16768 ( .A1(_03956_), .A2(_02828__PTR3), .ZN(_02828__PTR5) );
  AND2_X1 U16769 ( .A1(_03958_), .A2(_02828__PTR7), .ZN(_02828__PTR9) );
  AND2_X1 U16770 ( .A1(_03960_), .A2(_02828__PTR11), .ZN(_02828__PTR13) );
  AND2_X1 U16771 ( .A1(_03962_), .A2(_02828__PTR15), .ZN(_02828__PTR17) );
  AND2_X1 U16772 ( .A1(_03964_), .A2(_02828__PTR19), .ZN(_02828__PTR21) );
  AND2_X1 U16773 ( .A1(_03966_), .A2(_02828__PTR23), .ZN(_02828__PTR25) );
  AND2_X1 U16774 ( .A1(_03968_), .A2(_02828__PTR27), .ZN(_02828__PTR29) );
  AND2_X1 U16775 ( .A1(P1_EBX_PTR2), .A2(_02828__PTR1), .ZN(_02828__PTR2) );
  AND2_X1 U16776 ( .A1(P1_EBX_PTR4), .A2(_02828__PTR3), .ZN(_02828__PTR4) );
  AND2_X1 U16777 ( .A1(P1_EBX_PTR6), .A2(_02828__PTR5), .ZN(_02828__PTR6) );
  AND2_X1 U16778 ( .A1(P1_EBX_PTR8), .A2(_02828__PTR7), .ZN(_02828__PTR8) );
  AND2_X1 U16779 ( .A1(P1_EBX_PTR10), .A2(_02828__PTR9), .ZN(_02828__PTR10) );
  AND2_X1 U16780 ( .A1(P1_EBX_PTR12), .A2(_02828__PTR11), .ZN(_02828__PTR12) );
  AND2_X1 U16781 ( .A1(P1_EBX_PTR14), .A2(_02828__PTR13), .ZN(_02828__PTR14) );
  AND2_X1 U16782 ( .A1(P1_EBX_PTR16), .A2(_02828__PTR15), .ZN(_02828__PTR16) );
  AND2_X1 U16783 ( .A1(P1_EBX_PTR18), .A2(_02828__PTR17), .ZN(_02828__PTR18) );
  AND2_X1 U16784 ( .A1(P1_EBX_PTR20), .A2(_02828__PTR19), .ZN(_02828__PTR20) );
  AND2_X1 U16785 ( .A1(P1_EBX_PTR22), .A2(_02828__PTR21), .ZN(_02828__PTR22) );
  AND2_X1 U16786 ( .A1(P1_EBX_PTR24), .A2(_02828__PTR23), .ZN(_02828__PTR24) );
  AND2_X1 U16787 ( .A1(P1_EBX_PTR26), .A2(_02828__PTR25), .ZN(_02828__PTR26) );
  AND2_X1 U16788 ( .A1(P1_EBX_PTR28), .A2(_02828__PTR27), .ZN(_02828__PTR28) );
  AND2_X1 U16789 ( .A1(P1_EBX_PTR30), .A2(_02828__PTR29), .ZN(_02828__PTR30) );
  AND2_X1 U16790 ( .A1(P1_EAX_PTR1), .A2(P1_EAX_PTR0), .ZN(_02827__PTR1) );
  AND2_X1 U16791 ( .A1(_03941_), .A2(_02827__PTR1), .ZN(_02827__PTR3) );
  AND2_X1 U16792 ( .A1(_03949_), .A2(_02827__PTR3), .ZN(_02827__PTR7) );
  AND2_X1 U16793 ( .A1(_03953_), .A2(_02827__PTR7), .ZN(_02827__PTR15) );
  AND2_X1 U16794 ( .A1(P1_EAX_PTR3), .A2(P1_EAX_PTR2), .ZN(_03941_) );
  AND2_X1 U16795 ( .A1(P1_EAX_PTR5), .A2(P1_EAX_PTR4), .ZN(_03942_) );
  AND2_X1 U16796 ( .A1(P1_EAX_PTR7), .A2(P1_EAX_PTR6), .ZN(_03943_) );
  AND2_X1 U16797 ( .A1(P1_EAX_PTR9), .A2(P1_EAX_PTR8), .ZN(_03944_) );
  AND2_X1 U16798 ( .A1(P1_EAX_PTR11), .A2(P1_EAX_PTR10), .ZN(_03945_) );
  AND2_X1 U16799 ( .A1(P1_EAX_PTR13), .A2(P1_EAX_PTR12), .ZN(_03946_) );
  AND2_X1 U16800 ( .A1(P1_EAX_PTR15), .A2(P1_EAX_PTR14), .ZN(_03947_) );
  AND2_X1 U16801 ( .A1(P1_EAX_PTR17), .A2(P1_EAX_PTR16), .ZN(_03948_) );
  AND2_X1 U16802 ( .A1(_03943_), .A2(_03942_), .ZN(_03949_) );
  AND2_X1 U16803 ( .A1(_03945_), .A2(_03944_), .ZN(_03950_) );
  AND2_X1 U16804 ( .A1(_03947_), .A2(_03946_), .ZN(_03951_) );
  AND2_X1 U16805 ( .A1(_03933_), .A2(_03948_), .ZN(_03952_) );
  AND2_X1 U16806 ( .A1(_03951_), .A2(_03950_), .ZN(_03953_) );
  AND2_X1 U16807 ( .A1(_03939_), .A2(_03952_), .ZN(_03954_) );
  AND2_X1 U16808 ( .A1(_03954_), .A2(_02827__PTR15), .ZN(_02827__PTR23) );
  AND2_X1 U16809 ( .A1(_03950_), .A2(_02827__PTR7), .ZN(_02827__PTR11) );
  AND2_X1 U16810 ( .A1(_03952_), .A2(_02827__PTR15), .ZN(_02827__PTR19) );
  AND2_X1 U16811 ( .A1(_03940_), .A2(_02827__PTR23), .ZN(_02827__PTR27) );
  AND2_X1 U16812 ( .A1(_03942_), .A2(_02827__PTR3), .ZN(_02827__PTR5) );
  AND2_X1 U16813 ( .A1(_03944_), .A2(_02827__PTR7), .ZN(_02827__PTR9) );
  AND2_X1 U16814 ( .A1(_03946_), .A2(_02827__PTR11), .ZN(_02827__PTR13) );
  AND2_X1 U16815 ( .A1(_03948_), .A2(_02827__PTR15), .ZN(_02827__PTR17) );
  AND2_X1 U16816 ( .A1(_03934_), .A2(_02827__PTR19), .ZN(_02827__PTR21) );
  AND2_X1 U16817 ( .A1(_03936_), .A2(_02827__PTR23), .ZN(_02827__PTR25) );
  AND2_X1 U16818 ( .A1(_03938_), .A2(_02827__PTR27), .ZN(_02827__PTR29) );
  AND2_X1 U16819 ( .A1(P1_EAX_PTR2), .A2(_02827__PTR1), .ZN(_02827__PTR2) );
  AND2_X1 U16820 ( .A1(P1_EAX_PTR4), .A2(_02827__PTR3), .ZN(_02827__PTR4) );
  AND2_X1 U16821 ( .A1(P1_EAX_PTR6), .A2(_02827__PTR5), .ZN(_02827__PTR6) );
  AND2_X1 U16822 ( .A1(P1_EAX_PTR8), .A2(_02827__PTR7), .ZN(_02827__PTR8) );
  AND2_X1 U16823 ( .A1(P1_EAX_PTR10), .A2(_02827__PTR9), .ZN(_02827__PTR10) );
  AND2_X1 U16824 ( .A1(P1_EAX_PTR12), .A2(_02827__PTR11), .ZN(_02827__PTR12) );
  AND2_X1 U16825 ( .A1(P1_EAX_PTR14), .A2(_02827__PTR13), .ZN(_02827__PTR14) );
  AND2_X1 U16826 ( .A1(P1_EAX_PTR16), .A2(_02827__PTR15), .ZN(_02827__PTR16) );
  AND2_X1 U16827 ( .A1(P1_EAX_PTR18), .A2(_02827__PTR17), .ZN(_02827__PTR18) );
  AND2_X1 U16828 ( .A1(P1_EAX_PTR20), .A2(_02827__PTR19), .ZN(_02827__PTR20) );
  AND2_X1 U16829 ( .A1(P1_EAX_PTR22), .A2(_02827__PTR21), .ZN(_02827__PTR22) );
  AND2_X1 U16830 ( .A1(P1_EAX_PTR24), .A2(_02827__PTR23), .ZN(_02827__PTR24) );
  AND2_X1 U16831 ( .A1(P1_EAX_PTR26), .A2(_02827__PTR25), .ZN(_02827__PTR26) );
  AND2_X1 U16832 ( .A1(P1_EAX_PTR28), .A2(_02827__PTR27), .ZN(_02827__PTR28) );
  AND2_X1 U16833 ( .A1(P1_EAX_PTR30), .A2(_02827__PTR29), .ZN(_02827__PTR30) );
  AND2_X1 U16834 ( .A1(P1_EAX_PTR17), .A2(_02824__PTR0), .ZN(_02824__PTR1) );
  AND2_X1 U16835 ( .A1(_03933_), .A2(_02824__PTR1), .ZN(_02824__PTR3) );
  AND2_X1 U16836 ( .A1(_03939_), .A2(_02824__PTR3), .ZN(_02824__PTR7) );
  AND2_X1 U16837 ( .A1(P1_EAX_PTR19), .A2(P1_EAX_PTR18), .ZN(_03933_) );
  AND2_X1 U16838 ( .A1(P1_EAX_PTR21), .A2(P1_EAX_PTR20), .ZN(_03934_) );
  AND2_X1 U16839 ( .A1(P1_EAX_PTR23), .A2(P1_EAX_PTR22), .ZN(_03935_) );
  AND2_X1 U16840 ( .A1(P1_EAX_PTR25), .A2(P1_EAX_PTR24), .ZN(_03936_) );
  AND2_X1 U16841 ( .A1(P1_EAX_PTR27), .A2(P1_EAX_PTR26), .ZN(_03937_) );
  AND2_X1 U16842 ( .A1(P1_EAX_PTR29), .A2(P1_EAX_PTR28), .ZN(_03938_) );
  AND2_X1 U16843 ( .A1(_03935_), .A2(_03934_), .ZN(_03939_) );
  AND2_X1 U16844 ( .A1(_03937_), .A2(_03936_), .ZN(_03940_) );
  AND2_X1 U16845 ( .A1(_03940_), .A2(_02824__PTR7), .ZN(_02824__PTR11) );
  AND2_X1 U16846 ( .A1(_03934_), .A2(_02824__PTR3), .ZN(_02824__PTR5) );
  AND2_X1 U16847 ( .A1(_03936_), .A2(_02824__PTR7), .ZN(_02824__PTR9) );
  AND2_X1 U16848 ( .A1(_03938_), .A2(_02824__PTR11), .ZN(_02824__PTR13) );
  AND2_X1 U16849 ( .A1(P1_EAX_PTR18), .A2(_02824__PTR1), .ZN(_02824__PTR2) );
  AND2_X1 U16850 ( .A1(P1_EAX_PTR20), .A2(_02824__PTR3), .ZN(_02824__PTR4) );
  AND2_X1 U16851 ( .A1(P1_EAX_PTR22), .A2(_02824__PTR5), .ZN(_02824__PTR6) );
  AND2_X1 U16852 ( .A1(P1_EAX_PTR24), .A2(_02824__PTR7), .ZN(_02824__PTR8) );
  AND2_X1 U16853 ( .A1(P1_EAX_PTR26), .A2(_02824__PTR9), .ZN(_02824__PTR10) );
  AND2_X1 U16854 ( .A1(P1_EAX_PTR28), .A2(_02824__PTR11), .ZN(_02824__PTR12) );
  AND2_X1 U16855 ( .A1(P1_rEIP_PTR2), .A2(P1_rEIP_PTR1), .ZN(_02821__PTR1) );
  AND2_X1 U16856 ( .A1(_03716_), .A2(_02821__PTR1), .ZN(_02821__PTR3) );
  AND2_X1 U16857 ( .A1(_03730_), .A2(_02821__PTR3), .ZN(_02821__PTR7) );
  AND2_X1 U16858 ( .A1(_03736_), .A2(_02821__PTR7), .ZN(_02821__PTR15) );
  AND2_X1 U16859 ( .A1(P1_rEIP_PTR4), .A2(P1_rEIP_PTR3), .ZN(_03716_) );
  AND2_X1 U16860 ( .A1(P1_rEIP_PTR6), .A2(P1_rEIP_PTR5), .ZN(_03717_) );
  AND2_X1 U16861 ( .A1(P1_rEIP_PTR8), .A2(P1_rEIP_PTR7), .ZN(_03718_) );
  AND2_X1 U16862 ( .A1(P1_rEIP_PTR10), .A2(P1_rEIP_PTR9), .ZN(_03719_) );
  AND2_X1 U16863 ( .A1(P1_rEIP_PTR12), .A2(P1_rEIP_PTR11), .ZN(_03720_) );
  AND2_X1 U16864 ( .A1(P1_rEIP_PTR14), .A2(P1_rEIP_PTR13), .ZN(_03721_) );
  AND2_X1 U16865 ( .A1(P1_rEIP_PTR16), .A2(P1_rEIP_PTR15), .ZN(_03722_) );
  AND2_X1 U16866 ( .A1(P1_rEIP_PTR18), .A2(P1_rEIP_PTR17), .ZN(_03723_) );
  AND2_X1 U16867 ( .A1(P1_rEIP_PTR20), .A2(P1_rEIP_PTR19), .ZN(_03724_) );
  AND2_X1 U16868 ( .A1(P1_rEIP_PTR22), .A2(P1_rEIP_PTR21), .ZN(_03725_) );
  AND2_X1 U16869 ( .A1(P1_rEIP_PTR24), .A2(P1_rEIP_PTR23), .ZN(_03726_) );
  AND2_X1 U16870 ( .A1(P1_rEIP_PTR26), .A2(P1_rEIP_PTR25), .ZN(_03727_) );
  AND2_X1 U16871 ( .A1(P1_rEIP_PTR28), .A2(P1_rEIP_PTR27), .ZN(_03728_) );
  AND2_X1 U16872 ( .A1(P1_rEIP_PTR30), .A2(P1_rEIP_PTR29), .ZN(_03729_) );
  AND2_X1 U16873 ( .A1(_03722_), .A2(_03721_), .ZN(_03732_) );
  AND2_X1 U16874 ( .A1(_03724_), .A2(_03723_), .ZN(_03733_) );
  AND2_X1 U16875 ( .A1(_03726_), .A2(_03725_), .ZN(_03734_) );
  AND2_X1 U16876 ( .A1(_03737_), .A2(_02821__PTR15), .ZN(_02821__PTR23) );
  AND2_X1 U16877 ( .A1(_03731_), .A2(_02821__PTR7), .ZN(_02821__PTR11) );
  AND2_X1 U16878 ( .A1(_03733_), .A2(_02821__PTR15), .ZN(_02821__PTR19) );
  AND2_X1 U16879 ( .A1(_03735_), .A2(_02821__PTR23), .ZN(_02821__PTR27) );
  AND2_X1 U16880 ( .A1(_03717_), .A2(_02821__PTR3), .ZN(_02821__PTR5) );
  AND2_X1 U16881 ( .A1(_03719_), .A2(_02821__PTR7), .ZN(_02821__PTR9) );
  AND2_X1 U16882 ( .A1(_03721_), .A2(_02821__PTR11), .ZN(_02821__PTR13) );
  AND2_X1 U16883 ( .A1(_03723_), .A2(_02821__PTR15), .ZN(_02821__PTR17) );
  AND2_X1 U16884 ( .A1(_03725_), .A2(_02821__PTR19), .ZN(_02821__PTR21) );
  AND2_X1 U16885 ( .A1(_03727_), .A2(_02821__PTR23), .ZN(_02821__PTR25) );
  AND2_X1 U16886 ( .A1(_03729_), .A2(_02821__PTR27), .ZN(_02821__PTR29) );
  AND2_X1 U16887 ( .A1(P1_rEIP_PTR3), .A2(_02821__PTR1), .ZN(_02821__PTR2) );
  AND2_X1 U16888 ( .A1(P1_rEIP_PTR5), .A2(_02821__PTR3), .ZN(_02821__PTR4) );
  AND2_X1 U16889 ( .A1(P1_rEIP_PTR7), .A2(_02821__PTR5), .ZN(_02821__PTR6) );
  AND2_X1 U16890 ( .A1(P1_rEIP_PTR9), .A2(_02821__PTR7), .ZN(_02821__PTR8) );
  AND2_X1 U16891 ( .A1(P1_rEIP_PTR11), .A2(_02821__PTR9), .ZN(_02821__PTR10) );
  AND2_X1 U16892 ( .A1(P1_rEIP_PTR13), .A2(_02821__PTR11), .ZN(_02821__PTR12) );
  AND2_X1 U16893 ( .A1(P1_rEIP_PTR15), .A2(_02821__PTR13), .ZN(_02821__PTR14) );
  AND2_X1 U16894 ( .A1(P1_rEIP_PTR17), .A2(_02821__PTR15), .ZN(_02821__PTR16) );
  AND2_X1 U16895 ( .A1(P1_rEIP_PTR19), .A2(_02821__PTR17), .ZN(_02821__PTR18) );
  AND2_X1 U16896 ( .A1(P1_rEIP_PTR21), .A2(_02821__PTR19), .ZN(_02821__PTR20) );
  AND2_X1 U16897 ( .A1(P1_rEIP_PTR23), .A2(_02821__PTR21), .ZN(_02821__PTR22) );
  AND2_X1 U16898 ( .A1(P1_rEIP_PTR25), .A2(_02821__PTR23), .ZN(_02821__PTR24) );
  AND2_X1 U16899 ( .A1(P1_rEIP_PTR27), .A2(_02821__PTR25), .ZN(_02821__PTR26) );
  AND2_X1 U16900 ( .A1(P1_rEIP_PTR29), .A2(_02821__PTR27), .ZN(_02821__PTR28) );
  AND2_X1 U16901 ( .A1(_02734__PTR1), .A2(_02100__PTR32), .ZN(_02947__PTR1) );
  AND2_X1 U16902 ( .A1(_03554_), .A2(_02947__PTR1), .ZN(_02947__PTR3) );
  AND2_X1 U16903 ( .A1(_03583_), .A2(_02947__PTR3), .ZN(_02947__PTR7) );
  AND2_X1 U16904 ( .A1(_03590_), .A2(_02947__PTR7), .ZN(_02947__PTR15) );
  AND2_X1 U16905 ( .A1(_03591_), .A2(_02947__PTR15), .ZN(_02947__PTR23) );
  AND2_X1 U16906 ( .A1(_03584_), .A2(_02947__PTR7), .ZN(_02947__PTR11) );
  AND2_X1 U16907 ( .A1(_03586_), .A2(_02947__PTR15), .ZN(_02947__PTR19) );
  AND2_X1 U16908 ( .A1(_03588_), .A2(_02947__PTR23), .ZN(_02947__PTR27) );
  AND2_X1 U16909 ( .A1(_03569_), .A2(_02947__PTR3), .ZN(_02947__PTR5) );
  AND2_X1 U16910 ( .A1(_03571_), .A2(_02947__PTR7), .ZN(_02947__PTR9) );
  AND2_X1 U16911 ( .A1(_03573_), .A2(_02947__PTR11), .ZN(_02947__PTR13) );
  AND2_X1 U16912 ( .A1(_03575_), .A2(_02947__PTR15), .ZN(_02947__PTR17) );
  AND2_X1 U16913 ( .A1(_03577_), .A2(_02947__PTR19), .ZN(_02947__PTR21) );
  AND2_X1 U16914 ( .A1(_03579_), .A2(_02947__PTR23), .ZN(_02947__PTR25) );
  AND2_X1 U16915 ( .A1(_03581_), .A2(_02947__PTR27), .ZN(_02947__PTR29) );
  AND2_X1 U16916 ( .A1(_02734__PTR2), .A2(_02947__PTR1), .ZN(_02947__PTR2) );
  AND2_X1 U16917 ( .A1(_02734__PTR4), .A2(_02947__PTR3), .ZN(_02947__PTR4) );
  AND2_X1 U16918 ( .A1(_02734__PTR6), .A2(_02947__PTR5), .ZN(_02947__PTR6) );
  AND2_X1 U16919 ( .A1(_02734__PTR8), .A2(_02947__PTR7), .ZN(_02947__PTR8) );
  AND2_X1 U16920 ( .A1(_02734__PTR10), .A2(_02947__PTR9), .ZN(_02947__PTR10) );
  AND2_X1 U16921 ( .A1(_02734__PTR12), .A2(_02947__PTR11), .ZN(_02947__PTR12) );
  AND2_X1 U16922 ( .A1(_02734__PTR14), .A2(_02947__PTR13), .ZN(_02947__PTR14) );
  AND2_X1 U16923 ( .A1(_02734__PTR16), .A2(_02947__PTR15), .ZN(_02947__PTR16) );
  AND2_X1 U16924 ( .A1(_02734__PTR18), .A2(_02947__PTR17), .ZN(_02947__PTR18) );
  AND2_X1 U16925 ( .A1(_02734__PTR20), .A2(_02947__PTR19), .ZN(_02947__PTR20) );
  AND2_X1 U16926 ( .A1(_02734__PTR22), .A2(_02947__PTR21), .ZN(_02947__PTR22) );
  AND2_X1 U16927 ( .A1(_02734__PTR24), .A2(_02947__PTR23), .ZN(_02947__PTR24) );
  AND2_X1 U16928 ( .A1(_02734__PTR26), .A2(_02947__PTR25), .ZN(_02947__PTR26) );
  AND2_X1 U16929 ( .A1(_02734__PTR28), .A2(_02947__PTR27), .ZN(_02947__PTR28) );
  AND2_X1 U16930 ( .A1(_02734__PTR30), .A2(_02947__PTR29), .ZN(_02947__PTR30) );
  AND2_X1 U16931 ( .A1(_02734__PTR3), .A2(P1_EBX_PTR2), .ZN(_03539_) );
  AND2_X1 U16932 ( .A1(_02734__PTR5), .A2(P1_EBX_PTR4), .ZN(_03540_) );
  AND2_X1 U16933 ( .A1(_02734__PTR7), .A2(P1_EBX_PTR6), .ZN(_03541_) );
  AND2_X1 U16934 ( .A1(_02734__PTR9), .A2(P1_EBX_PTR8), .ZN(_03542_) );
  AND2_X1 U16935 ( .A1(_02734__PTR11), .A2(P1_EBX_PTR10), .ZN(_03543_) );
  AND2_X1 U16936 ( .A1(_02734__PTR13), .A2(P1_EBX_PTR12), .ZN(_03544_) );
  AND2_X1 U16937 ( .A1(_02734__PTR15), .A2(P1_EBX_PTR14), .ZN(_03545_) );
  AND2_X1 U16938 ( .A1(_02734__PTR17), .A2(P1_EBX_PTR16), .ZN(_03546_) );
  AND2_X1 U16939 ( .A1(_02734__PTR19), .A2(P1_EBX_PTR18), .ZN(_03547_) );
  AND2_X1 U16940 ( .A1(_02734__PTR21), .A2(P1_EBX_PTR20), .ZN(_03548_) );
  AND2_X1 U16941 ( .A1(_02734__PTR23), .A2(P1_EBX_PTR22), .ZN(_03549_) );
  AND2_X1 U16942 ( .A1(_02734__PTR25), .A2(P1_EBX_PTR24), .ZN(_03550_) );
  AND2_X1 U16943 ( .A1(_02734__PTR27), .A2(P1_EBX_PTR26), .ZN(_03551_) );
  AND2_X1 U16944 ( .A1(_02734__PTR29), .A2(P1_EBX_PTR28), .ZN(_03552_) );
  AND2_X1 U16945 ( .A1(_02732__PTR31), .A2(P1_EBX_PTR30), .ZN(_03553_) );
  AND2_X1 U16946 ( .A1(_03570_), .A2(_03595_), .ZN(_03555_) );
  AND2_X1 U16947 ( .A1(_03572_), .A2(_03597_), .ZN(_03556_) );
  AND2_X1 U16948 ( .A1(_03574_), .A2(_03599_), .ZN(_03557_) );
  AND2_X1 U16949 ( .A1(_03576_), .A2(_03601_), .ZN(_03558_) );
  AND2_X1 U16950 ( .A1(_03578_), .A2(_03603_), .ZN(_03559_) );
  AND2_X1 U16951 ( .A1(_03580_), .A2(_03605_), .ZN(_03560_) );
  AND2_X1 U16952 ( .A1(_03582_), .A2(_03607_), .ZN(_03561_) );
  AND2_X1 U16953 ( .A1(_03583_), .A2(_02733__PTR3), .ZN(_03562_) );
  AND2_X1 U16954 ( .A1(_03585_), .A2(_03609_), .ZN(_03563_) );
  AND2_X1 U16955 ( .A1(_03587_), .A2(_03611_), .ZN(_03564_) );
  AND2_X1 U16956 ( .A1(_03589_), .A2(_03613_), .ZN(_03565_) );
  AND2_X1 U16957 ( .A1(_03590_), .A2(_02733__PTR7), .ZN(_03566_) );
  AND2_X1 U16958 ( .A1(_03592_), .A2(_03616_), .ZN(_03567_) );
  AND2_X1 U16959 ( .A1(_03593_), .A2(_02733__PTR15), .ZN(_03568_) );
  AND2_X1 U16960 ( .A1(_02734__PTR3), .A2(_02734__PTR2), .ZN(_03554_) );
  AND2_X1 U16961 ( .A1(_02734__PTR5), .A2(_02734__PTR4), .ZN(_03569_) );
  AND2_X1 U16962 ( .A1(_02734__PTR7), .A2(_02734__PTR6), .ZN(_03570_) );
  AND2_X1 U16963 ( .A1(_02734__PTR9), .A2(_02734__PTR8), .ZN(_03571_) );
  AND2_X1 U16964 ( .A1(_02734__PTR11), .A2(_02734__PTR10), .ZN(_03572_) );
  AND2_X1 U16965 ( .A1(_02734__PTR13), .A2(_02734__PTR12), .ZN(_03573_) );
  AND2_X1 U16966 ( .A1(_02734__PTR15), .A2(_02734__PTR14), .ZN(_03574_) );
  AND2_X1 U16967 ( .A1(_02734__PTR17), .A2(_02734__PTR16), .ZN(_03575_) );
  AND2_X1 U16968 ( .A1(_02734__PTR19), .A2(_02734__PTR18), .ZN(_03576_) );
  AND2_X1 U16969 ( .A1(_02734__PTR21), .A2(_02734__PTR20), .ZN(_03577_) );
  AND2_X1 U16970 ( .A1(_02734__PTR23), .A2(_02734__PTR22), .ZN(_03578_) );
  AND2_X1 U16971 ( .A1(_02734__PTR25), .A2(_02734__PTR24), .ZN(_03579_) );
  AND2_X1 U16972 ( .A1(_02734__PTR27), .A2(_02734__PTR26), .ZN(_03580_) );
  AND2_X1 U16973 ( .A1(_02734__PTR29), .A2(_02734__PTR28), .ZN(_03581_) );
  AND2_X1 U16974 ( .A1(_02732__PTR31), .A2(_02734__PTR30), .ZN(_03582_) );
  AND2_X1 U16975 ( .A1(_03570_), .A2(_03569_), .ZN(_03583_) );
  AND2_X1 U16976 ( .A1(_03572_), .A2(_03571_), .ZN(_03584_) );
  AND2_X1 U16977 ( .A1(_03574_), .A2(_03573_), .ZN(_03585_) );
  AND2_X1 U16978 ( .A1(_03576_), .A2(_03575_), .ZN(_03586_) );
  AND2_X1 U16979 ( .A1(_03578_), .A2(_03577_), .ZN(_03587_) );
  AND2_X1 U16980 ( .A1(_03580_), .A2(_03579_), .ZN(_03588_) );
  AND2_X1 U16981 ( .A1(_03582_), .A2(_03581_), .ZN(_03589_) );
  AND2_X1 U16982 ( .A1(_03585_), .A2(_03584_), .ZN(_03590_) );
  AND2_X1 U16983 ( .A1(_03587_), .A2(_03586_), .ZN(_03591_) );
  AND2_X1 U16984 ( .A1(_03589_), .A2(_03588_), .ZN(_03592_) );
  AND2_X1 U16985 ( .A1(_03592_), .A2(_03591_), .ZN(_03593_) );
  OR2_X1 U16986 ( .A1(P1_EBX_PTR3), .A2(_03539_), .ZN(_03594_) );
  OR2_X1 U16987 ( .A1(P1_EBX_PTR5), .A2(_03540_), .ZN(_03595_) );
  OR2_X1 U16988 ( .A1(P1_EBX_PTR7), .A2(_03541_), .ZN(_03596_) );
  OR2_X1 U16989 ( .A1(P1_EBX_PTR9), .A2(_03542_), .ZN(_03597_) );
  OR2_X1 U16990 ( .A1(P1_EBX_PTR11), .A2(_03543_), .ZN(_03598_) );
  OR2_X1 U16991 ( .A1(P1_EBX_PTR13), .A2(_03544_), .ZN(_03599_) );
  OR2_X1 U16992 ( .A1(P1_EBX_PTR15), .A2(_03545_), .ZN(_03600_) );
  OR2_X1 U16993 ( .A1(P1_EBX_PTR17), .A2(_03546_), .ZN(_03601_) );
  OR2_X1 U16994 ( .A1(P1_EBX_PTR19), .A2(_03547_), .ZN(_03602_) );
  OR2_X1 U16995 ( .A1(P1_EBX_PTR21), .A2(_03548_), .ZN(_03603_) );
  OR2_X1 U16996 ( .A1(P1_EBX_PTR23), .A2(_03549_), .ZN(_03604_) );
  OR2_X1 U16997 ( .A1(P1_EBX_PTR25), .A2(_03550_), .ZN(_03605_) );
  OR2_X1 U16998 ( .A1(P1_EBX_PTR27), .A2(_03551_), .ZN(_03606_) );
  OR2_X1 U16999 ( .A1(P1_EBX_PTR29), .A2(_03552_), .ZN(_03607_) );
  OR2_X1 U17000 ( .A1(_03594_), .A2(_03554_), .ZN(_02733__PTR3) );
  OR2_X1 U17001 ( .A1(_03596_), .A2(_03555_), .ZN(_03608_) );
  OR2_X1 U17002 ( .A1(_03598_), .A2(_03556_), .ZN(_03609_) );
  OR2_X1 U17003 ( .A1(_03600_), .A2(_03557_), .ZN(_03610_) );
  OR2_X1 U17004 ( .A1(_03602_), .A2(_03558_), .ZN(_03611_) );
  OR2_X1 U17005 ( .A1(_03604_), .A2(_03559_), .ZN(_03612_) );
  OR2_X1 U17006 ( .A1(_03606_), .A2(_03560_), .ZN(_03613_) );
  OR2_X1 U17007 ( .A1(_03553_), .A2(_03561_), .ZN(_03614_) );
  OR2_X1 U17008 ( .A1(_03608_), .A2(_03562_), .ZN(_02733__PTR7) );
  OR2_X1 U17009 ( .A1(_03610_), .A2(_03563_), .ZN(_03615_) );
  OR2_X1 U17010 ( .A1(_03612_), .A2(_03564_), .ZN(_03616_) );
  OR2_X1 U17011 ( .A1(_03614_), .A2(_03565_), .ZN(_03617_) );
  OR2_X1 U17012 ( .A1(_03615_), .A2(_03566_), .ZN(_02733__PTR15) );
  OR2_X1 U17013 ( .A1(_03617_), .A2(_03567_), .ZN(_03618_) );
  OR2_X1 U17014 ( .A1(_03618_), .A2(_03568_), .ZN(_02733__PTR31) );
  AND2_X1 U17015 ( .A1(_02932__PTR1), .A2(_02931__PTR0), .ZN(_03977_) );
  AND2_X1 U17016 ( .A1(_02932__PTR3), .A2(_02933__PTR2), .ZN(_03978_) );
  AND2_X1 U17017 ( .A1(_03980_), .A2(_02931__PTR1), .ZN(_03979_) );
  AND2_X1 U17018 ( .A1(_02932__PTR3), .A2(_02932__PTR2), .ZN(_03980_) );
  AND2_X1 U17019 ( .A1(_02932__PTR2), .A2(_02931__PTR1), .ZN(_03982_) );
  AND2_X1 U17020 ( .A1(_02932__PTR4), .A2(_02931__PTR3), .ZN(_03981_) );
  OR2_X1 U17021 ( .A1(_02933__PTR0), .A2(_02718__PTR0), .ZN(_02931__PTR0) );
  OR2_X1 U17022 ( .A1(_02933__PTR1), .A2(_03977_), .ZN(_02931__PTR1) );
  OR2_X1 U17023 ( .A1(_02933__PTR3), .A2(_03978_), .ZN(_03983_) );
  OR2_X1 U17024 ( .A1(_03983_), .A2(_03979_), .ZN(_02931__PTR3) );
  OR2_X1 U17025 ( .A1(_02933__PTR4), .A2(_03981_), .ZN(_02720__PTR5) );
  OR2_X1 U17026 ( .A1(_02933__PTR2), .A2(_03982_), .ZN(_02931__PTR2) );
  AND2_X1 U17027 ( .A1(_02717__PTR1), .A2(_02718__PTR0), .ZN(_00618__PTR0) );
  AND2_X1 U17028 ( .A1(_02719__PTR3), .A2(_02729__PTR1), .ZN(_02729__PTR3) );
  AND2_X1 U17029 ( .A1(_00618__PTR2), .A2(_02729__PTR3), .ZN(_03538_) );
  OR2_X1 U17030 ( .A1(_02718__PTR1), .A2(_00618__PTR0), .ZN(_02729__PTR1) );
  OR2_X1 U17031 ( .A1(_02716__PTR5), .A2(_03538_), .ZN(_02729__PTR5) );
  AND2_X1 U17032 ( .A1(_01886__PTR5), .A2(_02750__PTR1), .ZN(_03932_) );
  OR2_X1 U17033 ( .A1(P1_P1_InstQueueRd_Addr_PTR2), .A2(_03932_), .ZN(_02819__PTR2) );
  AND2_X1 U17034 ( .A1(P1_P1_InstQueueRd_Addr_PTR2), .A2(P1_P1_InstQueueRd_Addr_PTR1), .ZN(_02817__PTR1) );
  AND2_X1 U17035 ( .A1(P1_P1_InstQueueRd_Addr_PTR3), .A2(_02817__PTR1), .ZN(_02817__PTR2) );
  AND2_X1 U17036 ( .A1(_01887__PTR1), .A2(_02814__PTR0), .ZN(_02814__PTR1) );
  AND2_X1 U17037 ( .A1(_03928_), .A2(_02814__PTR1), .ZN(_02814__PTR3) );
  AND2_X1 U17038 ( .A1(_03931_), .A2(_02814__PTR3), .ZN(_02814__PTR7) );
  AND2_X1 U17039 ( .A1(_01887__PTR3), .A2(_01887__PTR2), .ZN(_03928_) );
  AND2_X1 U17040 ( .A1(_01887__PTR5), .A2(_01887__PTR4), .ZN(_03929_) );
  AND2_X1 U17041 ( .A1(_01887__PTR7), .A2(_01887__PTR6), .ZN(_03930_) );
  AND2_X1 U17042 ( .A1(_03930_), .A2(_03929_), .ZN(_03931_) );
  AND2_X1 U17043 ( .A1(_03929_), .A2(_02814__PTR3), .ZN(_02814__PTR5) );
  AND2_X1 U17044 ( .A1(_01887__PTR2), .A2(_02814__PTR1), .ZN(_02814__PTR2) );
  AND2_X1 U17045 ( .A1(_01887__PTR4), .A2(_02814__PTR3), .ZN(_02814__PTR4) );
  AND2_X1 U17046 ( .A1(_01887__PTR6), .A2(_02814__PTR5), .ZN(_02814__PTR6) );
  AND2_X1 U17047 ( .A1(_01890__PTR4), .A2(P1_P1_InstQueueRd_Addr_PTR0), .ZN(_03927_) );
  AND2_X1 U17048 ( .A1(P1_P1_InstQueueRd_Addr_PTR2), .A2(_02813__PTR1), .ZN(_02813__PTR2) );
  OR2_X1 U17049 ( .A1(P1_P1_InstQueueRd_Addr_PTR1), .A2(_03927_), .ZN(_02813__PTR1) );
  AND2_X1 U17050 ( .A1(_03888_), .A2(_02798__PTR1), .ZN(_03887_) );
  AND2_X1 U17051 ( .A1(_03820_), .A2(_02806__PTR3), .ZN(_02806__PTR7) );
  AND2_X1 U17052 ( .A1(_03826_), .A2(_02806__PTR7), .ZN(_02806__PTR15) );
  AND2_X1 U17053 ( .A1(P1_P1_InstAddrPointer_PTR3), .A2(_02745__PTR2), .ZN(_03888_) );
  AND2_X1 U17054 ( .A1(_03808_), .A2(_03807_), .ZN(_03820_) );
  AND2_X1 U17055 ( .A1(_03810_), .A2(_03809_), .ZN(_03821_) );
  AND2_X1 U17056 ( .A1(_03812_), .A2(_03811_), .ZN(_03822_) );
  AND2_X1 U17057 ( .A1(_03814_), .A2(_03813_), .ZN(_03823_) );
  AND2_X1 U17058 ( .A1(_03816_), .A2(_03815_), .ZN(_03824_) );
  AND2_X1 U17059 ( .A1(_03818_), .A2(_03817_), .ZN(_03825_) );
  AND2_X1 U17060 ( .A1(_03822_), .A2(_03821_), .ZN(_03826_) );
  AND2_X1 U17061 ( .A1(_03824_), .A2(_03823_), .ZN(_03827_) );
  AND2_X1 U17062 ( .A1(_03827_), .A2(_02806__PTR15), .ZN(_02806__PTR23) );
  AND2_X1 U17063 ( .A1(_03821_), .A2(_02806__PTR7), .ZN(_02806__PTR11) );
  AND2_X1 U17064 ( .A1(_03823_), .A2(_02806__PTR15), .ZN(_02806__PTR19) );
  AND2_X1 U17065 ( .A1(_03825_), .A2(_02806__PTR23), .ZN(_02806__PTR27) );
  AND2_X1 U17066 ( .A1(_03807_), .A2(_02806__PTR3), .ZN(_02806__PTR5) );
  AND2_X1 U17067 ( .A1(_03809_), .A2(_02806__PTR7), .ZN(_02806__PTR9) );
  AND2_X1 U17068 ( .A1(_03811_), .A2(_02806__PTR11), .ZN(_02806__PTR13) );
  AND2_X1 U17069 ( .A1(_03813_), .A2(_02806__PTR15), .ZN(_02806__PTR17) );
  AND2_X1 U17070 ( .A1(_03815_), .A2(_02806__PTR19), .ZN(_02806__PTR21) );
  AND2_X1 U17071 ( .A1(_03817_), .A2(_02806__PTR23), .ZN(_02806__PTR25) );
  AND2_X1 U17072 ( .A1(_03819_), .A2(_02806__PTR27), .ZN(_02806__PTR29) );
  AND2_X1 U17073 ( .A1(_02745__PTR2), .A2(_02798__PTR1), .ZN(_03889_) );
  AND2_X1 U17074 ( .A1(P1_P1_InstAddrPointer_PTR4), .A2(_02806__PTR3), .ZN(_02806__PTR4) );
  AND2_X1 U17075 ( .A1(P1_P1_InstAddrPointer_PTR6), .A2(_02806__PTR5), .ZN(_02806__PTR6) );
  AND2_X1 U17076 ( .A1(P1_P1_InstAddrPointer_PTR8), .A2(_02806__PTR7), .ZN(_02806__PTR8) );
  AND2_X1 U17077 ( .A1(P1_P1_InstAddrPointer_PTR10), .A2(_02806__PTR9), .ZN(_02806__PTR10) );
  AND2_X1 U17078 ( .A1(P1_P1_InstAddrPointer_PTR12), .A2(_02806__PTR11), .ZN(_02806__PTR12) );
  AND2_X1 U17079 ( .A1(P1_P1_InstAddrPointer_PTR14), .A2(_02806__PTR13), .ZN(_02806__PTR14) );
  AND2_X1 U17080 ( .A1(P1_P1_InstAddrPointer_PTR16), .A2(_02806__PTR15), .ZN(_02806__PTR16) );
  AND2_X1 U17081 ( .A1(P1_P1_InstAddrPointer_PTR18), .A2(_02806__PTR17), .ZN(_02806__PTR18) );
  AND2_X1 U17082 ( .A1(P1_P1_InstAddrPointer_PTR20), .A2(_02806__PTR19), .ZN(_02806__PTR20) );
  AND2_X1 U17083 ( .A1(P1_P1_InstAddrPointer_PTR22), .A2(_02806__PTR21), .ZN(_02806__PTR22) );
  AND2_X1 U17084 ( .A1(P1_P1_InstAddrPointer_PTR24), .A2(_02806__PTR23), .ZN(_02806__PTR24) );
  AND2_X1 U17085 ( .A1(P1_P1_InstAddrPointer_PTR26), .A2(_02806__PTR25), .ZN(_02806__PTR26) );
  AND2_X1 U17086 ( .A1(P1_P1_InstAddrPointer_PTR28), .A2(_02806__PTR27), .ZN(_02806__PTR28) );
  AND2_X1 U17087 ( .A1(P1_P1_InstAddrPointer_PTR30), .A2(_02806__PTR29), .ZN(_02806__PTR30) );
  OR2_X1 U17088 ( .A1(_03806_), .A2(_03887_), .ZN(_02806__PTR3) );
  OR2_X1 U17089 ( .A1(P1_P1_InstAddrPointer_PTR2), .A2(_03889_), .ZN(_02806__PTR2) );
  AND2_X1 U17090 ( .A1(_02809__PTR1), .A2(_02808__PTR0), .ZN(_03890_) );
  AND2_X1 U17091 ( .A1(_02809__PTR3), .A2(_02811__PTR2), .ZN(_03891_) );
  AND2_X1 U17092 ( .A1(_02809__PTR5), .A2(_02811__PTR4), .ZN(_03892_) );
  AND2_X1 U17093 ( .A1(_02809__PTR7), .A2(_02811__PTR6), .ZN(_03893_) );
  AND2_X1 U17094 ( .A1(_03897_), .A2(_02808__PTR1), .ZN(_03894_) );
  AND2_X1 U17095 ( .A1(_03899_), .A2(_03924_), .ZN(_03895_) );
  AND2_X1 U17096 ( .A1(_03911_), .A2(_02808__PTR3), .ZN(_03896_) );
  AND2_X1 U17097 ( .A1(_03917_), .A2(_02808__PTR7), .ZN(_02808__PTR15) );
  AND2_X1 U17098 ( .A1(_02809__PTR3), .A2(_02809__PTR2), .ZN(_03897_) );
  AND2_X1 U17099 ( .A1(_02809__PTR5), .A2(_02809__PTR4), .ZN(_03898_) );
  AND2_X1 U17100 ( .A1(_02809__PTR7), .A2(_02809__PTR6), .ZN(_03899_) );
  AND2_X1 U17101 ( .A1(_02807__PTR9), .A2(_02807__PTR8), .ZN(_03900_) );
  AND2_X1 U17102 ( .A1(_02807__PTR11), .A2(_02807__PTR10), .ZN(_03901_) );
  AND2_X1 U17103 ( .A1(_02807__PTR13), .A2(_02807__PTR12), .ZN(_03902_) );
  AND2_X1 U17104 ( .A1(_02807__PTR15), .A2(_02807__PTR14), .ZN(_03903_) );
  AND2_X1 U17105 ( .A1(_02807__PTR17), .A2(_02807__PTR16), .ZN(_03904_) );
  AND2_X1 U17106 ( .A1(_02807__PTR19), .A2(_02807__PTR18), .ZN(_03905_) );
  AND2_X1 U17107 ( .A1(_02807__PTR21), .A2(_02807__PTR20), .ZN(_03906_) );
  AND2_X1 U17108 ( .A1(_02807__PTR23), .A2(_02807__PTR22), .ZN(_03907_) );
  AND2_X1 U17109 ( .A1(_02807__PTR25), .A2(_02807__PTR24), .ZN(_03908_) );
  AND2_X1 U17110 ( .A1(_02807__PTR27), .A2(_02807__PTR26), .ZN(_03909_) );
  AND2_X1 U17111 ( .A1(_02807__PTR29), .A2(_02807__PTR28), .ZN(_03910_) );
  AND2_X1 U17112 ( .A1(_03899_), .A2(_03898_), .ZN(_03911_) );
  AND2_X1 U17113 ( .A1(_03901_), .A2(_03900_), .ZN(_03912_) );
  AND2_X1 U17114 ( .A1(_03903_), .A2(_03902_), .ZN(_03913_) );
  AND2_X1 U17115 ( .A1(_03905_), .A2(_03904_), .ZN(_03914_) );
  AND2_X1 U17116 ( .A1(_03907_), .A2(_03906_), .ZN(_03915_) );
  AND2_X1 U17117 ( .A1(_03909_), .A2(_03908_), .ZN(_03916_) );
  AND2_X1 U17118 ( .A1(_03913_), .A2(_03912_), .ZN(_03917_) );
  AND2_X1 U17119 ( .A1(_03915_), .A2(_03914_), .ZN(_03918_) );
  AND2_X1 U17120 ( .A1(_03918_), .A2(_02808__PTR15), .ZN(_02808__PTR23) );
  AND2_X1 U17121 ( .A1(_03912_), .A2(_02808__PTR7), .ZN(_02808__PTR11) );
  AND2_X1 U17122 ( .A1(_03914_), .A2(_02808__PTR15), .ZN(_02808__PTR19) );
  AND2_X1 U17123 ( .A1(_03916_), .A2(_02808__PTR23), .ZN(_02808__PTR27) );
  AND2_X1 U17124 ( .A1(_03898_), .A2(_02808__PTR3), .ZN(_03919_) );
  AND2_X1 U17125 ( .A1(_03900_), .A2(_02808__PTR7), .ZN(_02808__PTR9) );
  AND2_X1 U17126 ( .A1(_03902_), .A2(_02808__PTR11), .ZN(_02808__PTR13) );
  AND2_X1 U17127 ( .A1(_03904_), .A2(_02808__PTR15), .ZN(_02808__PTR17) );
  AND2_X1 U17128 ( .A1(_03906_), .A2(_02808__PTR19), .ZN(_02808__PTR21) );
  AND2_X1 U17129 ( .A1(_03908_), .A2(_02808__PTR23), .ZN(_02808__PTR25) );
  AND2_X1 U17130 ( .A1(_03910_), .A2(_02808__PTR27), .ZN(_02808__PTR29) );
  AND2_X1 U17131 ( .A1(_02809__PTR2), .A2(_02808__PTR1), .ZN(_03920_) );
  AND2_X1 U17132 ( .A1(_02809__PTR4), .A2(_02808__PTR3), .ZN(_03921_) );
  AND2_X1 U17133 ( .A1(_02809__PTR6), .A2(_02808__PTR5), .ZN(_03922_) );
  AND2_X1 U17134 ( .A1(_02807__PTR8), .A2(_02808__PTR7), .ZN(_02808__PTR8) );
  AND2_X1 U17135 ( .A1(_02807__PTR10), .A2(_02808__PTR9), .ZN(_02808__PTR10) );
  AND2_X1 U17136 ( .A1(_02807__PTR12), .A2(_02808__PTR11), .ZN(_02808__PTR12) );
  AND2_X1 U17137 ( .A1(_02807__PTR14), .A2(_02808__PTR13), .ZN(_02808__PTR14) );
  AND2_X1 U17138 ( .A1(_02807__PTR16), .A2(_02808__PTR15), .ZN(_02808__PTR16) );
  AND2_X1 U17139 ( .A1(_02807__PTR18), .A2(_02808__PTR17), .ZN(_02808__PTR18) );
  AND2_X1 U17140 ( .A1(_02807__PTR20), .A2(_02808__PTR19), .ZN(_02808__PTR20) );
  AND2_X1 U17141 ( .A1(_02807__PTR22), .A2(_02808__PTR21), .ZN(_02808__PTR22) );
  AND2_X1 U17142 ( .A1(_02807__PTR24), .A2(_02808__PTR23), .ZN(_02808__PTR24) );
  AND2_X1 U17143 ( .A1(_02807__PTR26), .A2(_02808__PTR25), .ZN(_02808__PTR26) );
  AND2_X1 U17144 ( .A1(_02807__PTR28), .A2(_02808__PTR27), .ZN(_02808__PTR28) );
  AND2_X1 U17145 ( .A1(_02807__PTR30), .A2(_02808__PTR29), .ZN(_02808__PTR30) );
  OR2_X1 U17146 ( .A1(_02811__PTR1), .A2(_03890_), .ZN(_02808__PTR1) );
  OR2_X1 U17147 ( .A1(_02811__PTR3), .A2(_03891_), .ZN(_03923_) );
  OR2_X1 U17148 ( .A1(_02811__PTR5), .A2(_03892_), .ZN(_03924_) );
  OR2_X1 U17149 ( .A1(_02811__PTR7), .A2(_03893_), .ZN(_03925_) );
  OR2_X1 U17150 ( .A1(_03923_), .A2(_03894_), .ZN(_02808__PTR3) );
  OR2_X1 U17151 ( .A1(_03925_), .A2(_03895_), .ZN(_03926_) );
  OR2_X1 U17152 ( .A1(_03926_), .A2(_03896_), .ZN(_02808__PTR7) );
  OR2_X1 U17153 ( .A1(_03924_), .A2(_03919_), .ZN(_02808__PTR5) );
  OR2_X1 U17154 ( .A1(_02811__PTR2), .A2(_03920_), .ZN(_02808__PTR2) );
  OR2_X1 U17155 ( .A1(_02811__PTR4), .A2(_03921_), .ZN(_02808__PTR4) );
  OR2_X1 U17156 ( .A1(_02811__PTR6), .A2(_03922_), .ZN(_02808__PTR6) );
  AND2_X1 U17157 ( .A1(_00620__PTR1), .A2(_02718__PTR1), .ZN(_03536_) );
  AND2_X1 U17158 ( .A1(_02718__PTR3), .A2(_02717__PTR2), .ZN(_00620__PTR1) );
  AND2_X1 U17159 ( .A1(_00618__PTR2), .A2(_02726__PTR3), .ZN(_03537_) );
  OR2_X1 U17160 ( .A1(_02719__PTR3), .A2(_03536_), .ZN(_02726__PTR3) );
  OR2_X1 U17161 ( .A1(_02716__PTR5), .A2(_03537_), .ZN(_02726__PTR5) );
  AND2_X1 U17162 ( .A1(P1_P1_InstAddrPointer_PTR2), .A2(P1_P1_InstAddrPointer_PTR1), .ZN(_02801__PTR1) );
  AND2_X1 U17163 ( .A1(_03828_), .A2(_02801__PTR1), .ZN(_02801__PTR3) );
  AND2_X1 U17164 ( .A1(_03842_), .A2(_02801__PTR3), .ZN(_02801__PTR7) );
  AND2_X1 U17165 ( .A1(_03848_), .A2(_02801__PTR7), .ZN(_02801__PTR15) );
  AND2_X1 U17166 ( .A1(P1_P1_InstAddrPointer_PTR4), .A2(P1_P1_InstAddrPointer_PTR3), .ZN(_03828_) );
  AND2_X1 U17167 ( .A1(P1_P1_InstAddrPointer_PTR6), .A2(P1_P1_InstAddrPointer_PTR5), .ZN(_03829_) );
  AND2_X1 U17168 ( .A1(P1_P1_InstAddrPointer_PTR8), .A2(P1_P1_InstAddrPointer_PTR7), .ZN(_03830_) );
  AND2_X1 U17169 ( .A1(P1_P1_InstAddrPointer_PTR10), .A2(P1_P1_InstAddrPointer_PTR9), .ZN(_03831_) );
  AND2_X1 U17170 ( .A1(P1_P1_InstAddrPointer_PTR12), .A2(P1_P1_InstAddrPointer_PTR11), .ZN(_03832_) );
  AND2_X1 U17171 ( .A1(P1_P1_InstAddrPointer_PTR14), .A2(P1_P1_InstAddrPointer_PTR13), .ZN(_03833_) );
  AND2_X1 U17172 ( .A1(P1_P1_InstAddrPointer_PTR16), .A2(P1_P1_InstAddrPointer_PTR15), .ZN(_03834_) );
  AND2_X1 U17173 ( .A1(P1_P1_InstAddrPointer_PTR18), .A2(P1_P1_InstAddrPointer_PTR17), .ZN(_03835_) );
  AND2_X1 U17174 ( .A1(P1_P1_InstAddrPointer_PTR20), .A2(P1_P1_InstAddrPointer_PTR19), .ZN(_03836_) );
  AND2_X1 U17175 ( .A1(P1_P1_InstAddrPointer_PTR22), .A2(P1_P1_InstAddrPointer_PTR21), .ZN(_03837_) );
  AND2_X1 U17176 ( .A1(P1_P1_InstAddrPointer_PTR24), .A2(P1_P1_InstAddrPointer_PTR23), .ZN(_03838_) );
  AND2_X1 U17177 ( .A1(P1_P1_InstAddrPointer_PTR26), .A2(P1_P1_InstAddrPointer_PTR25), .ZN(_03839_) );
  AND2_X1 U17178 ( .A1(P1_P1_InstAddrPointer_PTR28), .A2(P1_P1_InstAddrPointer_PTR27), .ZN(_03840_) );
  AND2_X1 U17179 ( .A1(P1_P1_InstAddrPointer_PTR30), .A2(P1_P1_InstAddrPointer_PTR29), .ZN(_03841_) );
  AND2_X1 U17180 ( .A1(_03830_), .A2(_03829_), .ZN(_03842_) );
  AND2_X1 U17181 ( .A1(_03832_), .A2(_03831_), .ZN(_03843_) );
  AND2_X1 U17182 ( .A1(_03834_), .A2(_03833_), .ZN(_03844_) );
  AND2_X1 U17183 ( .A1(_03836_), .A2(_03835_), .ZN(_03845_) );
  AND2_X1 U17184 ( .A1(_03838_), .A2(_03837_), .ZN(_03846_) );
  AND2_X1 U17185 ( .A1(_03840_), .A2(_03839_), .ZN(_03847_) );
  AND2_X1 U17186 ( .A1(_03844_), .A2(_03843_), .ZN(_03848_) );
  AND2_X1 U17187 ( .A1(_03846_), .A2(_03845_), .ZN(_03849_) );
  AND2_X1 U17188 ( .A1(_03849_), .A2(_02801__PTR15), .ZN(_02801__PTR23) );
  AND2_X1 U17189 ( .A1(_03843_), .A2(_02801__PTR7), .ZN(_02801__PTR11) );
  AND2_X1 U17190 ( .A1(_03845_), .A2(_02801__PTR15), .ZN(_02801__PTR19) );
  AND2_X1 U17191 ( .A1(_03847_), .A2(_02801__PTR23), .ZN(_02801__PTR27) );
  AND2_X1 U17192 ( .A1(_03829_), .A2(_02801__PTR3), .ZN(_02801__PTR5) );
  AND2_X1 U17193 ( .A1(_03831_), .A2(_02801__PTR7), .ZN(_02801__PTR9) );
  AND2_X1 U17194 ( .A1(_03833_), .A2(_02801__PTR11), .ZN(_02801__PTR13) );
  AND2_X1 U17195 ( .A1(_03835_), .A2(_02801__PTR15), .ZN(_02801__PTR17) );
  AND2_X1 U17196 ( .A1(_03837_), .A2(_02801__PTR19), .ZN(_02801__PTR21) );
  AND2_X1 U17197 ( .A1(_03839_), .A2(_02801__PTR23), .ZN(_02801__PTR25) );
  AND2_X1 U17198 ( .A1(_03841_), .A2(_02801__PTR27), .ZN(_02801__PTR29) );
  AND2_X1 U17199 ( .A1(P1_P1_InstAddrPointer_PTR3), .A2(_02801__PTR1), .ZN(_02801__PTR2) );
  AND2_X1 U17200 ( .A1(P1_P1_InstAddrPointer_PTR5), .A2(_02801__PTR3), .ZN(_02801__PTR4) );
  AND2_X1 U17201 ( .A1(P1_P1_InstAddrPointer_PTR7), .A2(_02801__PTR5), .ZN(_02801__PTR6) );
  AND2_X1 U17202 ( .A1(P1_P1_InstAddrPointer_PTR9), .A2(_02801__PTR7), .ZN(_02801__PTR8) );
  AND2_X1 U17203 ( .A1(P1_P1_InstAddrPointer_PTR11), .A2(_02801__PTR9), .ZN(_02801__PTR10) );
  AND2_X1 U17204 ( .A1(P1_P1_InstAddrPointer_PTR13), .A2(_02801__PTR11), .ZN(_02801__PTR12) );
  AND2_X1 U17205 ( .A1(P1_P1_InstAddrPointer_PTR15), .A2(_02801__PTR13), .ZN(_02801__PTR14) );
  AND2_X1 U17206 ( .A1(P1_P1_InstAddrPointer_PTR17), .A2(_02801__PTR15), .ZN(_02801__PTR16) );
  AND2_X1 U17207 ( .A1(P1_P1_InstAddrPointer_PTR19), .A2(_02801__PTR17), .ZN(_02801__PTR18) );
  AND2_X1 U17208 ( .A1(P1_P1_InstAddrPointer_PTR21), .A2(_02801__PTR19), .ZN(_02801__PTR20) );
  AND2_X1 U17209 ( .A1(P1_P1_InstAddrPointer_PTR23), .A2(_02801__PTR21), .ZN(_02801__PTR22) );
  AND2_X1 U17210 ( .A1(P1_P1_InstAddrPointer_PTR25), .A2(_02801__PTR23), .ZN(_02801__PTR24) );
  AND2_X1 U17211 ( .A1(P1_P1_InstAddrPointer_PTR27), .A2(_02801__PTR25), .ZN(_02801__PTR26) );
  AND2_X1 U17212 ( .A1(P1_P1_InstAddrPointer_PTR29), .A2(_02801__PTR27), .ZN(_02801__PTR28) );
  AND2_X1 U17213 ( .A1(_02803__PTR1), .A2(_02802__PTR0), .ZN(_03850_) );
  AND2_X1 U17214 ( .A1(_02803__PTR3), .A2(_02805__PTR2), .ZN(_03851_) );
  AND2_X1 U17215 ( .A1(_02803__PTR5), .A2(_02805__PTR4), .ZN(_03852_) );
  AND2_X1 U17216 ( .A1(_02803__PTR7), .A2(_02805__PTR6), .ZN(_03853_) );
  AND2_X1 U17217 ( .A1(_03857_), .A2(_02802__PTR1), .ZN(_03854_) );
  AND2_X1 U17218 ( .A1(_03859_), .A2(_03884_), .ZN(_03855_) );
  AND2_X1 U17219 ( .A1(_03871_), .A2(_02802__PTR3), .ZN(_03856_) );
  AND2_X1 U17220 ( .A1(_03877_), .A2(_02802__PTR7), .ZN(_02802__PTR15) );
  AND2_X1 U17221 ( .A1(_02803__PTR3), .A2(_02803__PTR2), .ZN(_03857_) );
  AND2_X1 U17222 ( .A1(_02803__PTR5), .A2(_02803__PTR4), .ZN(_03858_) );
  AND2_X1 U17223 ( .A1(_02803__PTR7), .A2(_02803__PTR6), .ZN(_03859_) );
  AND2_X1 U17224 ( .A1(_02084__PTR41), .A2(_02084__PTR40), .ZN(_03860_) );
  AND2_X1 U17225 ( .A1(_02084__PTR43), .A2(_02084__PTR42), .ZN(_03861_) );
  AND2_X1 U17226 ( .A1(_02084__PTR45), .A2(_02084__PTR44), .ZN(_03862_) );
  AND2_X1 U17227 ( .A1(_02084__PTR47), .A2(_02084__PTR46), .ZN(_03863_) );
  AND2_X1 U17228 ( .A1(_02084__PTR49), .A2(_02084__PTR48), .ZN(_03864_) );
  AND2_X1 U17229 ( .A1(_02084__PTR51), .A2(_02084__PTR50), .ZN(_03865_) );
  AND2_X1 U17230 ( .A1(_02084__PTR53), .A2(_02084__PTR52), .ZN(_03866_) );
  AND2_X1 U17231 ( .A1(_02084__PTR55), .A2(_02084__PTR54), .ZN(_03867_) );
  AND2_X1 U17232 ( .A1(_02084__PTR57), .A2(_02084__PTR56), .ZN(_03868_) );
  AND2_X1 U17233 ( .A1(_02084__PTR59), .A2(_02084__PTR58), .ZN(_03869_) );
  AND2_X1 U17234 ( .A1(_02084__PTR61), .A2(_02084__PTR60), .ZN(_03870_) );
  AND2_X1 U17235 ( .A1(_03859_), .A2(_03858_), .ZN(_03871_) );
  AND2_X1 U17236 ( .A1(_03861_), .A2(_03860_), .ZN(_03872_) );
  AND2_X1 U17237 ( .A1(_03863_), .A2(_03862_), .ZN(_03873_) );
  AND2_X1 U17238 ( .A1(_03865_), .A2(_03864_), .ZN(_03874_) );
  AND2_X1 U17239 ( .A1(_03867_), .A2(_03866_), .ZN(_03875_) );
  AND2_X1 U17240 ( .A1(_03869_), .A2(_03868_), .ZN(_03876_) );
  AND2_X1 U17241 ( .A1(_03873_), .A2(_03872_), .ZN(_03877_) );
  AND2_X1 U17242 ( .A1(_03875_), .A2(_03874_), .ZN(_03878_) );
  AND2_X1 U17243 ( .A1(_03878_), .A2(_02802__PTR15), .ZN(_02802__PTR23) );
  AND2_X1 U17244 ( .A1(_03872_), .A2(_02802__PTR7), .ZN(_02802__PTR11) );
  AND2_X1 U17245 ( .A1(_03874_), .A2(_02802__PTR15), .ZN(_02802__PTR19) );
  AND2_X1 U17246 ( .A1(_03876_), .A2(_02802__PTR23), .ZN(_02802__PTR27) );
  AND2_X1 U17247 ( .A1(_03858_), .A2(_02802__PTR3), .ZN(_03879_) );
  AND2_X1 U17248 ( .A1(_03860_), .A2(_02802__PTR7), .ZN(_02802__PTR9) );
  AND2_X1 U17249 ( .A1(_03862_), .A2(_02802__PTR11), .ZN(_02802__PTR13) );
  AND2_X1 U17250 ( .A1(_03864_), .A2(_02802__PTR15), .ZN(_02802__PTR17) );
  AND2_X1 U17251 ( .A1(_03866_), .A2(_02802__PTR19), .ZN(_02802__PTR21) );
  AND2_X1 U17252 ( .A1(_03868_), .A2(_02802__PTR23), .ZN(_02802__PTR25) );
  AND2_X1 U17253 ( .A1(_03870_), .A2(_02802__PTR27), .ZN(_02802__PTR29) );
  AND2_X1 U17254 ( .A1(_02803__PTR2), .A2(_02802__PTR1), .ZN(_03880_) );
  AND2_X1 U17255 ( .A1(_02803__PTR4), .A2(_02802__PTR3), .ZN(_03881_) );
  AND2_X1 U17256 ( .A1(_02803__PTR6), .A2(_02802__PTR5), .ZN(_03882_) );
  AND2_X1 U17257 ( .A1(_02084__PTR40), .A2(_02802__PTR7), .ZN(_02802__PTR8) );
  AND2_X1 U17258 ( .A1(_02084__PTR42), .A2(_02802__PTR9), .ZN(_02802__PTR10) );
  AND2_X1 U17259 ( .A1(_02084__PTR44), .A2(_02802__PTR11), .ZN(_02802__PTR12) );
  AND2_X1 U17260 ( .A1(_02084__PTR46), .A2(_02802__PTR13), .ZN(_02802__PTR14) );
  AND2_X1 U17261 ( .A1(_02084__PTR48), .A2(_02802__PTR15), .ZN(_02802__PTR16) );
  AND2_X1 U17262 ( .A1(_02084__PTR50), .A2(_02802__PTR17), .ZN(_02802__PTR18) );
  AND2_X1 U17263 ( .A1(_02084__PTR52), .A2(_02802__PTR19), .ZN(_02802__PTR20) );
  AND2_X1 U17264 ( .A1(_02084__PTR54), .A2(_02802__PTR21), .ZN(_02802__PTR22) );
  AND2_X1 U17265 ( .A1(_02084__PTR56), .A2(_02802__PTR23), .ZN(_02802__PTR24) );
  AND2_X1 U17266 ( .A1(_02084__PTR58), .A2(_02802__PTR25), .ZN(_02802__PTR26) );
  AND2_X1 U17267 ( .A1(_02084__PTR60), .A2(_02802__PTR27), .ZN(_02802__PTR28) );
  AND2_X1 U17268 ( .A1(_02084__PTR62), .A2(_02802__PTR29), .ZN(_02802__PTR30) );
  OR2_X1 U17269 ( .A1(_02805__PTR1), .A2(_03850_), .ZN(_02802__PTR1) );
  OR2_X1 U17270 ( .A1(_02805__PTR3), .A2(_03851_), .ZN(_03883_) );
  OR2_X1 U17271 ( .A1(_02805__PTR5), .A2(_03852_), .ZN(_03884_) );
  OR2_X1 U17272 ( .A1(_02805__PTR7), .A2(_03853_), .ZN(_03885_) );
  OR2_X1 U17273 ( .A1(_03883_), .A2(_03854_), .ZN(_02802__PTR3) );
  OR2_X1 U17274 ( .A1(_03885_), .A2(_03855_), .ZN(_03886_) );
  OR2_X1 U17275 ( .A1(_03886_), .A2(_03856_), .ZN(_02802__PTR7) );
  OR2_X1 U17276 ( .A1(_03884_), .A2(_03879_), .ZN(_02802__PTR5) );
  OR2_X1 U17277 ( .A1(_02805__PTR2), .A2(_03880_), .ZN(_02802__PTR2) );
  OR2_X1 U17278 ( .A1(_02805__PTR4), .A2(_03881_), .ZN(_02802__PTR4) );
  OR2_X1 U17279 ( .A1(_02805__PTR6), .A2(_03882_), .ZN(_02802__PTR6) );
  AND2_X1 U17280 ( .A1(_01885__PTR7), .A2(_02723__PTR6), .ZN(_03984_) );
  AND2_X1 U17281 ( .A1(_03987_), .A2(_03534_), .ZN(_03985_) );
  AND2_X1 U17282 ( .A1(_03988_), .A2(_02724__PTR3), .ZN(_03986_) );
  AND2_X1 U17283 ( .A1(_01885__PTR7), .A2(_01885__PTR6), .ZN(_03987_) );
  AND2_X1 U17284 ( .A1(_03987_), .A2(_03527_), .ZN(_03988_) );
  OR2_X1 U17285 ( .A1(_02723__PTR7), .A2(_03984_), .ZN(_03989_) );
  OR2_X1 U17286 ( .A1(_03989_), .A2(_03985_), .ZN(_03990_) );
  OR2_X1 U17287 ( .A1(_03990_), .A2(_03986_), .ZN(_02934__PTR8) );
  AND2_X1 U17288 ( .A1(P1_P1_InstAddrPointer_PTR1), .A2(P1_P1_InstAddrPointer_PTR0), .ZN(_02798__PTR1) );
  AND2_X1 U17289 ( .A1(_03806_), .A2(_02798__PTR1), .ZN(_02798__PTR3) );
  AND2_X1 U17290 ( .A1(_03820_), .A2(_02798__PTR3), .ZN(_02798__PTR7) );
  AND2_X1 U17291 ( .A1(_03826_), .A2(_02798__PTR7), .ZN(_02798__PTR15) );
  AND2_X1 U17292 ( .A1(P1_P1_InstAddrPointer_PTR3), .A2(P1_P1_InstAddrPointer_PTR2), .ZN(_03806_) );
  AND2_X1 U17293 ( .A1(P1_P1_InstAddrPointer_PTR5), .A2(P1_P1_InstAddrPointer_PTR4), .ZN(_03807_) );
  AND2_X1 U17294 ( .A1(P1_P1_InstAddrPointer_PTR7), .A2(P1_P1_InstAddrPointer_PTR6), .ZN(_03808_) );
  AND2_X1 U17295 ( .A1(P1_P1_InstAddrPointer_PTR9), .A2(P1_P1_InstAddrPointer_PTR8), .ZN(_03809_) );
  AND2_X1 U17296 ( .A1(P1_P1_InstAddrPointer_PTR11), .A2(P1_P1_InstAddrPointer_PTR10), .ZN(_03810_) );
  AND2_X1 U17297 ( .A1(P1_P1_InstAddrPointer_PTR13), .A2(P1_P1_InstAddrPointer_PTR12), .ZN(_03811_) );
  AND2_X1 U17298 ( .A1(P1_P1_InstAddrPointer_PTR15), .A2(P1_P1_InstAddrPointer_PTR14), .ZN(_03812_) );
  AND2_X1 U17299 ( .A1(P1_P1_InstAddrPointer_PTR17), .A2(P1_P1_InstAddrPointer_PTR16), .ZN(_03813_) );
  AND2_X1 U17300 ( .A1(P1_P1_InstAddrPointer_PTR19), .A2(P1_P1_InstAddrPointer_PTR18), .ZN(_03814_) );
  AND2_X1 U17301 ( .A1(P1_P1_InstAddrPointer_PTR21), .A2(P1_P1_InstAddrPointer_PTR20), .ZN(_03815_) );
  AND2_X1 U17302 ( .A1(P1_P1_InstAddrPointer_PTR23), .A2(P1_P1_InstAddrPointer_PTR22), .ZN(_03816_) );
  AND2_X1 U17303 ( .A1(P1_P1_InstAddrPointer_PTR25), .A2(P1_P1_InstAddrPointer_PTR24), .ZN(_03817_) );
  AND2_X1 U17304 ( .A1(P1_P1_InstAddrPointer_PTR27), .A2(P1_P1_InstAddrPointer_PTR26), .ZN(_03818_) );
  AND2_X1 U17305 ( .A1(P1_P1_InstAddrPointer_PTR29), .A2(P1_P1_InstAddrPointer_PTR28), .ZN(_03819_) );
  AND2_X1 U17306 ( .A1(_03827_), .A2(_02798__PTR15), .ZN(_02798__PTR23) );
  AND2_X1 U17307 ( .A1(_03821_), .A2(_02798__PTR7), .ZN(_02798__PTR11) );
  AND2_X1 U17308 ( .A1(_03823_), .A2(_02798__PTR15), .ZN(_02798__PTR19) );
  AND2_X1 U17309 ( .A1(_03825_), .A2(_02798__PTR23), .ZN(_02798__PTR27) );
  AND2_X1 U17310 ( .A1(_03807_), .A2(_02798__PTR3), .ZN(_02798__PTR5) );
  AND2_X1 U17311 ( .A1(_03809_), .A2(_02798__PTR7), .ZN(_02798__PTR9) );
  AND2_X1 U17312 ( .A1(_03811_), .A2(_02798__PTR11), .ZN(_02798__PTR13) );
  AND2_X1 U17313 ( .A1(_03813_), .A2(_02798__PTR15), .ZN(_02798__PTR17) );
  AND2_X1 U17314 ( .A1(_03815_), .A2(_02798__PTR19), .ZN(_02798__PTR21) );
  AND2_X1 U17315 ( .A1(_03817_), .A2(_02798__PTR23), .ZN(_02798__PTR25) );
  AND2_X1 U17316 ( .A1(_03819_), .A2(_02798__PTR27), .ZN(_02798__PTR29) );
  AND2_X1 U17317 ( .A1(P1_P1_InstAddrPointer_PTR2), .A2(_02798__PTR1), .ZN(_02798__PTR2) );
  AND2_X1 U17318 ( .A1(P1_P1_InstAddrPointer_PTR4), .A2(_02798__PTR3), .ZN(_02798__PTR4) );
  AND2_X1 U17319 ( .A1(P1_P1_InstAddrPointer_PTR6), .A2(_02798__PTR5), .ZN(_02798__PTR6) );
  AND2_X1 U17320 ( .A1(P1_P1_InstAddrPointer_PTR8), .A2(_02798__PTR7), .ZN(_02798__PTR8) );
  AND2_X1 U17321 ( .A1(P1_P1_InstAddrPointer_PTR10), .A2(_02798__PTR9), .ZN(_02798__PTR10) );
  AND2_X1 U17322 ( .A1(P1_P1_InstAddrPointer_PTR12), .A2(_02798__PTR11), .ZN(_02798__PTR12) );
  AND2_X1 U17323 ( .A1(P1_P1_InstAddrPointer_PTR14), .A2(_02798__PTR13), .ZN(_02798__PTR14) );
  AND2_X1 U17324 ( .A1(P1_P1_InstAddrPointer_PTR16), .A2(_02798__PTR15), .ZN(_02798__PTR16) );
  AND2_X1 U17325 ( .A1(P1_P1_InstAddrPointer_PTR18), .A2(_02798__PTR17), .ZN(_02798__PTR18) );
  AND2_X1 U17326 ( .A1(P1_P1_InstAddrPointer_PTR20), .A2(_02798__PTR19), .ZN(_02798__PTR20) );
  AND2_X1 U17327 ( .A1(P1_P1_InstAddrPointer_PTR22), .A2(_02798__PTR21), .ZN(_02798__PTR22) );
  AND2_X1 U17328 ( .A1(P1_P1_InstAddrPointer_PTR24), .A2(_02798__PTR23), .ZN(_02798__PTR24) );
  AND2_X1 U17329 ( .A1(P1_P1_InstAddrPointer_PTR26), .A2(_02798__PTR25), .ZN(_02798__PTR26) );
  AND2_X1 U17330 ( .A1(P1_P1_InstAddrPointer_PTR28), .A2(_02798__PTR27), .ZN(_02798__PTR28) );
  AND2_X1 U17331 ( .A1(P1_P1_InstAddrPointer_PTR30), .A2(_02798__PTR29), .ZN(_02798__PTR30) );
  AND2_X1 U17332 ( .A1(_02809__PTR1), .A2(_02937__PTR0), .ZN(_03991_) );
  AND2_X1 U17333 ( .A1(_02938__PTR3), .A2(_02940__PTR2), .ZN(_03992_) );
  AND2_X1 U17334 ( .A1(_02938__PTR5), .A2(_02940__PTR4), .ZN(_03993_) );
  AND2_X1 U17335 ( .A1(_02938__PTR7), .A2(_02940__PTR6), .ZN(_03994_) );
  AND2_X1 U17336 ( .A1(_02938__PTR9), .A2(_02940__PTR8), .ZN(_03995_) );
  AND2_X1 U17337 ( .A1(_02938__PTR11), .A2(_02940__PTR10), .ZN(_03996_) );
  AND2_X1 U17338 ( .A1(_02938__PTR13), .A2(_02940__PTR12), .ZN(_03997_) );
  AND2_X1 U17339 ( .A1(_02938__PTR15), .A2(_02940__PTR14), .ZN(_03998_) );
  AND2_X1 U17340 ( .A1(_02938__PTR17), .A2(_02940__PTR16), .ZN(_03999_) );
  AND2_X1 U17341 ( .A1(_02938__PTR19), .A2(_02940__PTR18), .ZN(_04000_) );
  AND2_X1 U17342 ( .A1(_02938__PTR21), .A2(_02940__PTR20), .ZN(_04001_) );
  AND2_X1 U17343 ( .A1(_02938__PTR23), .A2(_02940__PTR22), .ZN(_04002_) );
  AND2_X1 U17344 ( .A1(_02938__PTR25), .A2(_02940__PTR24), .ZN(_04003_) );
  AND2_X1 U17345 ( .A1(_02938__PTR27), .A2(_02940__PTR26), .ZN(_04004_) );
  AND2_X1 U17346 ( .A1(_02938__PTR29), .A2(_02940__PTR28), .ZN(_04005_) );
  AND2_X1 U17347 ( .A1(_04017_), .A2(_02937__PTR1), .ZN(_04006_) );
  AND2_X1 U17348 ( .A1(_04019_), .A2(_04066_), .ZN(_04007_) );
  AND2_X1 U17349 ( .A1(_04021_), .A2(_04068_), .ZN(_04008_) );
  AND2_X1 U17350 ( .A1(_04023_), .A2(_04070_), .ZN(_04009_) );
  AND2_X1 U17351 ( .A1(_04025_), .A2(_04072_), .ZN(_04010_) );
  AND2_X1 U17352 ( .A1(_04027_), .A2(_04074_), .ZN(_04011_) );
  AND2_X1 U17353 ( .A1(_04029_), .A2(_04076_), .ZN(_04012_) );
  AND2_X1 U17354 ( .A1(_04031_), .A2(_02937__PTR3), .ZN(_04013_) );
  AND2_X1 U17355 ( .A1(_04033_), .A2(_04080_), .ZN(_04014_) );
  AND2_X1 U17356 ( .A1(_04035_), .A2(_04082_), .ZN(_04015_) );
  AND2_X1 U17357 ( .A1(_04037_), .A2(_02937__PTR7), .ZN(_04016_) );
  AND2_X1 U17358 ( .A1(_02938__PTR3), .A2(_02938__PTR2), .ZN(_04017_) );
  AND2_X1 U17359 ( .A1(_02938__PTR5), .A2(_02938__PTR4), .ZN(_04018_) );
  AND2_X1 U17360 ( .A1(_02938__PTR7), .A2(_02938__PTR6), .ZN(_04019_) );
  AND2_X1 U17361 ( .A1(_02938__PTR9), .A2(_02938__PTR8), .ZN(_04020_) );
  AND2_X1 U17362 ( .A1(_02938__PTR11), .A2(_02938__PTR10), .ZN(_04021_) );
  AND2_X1 U17363 ( .A1(_02938__PTR13), .A2(_02938__PTR12), .ZN(_04022_) );
  AND2_X1 U17364 ( .A1(_02938__PTR15), .A2(_02938__PTR14), .ZN(_04023_) );
  AND2_X1 U17365 ( .A1(_02938__PTR17), .A2(_02938__PTR16), .ZN(_04024_) );
  AND2_X1 U17366 ( .A1(_02938__PTR19), .A2(_02938__PTR18), .ZN(_04025_) );
  AND2_X1 U17367 ( .A1(_02938__PTR21), .A2(_02938__PTR20), .ZN(_04026_) );
  AND2_X1 U17368 ( .A1(_02938__PTR23), .A2(_02938__PTR22), .ZN(_04027_) );
  AND2_X1 U17369 ( .A1(_02938__PTR25), .A2(_02938__PTR24), .ZN(_04028_) );
  AND2_X1 U17370 ( .A1(_02938__PTR27), .A2(_02938__PTR26), .ZN(_04029_) );
  AND2_X1 U17371 ( .A1(_02938__PTR29), .A2(_02938__PTR28), .ZN(_04030_) );
  AND2_X1 U17372 ( .A1(_04019_), .A2(_04018_), .ZN(_04031_) );
  AND2_X1 U17373 ( .A1(_04021_), .A2(_04020_), .ZN(_04032_) );
  AND2_X1 U17374 ( .A1(_04023_), .A2(_04022_), .ZN(_04033_) );
  AND2_X1 U17375 ( .A1(_04025_), .A2(_04024_), .ZN(_04034_) );
  AND2_X1 U17376 ( .A1(_04027_), .A2(_04026_), .ZN(_04035_) );
  AND2_X1 U17377 ( .A1(_04029_), .A2(_04028_), .ZN(_04036_) );
  AND2_X1 U17378 ( .A1(_04033_), .A2(_04032_), .ZN(_04037_) );
  AND2_X1 U17379 ( .A1(_04035_), .A2(_04034_), .ZN(_04038_) );
  AND2_X1 U17380 ( .A1(_04038_), .A2(_02937__PTR15), .ZN(_04039_) );
  AND2_X1 U17381 ( .A1(_04032_), .A2(_02937__PTR7), .ZN(_04040_) );
  AND2_X1 U17382 ( .A1(_04034_), .A2(_02937__PTR15), .ZN(_04041_) );
  AND2_X1 U17383 ( .A1(_04036_), .A2(_02937__PTR23), .ZN(_04042_) );
  AND2_X1 U17384 ( .A1(_04018_), .A2(_02937__PTR3), .ZN(_04043_) );
  AND2_X1 U17385 ( .A1(_04020_), .A2(_02937__PTR7), .ZN(_04044_) );
  AND2_X1 U17386 ( .A1(_04022_), .A2(_02937__PTR11), .ZN(_04045_) );
  AND2_X1 U17387 ( .A1(_04024_), .A2(_02937__PTR15), .ZN(_04046_) );
  AND2_X1 U17388 ( .A1(_04026_), .A2(_02937__PTR19), .ZN(_04047_) );
  AND2_X1 U17389 ( .A1(_04028_), .A2(_02937__PTR23), .ZN(_04048_) );
  AND2_X1 U17390 ( .A1(_04030_), .A2(_02937__PTR27), .ZN(_04049_) );
  AND2_X1 U17391 ( .A1(_02938__PTR2), .A2(_02937__PTR1), .ZN(_04050_) );
  AND2_X1 U17392 ( .A1(_02938__PTR4), .A2(_02937__PTR3), .ZN(_04051_) );
  AND2_X1 U17393 ( .A1(_02938__PTR6), .A2(_02937__PTR5), .ZN(_04052_) );
  AND2_X1 U17394 ( .A1(_02938__PTR8), .A2(_02937__PTR7), .ZN(_04053_) );
  AND2_X1 U17395 ( .A1(_02938__PTR10), .A2(_02937__PTR9), .ZN(_04054_) );
  AND2_X1 U17396 ( .A1(_02938__PTR12), .A2(_02937__PTR11), .ZN(_04055_) );
  AND2_X1 U17397 ( .A1(_02938__PTR14), .A2(_02937__PTR13), .ZN(_04056_) );
  AND2_X1 U17398 ( .A1(_02938__PTR16), .A2(_02937__PTR15), .ZN(_04057_) );
  AND2_X1 U17399 ( .A1(_02938__PTR18), .A2(_02937__PTR17), .ZN(_04058_) );
  AND2_X1 U17400 ( .A1(_02938__PTR20), .A2(_02937__PTR19), .ZN(_04059_) );
  AND2_X1 U17401 ( .A1(_02938__PTR22), .A2(_02937__PTR21), .ZN(_04060_) );
  AND2_X1 U17402 ( .A1(_02938__PTR24), .A2(_02937__PTR23), .ZN(_04061_) );
  AND2_X1 U17403 ( .A1(_02938__PTR26), .A2(_02937__PTR25), .ZN(_04062_) );
  AND2_X1 U17404 ( .A1(_02938__PTR28), .A2(_02937__PTR27), .ZN(_04063_) );
  AND2_X1 U17405 ( .A1(_02938__PTR30), .A2(_02937__PTR29), .ZN(_04064_) );
  OR2_X1 U17406 ( .A1(_02808__PTR0), .A2(_02809__PTR0), .ZN(_02937__PTR0) );
  OR2_X1 U17407 ( .A1(_02811__PTR1), .A2(_03991_), .ZN(_02937__PTR1) );
  OR2_X1 U17408 ( .A1(_02940__PTR3), .A2(_03992_), .ZN(_04065_) );
  OR2_X1 U17409 ( .A1(_02940__PTR5), .A2(_03993_), .ZN(_04066_) );
  OR2_X1 U17410 ( .A1(_02940__PTR7), .A2(_03994_), .ZN(_04067_) );
  OR2_X1 U17411 ( .A1(_02940__PTR9), .A2(_03995_), .ZN(_04068_) );
  OR2_X1 U17412 ( .A1(_02940__PTR11), .A2(_03996_), .ZN(_04069_) );
  OR2_X1 U17413 ( .A1(_02940__PTR13), .A2(_03997_), .ZN(_04070_) );
  OR2_X1 U17414 ( .A1(_02940__PTR15), .A2(_03998_), .ZN(_04071_) );
  OR2_X1 U17415 ( .A1(_02940__PTR17), .A2(_03999_), .ZN(_04072_) );
  OR2_X1 U17416 ( .A1(_02940__PTR19), .A2(_04000_), .ZN(_04073_) );
  OR2_X1 U17417 ( .A1(_02940__PTR21), .A2(_04001_), .ZN(_04074_) );
  OR2_X1 U17418 ( .A1(_02940__PTR23), .A2(_04002_), .ZN(_04075_) );
  OR2_X1 U17419 ( .A1(_02940__PTR25), .A2(_04003_), .ZN(_04076_) );
  OR2_X1 U17420 ( .A1(_02940__PTR27), .A2(_04004_), .ZN(_04077_) );
  OR2_X1 U17421 ( .A1(_02940__PTR29), .A2(_04005_), .ZN(_04078_) );
  OR2_X1 U17422 ( .A1(_04065_), .A2(_04006_), .ZN(_02937__PTR3) );
  OR2_X1 U17423 ( .A1(_04067_), .A2(_04007_), .ZN(_04079_) );
  OR2_X1 U17424 ( .A1(_04069_), .A2(_04008_), .ZN(_04080_) );
  OR2_X1 U17425 ( .A1(_04071_), .A2(_04009_), .ZN(_04081_) );
  OR2_X1 U17426 ( .A1(_04073_), .A2(_04010_), .ZN(_04082_) );
  OR2_X1 U17427 ( .A1(_04075_), .A2(_04011_), .ZN(_04083_) );
  OR2_X1 U17428 ( .A1(_04077_), .A2(_04012_), .ZN(_04084_) );
  OR2_X1 U17429 ( .A1(_04079_), .A2(_04013_), .ZN(_02937__PTR7) );
  OR2_X1 U17430 ( .A1(_04081_), .A2(_04014_), .ZN(_04085_) );
  OR2_X1 U17431 ( .A1(_04083_), .A2(_04015_), .ZN(_04086_) );
  OR2_X1 U17432 ( .A1(_04085_), .A2(_04016_), .ZN(_02937__PTR15) );
  OR2_X1 U17433 ( .A1(_04086_), .A2(_04039_), .ZN(_02937__PTR23) );
  OR2_X1 U17434 ( .A1(_04080_), .A2(_04040_), .ZN(_02937__PTR11) );
  OR2_X1 U17435 ( .A1(_04082_), .A2(_04041_), .ZN(_02937__PTR19) );
  OR2_X1 U17436 ( .A1(_04084_), .A2(_04042_), .ZN(_02937__PTR27) );
  OR2_X1 U17437 ( .A1(_04066_), .A2(_04043_), .ZN(_02937__PTR5) );
  OR2_X1 U17438 ( .A1(_04068_), .A2(_04044_), .ZN(_02937__PTR9) );
  OR2_X1 U17439 ( .A1(_04070_), .A2(_04045_), .ZN(_02937__PTR13) );
  OR2_X1 U17440 ( .A1(_04072_), .A2(_04046_), .ZN(_02937__PTR17) );
  OR2_X1 U17441 ( .A1(_04074_), .A2(_04047_), .ZN(_02937__PTR21) );
  OR2_X1 U17442 ( .A1(_04076_), .A2(_04048_), .ZN(_02937__PTR25) );
  OR2_X1 U17443 ( .A1(_04078_), .A2(_04049_), .ZN(_02937__PTR29) );
  OR2_X1 U17444 ( .A1(_02940__PTR2), .A2(_04050_), .ZN(_02937__PTR2) );
  OR2_X1 U17445 ( .A1(_02940__PTR4), .A2(_04051_), .ZN(_02937__PTR4) );
  OR2_X1 U17446 ( .A1(_02940__PTR6), .A2(_04052_), .ZN(_02937__PTR6) );
  OR2_X1 U17447 ( .A1(_02940__PTR8), .A2(_04053_), .ZN(_02937__PTR8) );
  OR2_X1 U17448 ( .A1(_02940__PTR10), .A2(_04054_), .ZN(_02937__PTR10) );
  OR2_X1 U17449 ( .A1(_02940__PTR12), .A2(_04055_), .ZN(_02937__PTR12) );
  OR2_X1 U17450 ( .A1(_02940__PTR14), .A2(_04056_), .ZN(_02937__PTR14) );
  OR2_X1 U17451 ( .A1(_02940__PTR16), .A2(_04057_), .ZN(_02937__PTR16) );
  OR2_X1 U17452 ( .A1(_02940__PTR18), .A2(_04058_), .ZN(_02937__PTR18) );
  OR2_X1 U17453 ( .A1(_02940__PTR20), .A2(_04059_), .ZN(_02937__PTR20) );
  OR2_X1 U17454 ( .A1(_02940__PTR22), .A2(_04060_), .ZN(_02937__PTR22) );
  OR2_X1 U17455 ( .A1(_02940__PTR24), .A2(_04061_), .ZN(_02937__PTR24) );
  OR2_X1 U17456 ( .A1(_02940__PTR26), .A2(_04062_), .ZN(_02937__PTR26) );
  OR2_X1 U17457 ( .A1(_02940__PTR28), .A2(_04063_), .ZN(_02937__PTR28) );
  OR2_X1 U17458 ( .A1(_02940__PTR30), .A2(_04064_), .ZN(_02937__PTR30) );
  AND2_X1 U17459 ( .A1(_01885__PTR3), .A2(_02723__PTR2), .ZN(_03521_) );
  AND2_X1 U17460 ( .A1(_01885__PTR5), .A2(_02723__PTR4), .ZN(_03522_) );
  AND2_X1 U17461 ( .A1(_02723__PTR7), .A2(_02723__PTR6), .ZN(_03523_) );
  AND2_X1 U17462 ( .A1(_03528_), .A2(_03534_), .ZN(_03525_) );
  AND2_X1 U17463 ( .A1(_03529_), .A2(_02724__PTR3), .ZN(_03526_) );
  AND2_X1 U17464 ( .A1(_01885__PTR3), .A2(_01885__PTR2), .ZN(_03524_) );
  AND2_X1 U17465 ( .A1(_01885__PTR5), .A2(_01885__PTR4), .ZN(_03527_) );
  AND2_X1 U17466 ( .A1(_02723__PTR7), .A2(_01885__PTR6), .ZN(_03528_) );
  AND2_X1 U17467 ( .A1(_03528_), .A2(_03527_), .ZN(_03529_) );
  AND2_X1 U17468 ( .A1(_03527_), .A2(_02724__PTR3), .ZN(_03530_) );
  AND2_X1 U17469 ( .A1(_01885__PTR4), .A2(_02724__PTR3), .ZN(_03531_) );
  AND2_X1 U17470 ( .A1(_01885__PTR6), .A2(_02724__PTR5), .ZN(_03532_) );
  OR2_X1 U17471 ( .A1(_02723__PTR3), .A2(_03521_), .ZN(_03533_) );
  OR2_X1 U17472 ( .A1(_02723__PTR5), .A2(_03522_), .ZN(_03534_) );
  OR2_X1 U17473 ( .A1(_03533_), .A2(_03524_), .ZN(_02724__PTR3) );
  OR2_X1 U17474 ( .A1(_03523_), .A2(_03525_), .ZN(_03535_) );
  OR2_X1 U17475 ( .A1(_03535_), .A2(_03526_), .ZN(_02724__PTR7) );
  OR2_X1 U17476 ( .A1(_03534_), .A2(_03530_), .ZN(_02724__PTR5) );
  OR2_X1 U17477 ( .A1(_02723__PTR4), .A2(_03531_), .ZN(_02724__PTR4) );
  OR2_X1 U17478 ( .A1(_02723__PTR6), .A2(_03532_), .ZN(_02724__PTR6) );
  AND2_X1 U17479 ( .A1(_02718__PTR3), .A2(_02718__PTR2), .ZN(_02719__PTR3) );
  AND2_X1 U17480 ( .A1(_00618__PTR2), .A2(_02719__PTR3), .ZN(_03520_) );
  OR2_X1 U17481 ( .A1(_02716__PTR5), .A2(_03520_), .ZN(_02719__PTR5) );
  AND2_X1 U17482 ( .A1(P1_P1_InstQueueRd_Addr_PTR1), .A2(P1_P1_InstQueueRd_Addr_PTR0), .ZN(_02750__PTR1) );
  AND2_X1 U17483 ( .A1(P1_P1_InstQueueRd_Addr_PTR3), .A2(P1_P1_InstQueueRd_Addr_PTR2), .ZN(_02812__PTR1) );
  AND2_X1 U17484 ( .A1(P1_P1_InstQueueRd_Addr_PTR4), .A2(_02750__PTR3), .ZN(_02799__PTR4) );
  AND2_X1 U17485 ( .A1(P1_P1_PhyAddrPointer_PTR2), .A2(P1_P1_PhyAddrPointer_PTR1), .ZN(_02797__PTR1) );
  AND2_X1 U17486 ( .A1(_03784_), .A2(_02797__PTR1), .ZN(_02797__PTR3) );
  AND2_X1 U17487 ( .A1(_03798_), .A2(_02797__PTR3), .ZN(_02797__PTR7) );
  AND2_X1 U17488 ( .A1(_03804_), .A2(_02797__PTR7), .ZN(_02797__PTR15) );
  AND2_X1 U17489 ( .A1(P1_P1_PhyAddrPointer_PTR4), .A2(P1_P1_PhyAddrPointer_PTR3), .ZN(_03784_) );
  AND2_X1 U17490 ( .A1(P1_P1_PhyAddrPointer_PTR6), .A2(P1_P1_PhyAddrPointer_PTR5), .ZN(_03785_) );
  AND2_X1 U17491 ( .A1(P1_P1_PhyAddrPointer_PTR8), .A2(P1_P1_PhyAddrPointer_PTR7), .ZN(_03786_) );
  AND2_X1 U17492 ( .A1(P1_P1_PhyAddrPointer_PTR10), .A2(P1_P1_PhyAddrPointer_PTR9), .ZN(_03787_) );
  AND2_X1 U17493 ( .A1(P1_P1_PhyAddrPointer_PTR12), .A2(P1_P1_PhyAddrPointer_PTR11), .ZN(_03788_) );
  AND2_X1 U17494 ( .A1(P1_P1_PhyAddrPointer_PTR14), .A2(P1_P1_PhyAddrPointer_PTR13), .ZN(_03789_) );
  AND2_X1 U17495 ( .A1(P1_P1_PhyAddrPointer_PTR16), .A2(P1_P1_PhyAddrPointer_PTR15), .ZN(_03790_) );
  AND2_X1 U17496 ( .A1(P1_P1_PhyAddrPointer_PTR18), .A2(P1_P1_PhyAddrPointer_PTR17), .ZN(_03791_) );
  AND2_X1 U17497 ( .A1(P1_P1_PhyAddrPointer_PTR20), .A2(P1_P1_PhyAddrPointer_PTR19), .ZN(_03792_) );
  AND2_X1 U17498 ( .A1(P1_P1_PhyAddrPointer_PTR22), .A2(P1_P1_PhyAddrPointer_PTR21), .ZN(_03793_) );
  AND2_X1 U17499 ( .A1(P1_P1_PhyAddrPointer_PTR24), .A2(P1_P1_PhyAddrPointer_PTR23), .ZN(_03794_) );
  AND2_X1 U17500 ( .A1(P1_P1_PhyAddrPointer_PTR26), .A2(P1_P1_PhyAddrPointer_PTR25), .ZN(_03795_) );
  AND2_X1 U17501 ( .A1(P1_P1_PhyAddrPointer_PTR28), .A2(P1_P1_PhyAddrPointer_PTR27), .ZN(_03796_) );
  AND2_X1 U17502 ( .A1(P1_P1_PhyAddrPointer_PTR30), .A2(P1_P1_PhyAddrPointer_PTR29), .ZN(_03797_) );
  AND2_X1 U17503 ( .A1(_03786_), .A2(_03785_), .ZN(_03798_) );
  AND2_X1 U17504 ( .A1(_03788_), .A2(_03787_), .ZN(_03799_) );
  AND2_X1 U17505 ( .A1(_03790_), .A2(_03789_), .ZN(_03800_) );
  AND2_X1 U17506 ( .A1(_03792_), .A2(_03791_), .ZN(_03801_) );
  AND2_X1 U17507 ( .A1(_03794_), .A2(_03793_), .ZN(_03802_) );
  AND2_X1 U17508 ( .A1(_03796_), .A2(_03795_), .ZN(_03803_) );
  AND2_X1 U17509 ( .A1(_03800_), .A2(_03799_), .ZN(_03804_) );
  AND2_X1 U17510 ( .A1(_03802_), .A2(_03801_), .ZN(_03805_) );
  AND2_X1 U17511 ( .A1(_03805_), .A2(_02797__PTR15), .ZN(_02797__PTR23) );
  AND2_X1 U17512 ( .A1(_03799_), .A2(_02797__PTR7), .ZN(_02797__PTR11) );
  AND2_X1 U17513 ( .A1(_03801_), .A2(_02797__PTR15), .ZN(_02797__PTR19) );
  AND2_X1 U17514 ( .A1(_03803_), .A2(_02797__PTR23), .ZN(_02797__PTR27) );
  AND2_X1 U17515 ( .A1(_03785_), .A2(_02797__PTR3), .ZN(_02797__PTR5) );
  AND2_X1 U17516 ( .A1(_03787_), .A2(_02797__PTR7), .ZN(_02797__PTR9) );
  AND2_X1 U17517 ( .A1(_03789_), .A2(_02797__PTR11), .ZN(_02797__PTR13) );
  AND2_X1 U17518 ( .A1(_03791_), .A2(_02797__PTR15), .ZN(_02797__PTR17) );
  AND2_X1 U17519 ( .A1(_03793_), .A2(_02797__PTR19), .ZN(_02797__PTR21) );
  AND2_X1 U17520 ( .A1(_03795_), .A2(_02797__PTR23), .ZN(_02797__PTR25) );
  AND2_X1 U17521 ( .A1(_03797_), .A2(_02797__PTR27), .ZN(_02797__PTR29) );
  AND2_X1 U17522 ( .A1(P1_P1_PhyAddrPointer_PTR3), .A2(_02797__PTR1), .ZN(_02797__PTR2) );
  AND2_X1 U17523 ( .A1(P1_P1_PhyAddrPointer_PTR5), .A2(_02797__PTR3), .ZN(_02797__PTR4) );
  AND2_X1 U17524 ( .A1(P1_P1_PhyAddrPointer_PTR7), .A2(_02797__PTR5), .ZN(_02797__PTR6) );
  AND2_X1 U17525 ( .A1(P1_P1_PhyAddrPointer_PTR9), .A2(_02797__PTR7), .ZN(_02797__PTR8) );
  AND2_X1 U17526 ( .A1(P1_P1_PhyAddrPointer_PTR11), .A2(_02797__PTR9), .ZN(_02797__PTR10) );
  AND2_X1 U17527 ( .A1(P1_P1_PhyAddrPointer_PTR13), .A2(_02797__PTR11), .ZN(_02797__PTR12) );
  AND2_X1 U17528 ( .A1(P1_P1_PhyAddrPointer_PTR15), .A2(_02797__PTR13), .ZN(_02797__PTR14) );
  AND2_X1 U17529 ( .A1(P1_P1_PhyAddrPointer_PTR17), .A2(_02797__PTR15), .ZN(_02797__PTR16) );
  AND2_X1 U17530 ( .A1(P1_P1_PhyAddrPointer_PTR19), .A2(_02797__PTR17), .ZN(_02797__PTR18) );
  AND2_X1 U17531 ( .A1(P1_P1_PhyAddrPointer_PTR21), .A2(_02797__PTR19), .ZN(_02797__PTR20) );
  AND2_X1 U17532 ( .A1(P1_P1_PhyAddrPointer_PTR23), .A2(_02797__PTR21), .ZN(_02797__PTR22) );
  AND2_X1 U17533 ( .A1(P1_P1_PhyAddrPointer_PTR25), .A2(_02797__PTR23), .ZN(_02797__PTR24) );
  AND2_X1 U17534 ( .A1(P1_P1_PhyAddrPointer_PTR27), .A2(_02797__PTR25), .ZN(_02797__PTR26) );
  AND2_X1 U17535 ( .A1(P1_P1_PhyAddrPointer_PTR29), .A2(_02797__PTR27), .ZN(_02797__PTR28) );
  AND2_X1 U17536 ( .A1(P1_P1_PhyAddrPointer_PTR1), .A2(_02715__PTR0), .ZN(_02945__PTR1) );
  AND2_X1 U17537 ( .A1(_03455_), .A2(_02945__PTR1), .ZN(_02945__PTR3) );
  AND2_X1 U17538 ( .A1(_03484_), .A2(_02945__PTR3), .ZN(_02945__PTR7) );
  AND2_X1 U17539 ( .A1(_03491_), .A2(_02945__PTR7), .ZN(_02945__PTR15) );
  AND2_X1 U17540 ( .A1(_03492_), .A2(_02945__PTR15), .ZN(_02945__PTR23) );
  AND2_X1 U17541 ( .A1(_03485_), .A2(_02945__PTR7), .ZN(_02945__PTR11) );
  AND2_X1 U17542 ( .A1(_03487_), .A2(_02945__PTR15), .ZN(_02945__PTR19) );
  AND2_X1 U17543 ( .A1(_03489_), .A2(_02945__PTR23), .ZN(_02945__PTR27) );
  AND2_X1 U17544 ( .A1(_03470_), .A2(_02945__PTR3), .ZN(_02945__PTR5) );
  AND2_X1 U17545 ( .A1(_03472_), .A2(_02945__PTR7), .ZN(_02945__PTR9) );
  AND2_X1 U17546 ( .A1(_03474_), .A2(_02945__PTR11), .ZN(_02945__PTR13) );
  AND2_X1 U17547 ( .A1(_03476_), .A2(_02945__PTR15), .ZN(_02945__PTR17) );
  AND2_X1 U17548 ( .A1(_03478_), .A2(_02945__PTR19), .ZN(_02945__PTR21) );
  AND2_X1 U17549 ( .A1(_03480_), .A2(_02945__PTR23), .ZN(_02945__PTR25) );
  AND2_X1 U17550 ( .A1(_03482_), .A2(_02945__PTR27), .ZN(_02945__PTR29) );
  AND2_X1 U17551 ( .A1(_02715__PTR2), .A2(_02945__PTR1), .ZN(_02945__PTR2) );
  AND2_X1 U17552 ( .A1(_02715__PTR4), .A2(_02945__PTR3), .ZN(_02945__PTR4) );
  AND2_X1 U17553 ( .A1(_02715__PTR6), .A2(_02945__PTR5), .ZN(_02945__PTR6) );
  AND2_X1 U17554 ( .A1(_02715__PTR8), .A2(_02945__PTR7), .ZN(_02945__PTR8) );
  AND2_X1 U17555 ( .A1(_02715__PTR10), .A2(_02945__PTR9), .ZN(_02945__PTR10) );
  AND2_X1 U17556 ( .A1(_02715__PTR12), .A2(_02945__PTR11), .ZN(_02945__PTR12) );
  AND2_X1 U17557 ( .A1(_02715__PTR14), .A2(_02945__PTR13), .ZN(_02945__PTR14) );
  AND2_X1 U17558 ( .A1(_02715__PTR16), .A2(_02945__PTR15), .ZN(_02945__PTR16) );
  AND2_X1 U17559 ( .A1(_02715__PTR18), .A2(_02945__PTR17), .ZN(_02945__PTR18) );
  AND2_X1 U17560 ( .A1(_02715__PTR20), .A2(_02945__PTR19), .ZN(_02945__PTR20) );
  AND2_X1 U17561 ( .A1(_02715__PTR22), .A2(_02945__PTR21), .ZN(_02945__PTR22) );
  AND2_X1 U17562 ( .A1(_02715__PTR24), .A2(_02945__PTR23), .ZN(_02945__PTR24) );
  AND2_X1 U17563 ( .A1(_02715__PTR26), .A2(_02945__PTR25), .ZN(_02945__PTR26) );
  AND2_X1 U17564 ( .A1(_02715__PTR28), .A2(_02945__PTR27), .ZN(_02945__PTR28) );
  AND2_X1 U17565 ( .A1(_02715__PTR30), .A2(_02945__PTR29), .ZN(_02945__PTR30) );
  AND2_X1 U17566 ( .A1(_02715__PTR3), .A2(_01892__PTR130), .ZN(_03440_) );
  AND2_X1 U17567 ( .A1(_02715__PTR5), .A2(_01892__PTR132), .ZN(_03441_) );
  AND2_X1 U17568 ( .A1(_02715__PTR7), .A2(_01892__PTR134), .ZN(_03442_) );
  AND2_X1 U17569 ( .A1(_02715__PTR9), .A2(_01892__PTR136), .ZN(_03443_) );
  AND2_X1 U17570 ( .A1(_02715__PTR11), .A2(_01892__PTR138), .ZN(_03444_) );
  AND2_X1 U17571 ( .A1(_02715__PTR13), .A2(_01892__PTR140), .ZN(_03445_) );
  AND2_X1 U17572 ( .A1(_02715__PTR15), .A2(_01892__PTR142), .ZN(_03446_) );
  AND2_X1 U17573 ( .A1(_02715__PTR17), .A2(_01892__PTR144), .ZN(_03447_) );
  AND2_X1 U17574 ( .A1(_02715__PTR19), .A2(_01892__PTR146), .ZN(_03448_) );
  AND2_X1 U17575 ( .A1(_02715__PTR21), .A2(_01892__PTR148), .ZN(_03449_) );
  AND2_X1 U17576 ( .A1(_02715__PTR23), .A2(_01892__PTR150), .ZN(_03450_) );
  AND2_X1 U17577 ( .A1(_02715__PTR25), .A2(_01892__PTR152), .ZN(_03451_) );
  AND2_X1 U17578 ( .A1(_02715__PTR27), .A2(_01892__PTR154), .ZN(_03452_) );
  AND2_X1 U17579 ( .A1(_02715__PTR29), .A2(_01892__PTR156), .ZN(_03453_) );
  AND2_X1 U17580 ( .A1(_02713__PTR31), .A2(_01892__PTR158), .ZN(_03454_) );
  AND2_X1 U17581 ( .A1(_03471_), .A2(_03496_), .ZN(_03456_) );
  AND2_X1 U17582 ( .A1(_03473_), .A2(_03498_), .ZN(_03457_) );
  AND2_X1 U17583 ( .A1(_03475_), .A2(_03500_), .ZN(_03458_) );
  AND2_X1 U17584 ( .A1(_03477_), .A2(_03502_), .ZN(_03459_) );
  AND2_X1 U17585 ( .A1(_03479_), .A2(_03504_), .ZN(_03460_) );
  AND2_X1 U17586 ( .A1(_03481_), .A2(_03506_), .ZN(_03461_) );
  AND2_X1 U17587 ( .A1(_03483_), .A2(_03508_), .ZN(_03462_) );
  AND2_X1 U17588 ( .A1(_03484_), .A2(_02714__PTR3), .ZN(_03463_) );
  AND2_X1 U17589 ( .A1(_03486_), .A2(_03510_), .ZN(_03464_) );
  AND2_X1 U17590 ( .A1(_03488_), .A2(_03512_), .ZN(_03465_) );
  AND2_X1 U17591 ( .A1(_03490_), .A2(_03514_), .ZN(_03466_) );
  AND2_X1 U17592 ( .A1(_03491_), .A2(_02714__PTR7), .ZN(_03467_) );
  AND2_X1 U17593 ( .A1(_03493_), .A2(_03517_), .ZN(_03468_) );
  AND2_X1 U17594 ( .A1(_03494_), .A2(_02714__PTR15), .ZN(_03469_) );
  AND2_X1 U17595 ( .A1(_02715__PTR3), .A2(_02715__PTR2), .ZN(_03455_) );
  AND2_X1 U17596 ( .A1(_02715__PTR5), .A2(_02715__PTR4), .ZN(_03470_) );
  AND2_X1 U17597 ( .A1(_02715__PTR7), .A2(_02715__PTR6), .ZN(_03471_) );
  AND2_X1 U17598 ( .A1(_02715__PTR9), .A2(_02715__PTR8), .ZN(_03472_) );
  AND2_X1 U17599 ( .A1(_02715__PTR11), .A2(_02715__PTR10), .ZN(_03473_) );
  AND2_X1 U17600 ( .A1(_02715__PTR13), .A2(_02715__PTR12), .ZN(_03474_) );
  AND2_X1 U17601 ( .A1(_02715__PTR15), .A2(_02715__PTR14), .ZN(_03475_) );
  AND2_X1 U17602 ( .A1(_02715__PTR17), .A2(_02715__PTR16), .ZN(_03476_) );
  AND2_X1 U17603 ( .A1(_02715__PTR19), .A2(_02715__PTR18), .ZN(_03477_) );
  AND2_X1 U17604 ( .A1(_02715__PTR21), .A2(_02715__PTR20), .ZN(_03478_) );
  AND2_X1 U17605 ( .A1(_02715__PTR23), .A2(_02715__PTR22), .ZN(_03479_) );
  AND2_X1 U17606 ( .A1(_02715__PTR25), .A2(_02715__PTR24), .ZN(_03480_) );
  AND2_X1 U17607 ( .A1(_02715__PTR27), .A2(_02715__PTR26), .ZN(_03481_) );
  AND2_X1 U17608 ( .A1(_02715__PTR29), .A2(_02715__PTR28), .ZN(_03482_) );
  AND2_X1 U17609 ( .A1(_02713__PTR31), .A2(_02715__PTR30), .ZN(_03483_) );
  AND2_X1 U17610 ( .A1(_03471_), .A2(_03470_), .ZN(_03484_) );
  AND2_X1 U17611 ( .A1(_03473_), .A2(_03472_), .ZN(_03485_) );
  AND2_X1 U17612 ( .A1(_03475_), .A2(_03474_), .ZN(_03486_) );
  AND2_X1 U17613 ( .A1(_03477_), .A2(_03476_), .ZN(_03487_) );
  AND2_X1 U17614 ( .A1(_03479_), .A2(_03478_), .ZN(_03488_) );
  AND2_X1 U17615 ( .A1(_03481_), .A2(_03480_), .ZN(_03489_) );
  AND2_X1 U17616 ( .A1(_03483_), .A2(_03482_), .ZN(_03490_) );
  AND2_X1 U17617 ( .A1(_03486_), .A2(_03485_), .ZN(_03491_) );
  AND2_X1 U17618 ( .A1(_03488_), .A2(_03487_), .ZN(_03492_) );
  AND2_X1 U17619 ( .A1(_03490_), .A2(_03489_), .ZN(_03493_) );
  AND2_X1 U17620 ( .A1(_03493_), .A2(_03492_), .ZN(_03494_) );
  OR2_X1 U17621 ( .A1(_01892__PTR131), .A2(_03440_), .ZN(_03495_) );
  OR2_X1 U17622 ( .A1(_01892__PTR133), .A2(_03441_), .ZN(_03496_) );
  OR2_X1 U17623 ( .A1(_01892__PTR135), .A2(_03442_), .ZN(_03497_) );
  OR2_X1 U17624 ( .A1(_01892__PTR137), .A2(_03443_), .ZN(_03498_) );
  OR2_X1 U17625 ( .A1(_01892__PTR139), .A2(_03444_), .ZN(_03499_) );
  OR2_X1 U17626 ( .A1(_01892__PTR141), .A2(_03445_), .ZN(_03500_) );
  OR2_X1 U17627 ( .A1(_01892__PTR143), .A2(_03446_), .ZN(_03501_) );
  OR2_X1 U17628 ( .A1(_01892__PTR145), .A2(_03447_), .ZN(_03502_) );
  OR2_X1 U17629 ( .A1(_01892__PTR147), .A2(_03448_), .ZN(_03503_) );
  OR2_X1 U17630 ( .A1(_01892__PTR149), .A2(_03449_), .ZN(_03504_) );
  OR2_X1 U17631 ( .A1(_01892__PTR151), .A2(_03450_), .ZN(_03505_) );
  OR2_X1 U17632 ( .A1(_01892__PTR153), .A2(_03451_), .ZN(_03506_) );
  OR2_X1 U17633 ( .A1(_01892__PTR155), .A2(_03452_), .ZN(_03507_) );
  OR2_X1 U17634 ( .A1(_01892__PTR157), .A2(_03453_), .ZN(_03508_) );
  OR2_X1 U17635 ( .A1(_03495_), .A2(_03455_), .ZN(_02714__PTR3) );
  OR2_X1 U17636 ( .A1(_03497_), .A2(_03456_), .ZN(_03509_) );
  OR2_X1 U17637 ( .A1(_03499_), .A2(_03457_), .ZN(_03510_) );
  OR2_X1 U17638 ( .A1(_03501_), .A2(_03458_), .ZN(_03511_) );
  OR2_X1 U17639 ( .A1(_03503_), .A2(_03459_), .ZN(_03512_) );
  OR2_X1 U17640 ( .A1(_03505_), .A2(_03460_), .ZN(_03513_) );
  OR2_X1 U17641 ( .A1(_03507_), .A2(_03461_), .ZN(_03514_) );
  OR2_X1 U17642 ( .A1(_03454_), .A2(_03462_), .ZN(_03515_) );
  OR2_X1 U17643 ( .A1(_03509_), .A2(_03463_), .ZN(_02714__PTR7) );
  OR2_X1 U17644 ( .A1(_03511_), .A2(_03464_), .ZN(_03516_) );
  OR2_X1 U17645 ( .A1(_03513_), .A2(_03465_), .ZN(_03517_) );
  OR2_X1 U17646 ( .A1(_03515_), .A2(_03466_), .ZN(_03518_) );
  OR2_X1 U17647 ( .A1(_03516_), .A2(_03467_), .ZN(_02714__PTR15) );
  OR2_X1 U17648 ( .A1(_03518_), .A2(_03468_), .ZN(_03519_) );
  OR2_X1 U17649 ( .A1(_03519_), .A2(_03469_), .ZN(_02714__PTR31) );
  AND2_X1 U17650 ( .A1(P1_P1_PhyAddrPointer_PTR3), .A2(P1_P1_PhyAddrPointer_PTR2), .ZN(_02794__PTR1) );
  AND2_X1 U17651 ( .A1(_03763_), .A2(_02794__PTR1), .ZN(_02794__PTR3) );
  AND2_X1 U17652 ( .A1(_03776_), .A2(_02794__PTR3), .ZN(_02794__PTR7) );
  AND2_X1 U17653 ( .A1(_03782_), .A2(_02794__PTR7), .ZN(_02794__PTR15) );
  AND2_X1 U17654 ( .A1(P1_P1_PhyAddrPointer_PTR5), .A2(P1_P1_PhyAddrPointer_PTR4), .ZN(_03763_) );
  AND2_X1 U17655 ( .A1(P1_P1_PhyAddrPointer_PTR7), .A2(P1_P1_PhyAddrPointer_PTR6), .ZN(_03764_) );
  AND2_X1 U17656 ( .A1(P1_P1_PhyAddrPointer_PTR9), .A2(P1_P1_PhyAddrPointer_PTR8), .ZN(_03765_) );
  AND2_X1 U17657 ( .A1(P1_P1_PhyAddrPointer_PTR11), .A2(P1_P1_PhyAddrPointer_PTR10), .ZN(_03766_) );
  AND2_X1 U17658 ( .A1(P1_P1_PhyAddrPointer_PTR13), .A2(P1_P1_PhyAddrPointer_PTR12), .ZN(_03767_) );
  AND2_X1 U17659 ( .A1(P1_P1_PhyAddrPointer_PTR15), .A2(P1_P1_PhyAddrPointer_PTR14), .ZN(_03768_) );
  AND2_X1 U17660 ( .A1(P1_P1_PhyAddrPointer_PTR17), .A2(P1_P1_PhyAddrPointer_PTR16), .ZN(_03769_) );
  AND2_X1 U17661 ( .A1(P1_P1_PhyAddrPointer_PTR19), .A2(P1_P1_PhyAddrPointer_PTR18), .ZN(_03770_) );
  AND2_X1 U17662 ( .A1(P1_P1_PhyAddrPointer_PTR21), .A2(P1_P1_PhyAddrPointer_PTR20), .ZN(_03771_) );
  AND2_X1 U17663 ( .A1(P1_P1_PhyAddrPointer_PTR23), .A2(P1_P1_PhyAddrPointer_PTR22), .ZN(_03772_) );
  AND2_X1 U17664 ( .A1(P1_P1_PhyAddrPointer_PTR25), .A2(P1_P1_PhyAddrPointer_PTR24), .ZN(_03773_) );
  AND2_X1 U17665 ( .A1(P1_P1_PhyAddrPointer_PTR27), .A2(P1_P1_PhyAddrPointer_PTR26), .ZN(_03774_) );
  AND2_X1 U17666 ( .A1(P1_P1_PhyAddrPointer_PTR29), .A2(P1_P1_PhyAddrPointer_PTR28), .ZN(_03775_) );
  AND2_X1 U17667 ( .A1(_03765_), .A2(_03764_), .ZN(_03776_) );
  AND2_X1 U17668 ( .A1(_03767_), .A2(_03766_), .ZN(_03777_) );
  AND2_X1 U17669 ( .A1(_03769_), .A2(_03768_), .ZN(_03778_) );
  AND2_X1 U17670 ( .A1(_03771_), .A2(_03770_), .ZN(_03779_) );
  AND2_X1 U17671 ( .A1(_03773_), .A2(_03772_), .ZN(_03780_) );
  AND2_X1 U17672 ( .A1(_03775_), .A2(_03774_), .ZN(_03781_) );
  AND2_X1 U17673 ( .A1(_03778_), .A2(_03777_), .ZN(_03782_) );
  AND2_X1 U17674 ( .A1(_03780_), .A2(_03779_), .ZN(_03783_) );
  AND2_X1 U17675 ( .A1(_03783_), .A2(_02794__PTR15), .ZN(_02794__PTR23) );
  AND2_X1 U17676 ( .A1(_03777_), .A2(_02794__PTR7), .ZN(_02794__PTR11) );
  AND2_X1 U17677 ( .A1(_03779_), .A2(_02794__PTR15), .ZN(_02794__PTR19) );
  AND2_X1 U17678 ( .A1(_03781_), .A2(_02794__PTR23), .ZN(_02794__PTR27) );
  AND2_X1 U17679 ( .A1(_03764_), .A2(_02794__PTR3), .ZN(_02794__PTR5) );
  AND2_X1 U17680 ( .A1(_03766_), .A2(_02794__PTR7), .ZN(_02794__PTR9) );
  AND2_X1 U17681 ( .A1(_03768_), .A2(_02794__PTR11), .ZN(_02794__PTR13) );
  AND2_X1 U17682 ( .A1(_03770_), .A2(_02794__PTR15), .ZN(_02794__PTR17) );
  AND2_X1 U17683 ( .A1(_03772_), .A2(_02794__PTR19), .ZN(_02794__PTR21) );
  AND2_X1 U17684 ( .A1(_03774_), .A2(_02794__PTR23), .ZN(_02794__PTR25) );
  AND2_X1 U17685 ( .A1(P1_P1_PhyAddrPointer_PTR4), .A2(_02794__PTR1), .ZN(_02794__PTR2) );
  AND2_X1 U17686 ( .A1(P1_P1_PhyAddrPointer_PTR6), .A2(_02794__PTR3), .ZN(_02794__PTR4) );
  AND2_X1 U17687 ( .A1(P1_P1_PhyAddrPointer_PTR8), .A2(_02794__PTR5), .ZN(_02794__PTR6) );
  AND2_X1 U17688 ( .A1(P1_P1_PhyAddrPointer_PTR10), .A2(_02794__PTR7), .ZN(_02794__PTR8) );
  AND2_X1 U17689 ( .A1(P1_P1_PhyAddrPointer_PTR12), .A2(_02794__PTR9), .ZN(_02794__PTR10) );
  AND2_X1 U17690 ( .A1(P1_P1_PhyAddrPointer_PTR14), .A2(_02794__PTR11), .ZN(_02794__PTR12) );
  AND2_X1 U17691 ( .A1(P1_P1_PhyAddrPointer_PTR16), .A2(_02794__PTR13), .ZN(_02794__PTR14) );
  AND2_X1 U17692 ( .A1(P1_P1_PhyAddrPointer_PTR18), .A2(_02794__PTR15), .ZN(_02794__PTR16) );
  AND2_X1 U17693 ( .A1(P1_P1_PhyAddrPointer_PTR20), .A2(_02794__PTR17), .ZN(_02794__PTR18) );
  AND2_X1 U17694 ( .A1(P1_P1_PhyAddrPointer_PTR22), .A2(_02794__PTR19), .ZN(_02794__PTR20) );
  AND2_X1 U17695 ( .A1(P1_P1_PhyAddrPointer_PTR24), .A2(_02794__PTR21), .ZN(_02794__PTR22) );
  AND2_X1 U17696 ( .A1(P1_P1_PhyAddrPointer_PTR26), .A2(_02794__PTR23), .ZN(_02794__PTR24) );
  AND2_X1 U17697 ( .A1(P1_P1_PhyAddrPointer_PTR28), .A2(_02794__PTR25), .ZN(_02794__PTR26) );
  AND2_X1 U17698 ( .A1(P1_P1_PhyAddrPointer_PTR30), .A2(_02794__PTR27), .ZN(_02794__PTR28) );
  AND2_X1 U17699 ( .A1(P1_P1_InstQueueWr_Addr_PTR1), .A2(P1_P1_InstQueueWr_Addr_PTR0), .ZN(_02779__PTR1) );
  AND2_X1 U17700 ( .A1(P1_P1_InstQueueWr_Addr_PTR2), .A2(_02779__PTR1), .ZN(_02779__PTR2) );
  AND2_X1 U17701 ( .A1(_01836__PTR1), .A2(_01836__PTR0), .ZN(_02780__PTR1) );
  AND2_X1 U17702 ( .A1(_01836__PTR2), .A2(_02780__PTR1), .ZN(_02780__PTR2) );
  AND2_X1 U17703 ( .A1(_01838__PTR1), .A2(P1_P1_InstQueueWr_Addr_PTR0), .ZN(_02785__PTR1) );
  AND2_X1 U17704 ( .A1(_01838__PTR2), .A2(_02785__PTR1), .ZN(_02785__PTR2) );
  AND2_X1 U17705 ( .A1(_01840__PTR1), .A2(_01836__PTR0), .ZN(_02790__PTR1) );
  AND2_X1 U17706 ( .A1(_01840__PTR2), .A2(_02790__PTR1), .ZN(_02790__PTR2) );
  AND2_X1 U17707 ( .A1(di1_PTR25), .A2(_02787__PTR0), .ZN(_02787__PTR1) );
  AND2_X1 U17708 ( .A1(_03740_), .A2(_02787__PTR1), .ZN(_02787__PTR3) );
  AND2_X1 U17709 ( .A1(_03741_), .A2(_02787__PTR3), .ZN(_02787__PTR5) );
  AND2_X1 U17710 ( .A1(di1_PTR26), .A2(_02787__PTR1), .ZN(_02787__PTR2) );
  AND2_X1 U17711 ( .A1(di1_PTR28), .A2(_02787__PTR3), .ZN(_02787__PTR4) );
  AND2_X1 U17712 ( .A1(di1_PTR30), .A2(_02787__PTR5), .ZN(_02787__PTR6) );
  AND2_X1 U17713 ( .A1(di1_PTR17), .A2(_02782__PTR0), .ZN(_02782__PTR1) );
  AND2_X1 U17714 ( .A1(_03738_), .A2(_02782__PTR1), .ZN(_02782__PTR3) );
  AND2_X1 U17715 ( .A1(di1_PTR19), .A2(di1_PTR18), .ZN(_03738_) );
  AND2_X1 U17716 ( .A1(di1_PTR21), .A2(di1_PTR20), .ZN(_03739_) );
  AND2_X1 U17717 ( .A1(di1_PTR27), .A2(di1_PTR26), .ZN(_03740_) );
  AND2_X1 U17718 ( .A1(di1_PTR29), .A2(di1_PTR28), .ZN(_03741_) );
  AND2_X1 U17719 ( .A1(_03739_), .A2(_02782__PTR3), .ZN(_02782__PTR5) );
  AND2_X1 U17720 ( .A1(di1_PTR18), .A2(_02782__PTR1), .ZN(_02782__PTR2) );
  AND2_X1 U17721 ( .A1(di1_PTR20), .A2(_02782__PTR3), .ZN(_02782__PTR4) );
  AND2_X1 U17722 ( .A1(di1_PTR22), .A2(_02782__PTR5), .ZN(_02782__PTR6) );
  AND2_X1 U17723 ( .A1(P1_rEIP_PTR2), .A2(_02778__PTR0), .ZN(_02778__PTR1) );
  AND2_X1 U17724 ( .A1(_03716_), .A2(_02778__PTR1), .ZN(_02778__PTR3) );
  AND2_X1 U17725 ( .A1(_03730_), .A2(_02778__PTR3), .ZN(_02778__PTR7) );
  AND2_X1 U17726 ( .A1(_03736_), .A2(_02778__PTR7), .ZN(_02778__PTR15) );
  AND2_X1 U17727 ( .A1(_03718_), .A2(_03717_), .ZN(_03730_) );
  AND2_X1 U17728 ( .A1(_03720_), .A2(_03719_), .ZN(_03731_) );
  AND2_X1 U17729 ( .A1(_03728_), .A2(_03727_), .ZN(_03735_) );
  AND2_X1 U17730 ( .A1(_03732_), .A2(_03731_), .ZN(_03736_) );
  AND2_X1 U17731 ( .A1(_03734_), .A2(_03733_), .ZN(_03737_) );
  AND2_X1 U17732 ( .A1(_03737_), .A2(_02778__PTR15), .ZN(_02778__PTR23) );
  AND2_X1 U17733 ( .A1(_03731_), .A2(_02778__PTR7), .ZN(_02778__PTR11) );
  AND2_X1 U17734 ( .A1(_03733_), .A2(_02778__PTR15), .ZN(_02778__PTR19) );
  AND2_X1 U17735 ( .A1(_03735_), .A2(_02778__PTR23), .ZN(_02778__PTR27) );
  AND2_X1 U17736 ( .A1(_03717_), .A2(_02778__PTR3), .ZN(_02778__PTR5) );
  AND2_X1 U17737 ( .A1(_03719_), .A2(_02778__PTR7), .ZN(_02778__PTR9) );
  AND2_X1 U17738 ( .A1(_03721_), .A2(_02778__PTR11), .ZN(_02778__PTR13) );
  AND2_X1 U17739 ( .A1(_03723_), .A2(_02778__PTR15), .ZN(_02778__PTR17) );
  AND2_X1 U17740 ( .A1(_03725_), .A2(_02778__PTR19), .ZN(_02778__PTR21) );
  AND2_X1 U17741 ( .A1(_03727_), .A2(_02778__PTR23), .ZN(_02778__PTR25) );
  AND2_X1 U17742 ( .A1(P1_rEIP_PTR3), .A2(_02778__PTR1), .ZN(_02778__PTR2) );
  AND2_X1 U17743 ( .A1(P1_rEIP_PTR5), .A2(_02778__PTR3), .ZN(_02778__PTR4) );
  AND2_X1 U17744 ( .A1(P1_rEIP_PTR7), .A2(_02778__PTR5), .ZN(_02778__PTR6) );
  AND2_X1 U17745 ( .A1(P1_rEIP_PTR9), .A2(_02778__PTR7), .ZN(_02778__PTR8) );
  AND2_X1 U17746 ( .A1(P1_rEIP_PTR11), .A2(_02778__PTR9), .ZN(_02778__PTR10) );
  AND2_X1 U17747 ( .A1(P1_rEIP_PTR13), .A2(_02778__PTR11), .ZN(_02778__PTR12) );
  AND2_X1 U17748 ( .A1(P1_rEIP_PTR15), .A2(_02778__PTR13), .ZN(_02778__PTR14) );
  AND2_X1 U17749 ( .A1(P1_rEIP_PTR17), .A2(_02778__PTR15), .ZN(_02778__PTR16) );
  AND2_X1 U17750 ( .A1(P1_rEIP_PTR19), .A2(_02778__PTR17), .ZN(_02778__PTR18) );
  AND2_X1 U17751 ( .A1(P1_rEIP_PTR21), .A2(_02778__PTR19), .ZN(_02778__PTR20) );
  AND2_X1 U17752 ( .A1(P1_rEIP_PTR23), .A2(_02778__PTR21), .ZN(_02778__PTR22) );
  AND2_X1 U17753 ( .A1(P1_rEIP_PTR25), .A2(_02778__PTR23), .ZN(_02778__PTR24) );
  AND2_X1 U17754 ( .A1(P1_rEIP_PTR27), .A2(_02778__PTR25), .ZN(_02778__PTR26) );
  AND2_X1 U17755 ( .A1(P1_rEIP_PTR29), .A2(_02778__PTR27), .ZN(_02778__PTR28) );
  AND2_X1 U17756 ( .A1(P1_rEIP_PTR3), .A2(_02793__PTR0), .ZN(_02793__PTR1) );
  AND2_X1 U17757 ( .A1(_03742_), .A2(_02793__PTR1), .ZN(_02793__PTR3) );
  AND2_X1 U17758 ( .A1(_03755_), .A2(_02793__PTR3), .ZN(_02793__PTR7) );
  AND2_X1 U17759 ( .A1(_03761_), .A2(_02793__PTR7), .ZN(_02793__PTR15) );
  AND2_X1 U17760 ( .A1(P1_rEIP_PTR5), .A2(P1_rEIP_PTR4), .ZN(_03742_) );
  AND2_X1 U17761 ( .A1(P1_rEIP_PTR7), .A2(P1_rEIP_PTR6), .ZN(_03743_) );
  AND2_X1 U17762 ( .A1(P1_rEIP_PTR9), .A2(P1_rEIP_PTR8), .ZN(_03744_) );
  AND2_X1 U17763 ( .A1(P1_rEIP_PTR11), .A2(P1_rEIP_PTR10), .ZN(_03745_) );
  AND2_X1 U17764 ( .A1(P1_rEIP_PTR13), .A2(P1_rEIP_PTR12), .ZN(_03746_) );
  AND2_X1 U17765 ( .A1(P1_rEIP_PTR15), .A2(P1_rEIP_PTR14), .ZN(_03747_) );
  AND2_X1 U17766 ( .A1(P1_rEIP_PTR17), .A2(P1_rEIP_PTR16), .ZN(_03748_) );
  AND2_X1 U17767 ( .A1(P1_rEIP_PTR19), .A2(P1_rEIP_PTR18), .ZN(_03749_) );
  AND2_X1 U17768 ( .A1(P1_rEIP_PTR21), .A2(P1_rEIP_PTR20), .ZN(_03750_) );
  AND2_X1 U17769 ( .A1(P1_rEIP_PTR23), .A2(P1_rEIP_PTR22), .ZN(_03751_) );
  AND2_X1 U17770 ( .A1(P1_rEIP_PTR25), .A2(P1_rEIP_PTR24), .ZN(_03752_) );
  AND2_X1 U17771 ( .A1(P1_rEIP_PTR27), .A2(P1_rEIP_PTR26), .ZN(_03753_) );
  AND2_X1 U17772 ( .A1(P1_rEIP_PTR29), .A2(P1_rEIP_PTR28), .ZN(_03754_) );
  AND2_X1 U17773 ( .A1(_03744_), .A2(_03743_), .ZN(_03755_) );
  AND2_X1 U17774 ( .A1(_03746_), .A2(_03745_), .ZN(_03756_) );
  AND2_X1 U17775 ( .A1(_03748_), .A2(_03747_), .ZN(_03757_) );
  AND2_X1 U17776 ( .A1(_03750_), .A2(_03749_), .ZN(_03758_) );
  AND2_X1 U17777 ( .A1(_03752_), .A2(_03751_), .ZN(_03759_) );
  AND2_X1 U17778 ( .A1(_03754_), .A2(_03753_), .ZN(_03760_) );
  AND2_X1 U17779 ( .A1(_03757_), .A2(_03756_), .ZN(_03761_) );
  AND2_X1 U17780 ( .A1(_03759_), .A2(_03758_), .ZN(_03762_) );
  AND2_X1 U17781 ( .A1(_03762_), .A2(_02793__PTR15), .ZN(_02793__PTR23) );
  AND2_X1 U17782 ( .A1(_03756_), .A2(_02793__PTR7), .ZN(_02793__PTR11) );
  AND2_X1 U17783 ( .A1(_03758_), .A2(_02793__PTR15), .ZN(_02793__PTR19) );
  AND2_X1 U17784 ( .A1(_03760_), .A2(_02793__PTR23), .ZN(_02793__PTR27) );
  AND2_X1 U17785 ( .A1(_03743_), .A2(_02793__PTR3), .ZN(_02793__PTR5) );
  AND2_X1 U17786 ( .A1(_03745_), .A2(_02793__PTR7), .ZN(_02793__PTR9) );
  AND2_X1 U17787 ( .A1(_03747_), .A2(_02793__PTR11), .ZN(_02793__PTR13) );
  AND2_X1 U17788 ( .A1(_03749_), .A2(_02793__PTR15), .ZN(_02793__PTR17) );
  AND2_X1 U17789 ( .A1(_03751_), .A2(_02793__PTR19), .ZN(_02793__PTR21) );
  AND2_X1 U17790 ( .A1(_03753_), .A2(_02793__PTR23), .ZN(_02793__PTR25) );
  AND2_X1 U17791 ( .A1(P1_rEIP_PTR4), .A2(_02793__PTR1), .ZN(_02793__PTR2) );
  AND2_X1 U17792 ( .A1(P1_rEIP_PTR6), .A2(_02793__PTR3), .ZN(_02793__PTR4) );
  AND2_X1 U17793 ( .A1(P1_rEIP_PTR8), .A2(_02793__PTR5), .ZN(_02793__PTR6) );
  AND2_X1 U17794 ( .A1(P1_rEIP_PTR10), .A2(_02793__PTR7), .ZN(_02793__PTR8) );
  AND2_X1 U17795 ( .A1(P1_rEIP_PTR12), .A2(_02793__PTR9), .ZN(_02793__PTR10) );
  AND2_X1 U17796 ( .A1(P1_rEIP_PTR14), .A2(_02793__PTR11), .ZN(_02793__PTR12) );
  AND2_X1 U17797 ( .A1(P1_rEIP_PTR16), .A2(_02793__PTR13), .ZN(_02793__PTR14) );
  AND2_X1 U17798 ( .A1(P1_rEIP_PTR18), .A2(_02793__PTR15), .ZN(_02793__PTR16) );
  AND2_X1 U17799 ( .A1(P1_rEIP_PTR20), .A2(_02793__PTR17), .ZN(_02793__PTR18) );
  AND2_X1 U17800 ( .A1(P1_rEIP_PTR22), .A2(_02793__PTR19), .ZN(_02793__PTR20) );
  AND2_X1 U17801 ( .A1(P1_rEIP_PTR24), .A2(_02793__PTR21), .ZN(_02793__PTR22) );
  AND2_X1 U17802 ( .A1(P1_rEIP_PTR26), .A2(_02793__PTR23), .ZN(_02793__PTR24) );
  AND2_X1 U17803 ( .A1(P1_rEIP_PTR28), .A2(_02793__PTR25), .ZN(_02793__PTR26) );
  AND2_X1 U17804 ( .A1(P1_rEIP_PTR30), .A2(_02793__PTR27), .ZN(_02793__PTR28) );
  AND2_X1 U17805 ( .A1(_02996__PTR4), .A2(_02995__PTR3), .ZN(_02998_) );
  OR2_X1 U17806 ( .A1(P2_P1_InstQueueRd_Addr_PTR4), .A2(_02998_), .ZN(_02995__PTR4) );
  AND2_X1 U17807 ( .A1(_02224__PTR59), .A2(_02991__PTR2), .ZN(_04357_) );
  AND2_X1 U17808 ( .A1(_03188__PTR4), .A2(_03189__PTR3), .ZN(_02992__PTR5) );
  OR2_X1 U17809 ( .A1(_04363_), .A2(_04360_), .ZN(_03189__PTR3) );
  AND2_X1 U17810 ( .A1(_02991__PTR1), .A2(_02991__PTR0), .ZN(_02993__PTR1) );
  AND2_X1 U17811 ( .A1(_02992__PTR5), .A2(_02991__PTR4), .ZN(_04358_) );
  AND2_X1 U17812 ( .A1(_04360_), .A2(_02993__PTR1), .ZN(_04359_) );
  AND2_X1 U17813 ( .A1(_02224__PTR59), .A2(_02224__PTR58), .ZN(_04360_) );
  AND2_X1 U17814 ( .A1(_02992__PTR5), .A2(_02994__PTR4), .ZN(_04361_) );
  AND2_X1 U17815 ( .A1(_04361_), .A2(_02993__PTR3), .ZN(_04362_) );
  OR2_X1 U17816 ( .A1(_02991__PTR3), .A2(_04357_), .ZN(_04363_) );
  OR2_X1 U17817 ( .A1(_04363_), .A2(_04359_), .ZN(_02993__PTR3) );
  OR2_X1 U17818 ( .A1(_04358_), .A2(_04362_), .ZN(_02186__PTR28) );
  AND2_X1 U17819 ( .A1(_03074__PTR1), .A2(P2_P1_InstAddrPointer_PTR0), .ZN(_03075__PTR1) );
  AND2_X1 U17820 ( .A1(_02990__PTR3), .A2(_02990__PTR2), .ZN(_04292_) );
  AND2_X1 U17821 ( .A1(_02990__PTR5), .A2(_02990__PTR4), .ZN(_04307_) );
  AND2_X1 U17822 ( .A1(_02990__PTR7), .A2(_02990__PTR6), .ZN(_04308_) );
  AND2_X1 U17823 ( .A1(_02990__PTR9), .A2(_02990__PTR8), .ZN(_04309_) );
  AND2_X1 U17824 ( .A1(_02990__PTR15), .A2(_02990__PTR14), .ZN(_04312_) );
  AND2_X1 U17825 ( .A1(_02990__PTR17), .A2(_02990__PTR16), .ZN(_04313_) );
  AND2_X1 U17826 ( .A1(_02990__PTR19), .A2(_02990__PTR18), .ZN(_04314_) );
  AND2_X1 U17827 ( .A1(_02990__PTR21), .A2(_02990__PTR20), .ZN(_04315_) );
  AND2_X1 U17828 ( .A1(_02990__PTR23), .A2(_02990__PTR22), .ZN(_04316_) );
  AND2_X1 U17829 ( .A1(_02990__PTR25), .A2(_02990__PTR24), .ZN(_04317_) );
  AND2_X1 U17830 ( .A1(_02990__PTR27), .A2(_02990__PTR26), .ZN(_04318_) );
  AND2_X1 U17831 ( .A1(_02990__PTR29), .A2(_02990__PTR28), .ZN(_04319_) );
  AND2_X1 U17832 ( .A1(_02988__PTR31), .A2(_02990__PTR30), .ZN(_04320_) );
  AND2_X1 U17833 ( .A1(_04308_), .A2(_04307_), .ZN(_04321_) );
  AND2_X1 U17834 ( .A1(_04312_), .A2(_04311_), .ZN(_04323_) );
  AND2_X1 U17835 ( .A1(_04314_), .A2(_04313_), .ZN(_04324_) );
  AND2_X1 U17836 ( .A1(_04316_), .A2(_04315_), .ZN(_04325_) );
  AND2_X1 U17837 ( .A1(_04318_), .A2(_04317_), .ZN(_04326_) );
  AND2_X1 U17838 ( .A1(_04320_), .A2(_04319_), .ZN(_04327_) );
  AND2_X1 U17839 ( .A1(_04323_), .A2(_04322_), .ZN(_04328_) );
  AND2_X1 U17840 ( .A1(_04325_), .A2(_04324_), .ZN(_04329_) );
  AND2_X1 U17841 ( .A1(_02990__PTR3), .A2(P2_P1_InstAddrPointer_PTR2), .ZN(_04277_) );
  AND2_X1 U17842 ( .A1(_02990__PTR5), .A2(P2_P1_InstAddrPointer_PTR4), .ZN(_04278_) );
  AND2_X1 U17843 ( .A1(_02990__PTR7), .A2(P2_P1_InstAddrPointer_PTR6), .ZN(_04279_) );
  AND2_X1 U17844 ( .A1(_02990__PTR9), .A2(P2_P1_InstAddrPointer_PTR8), .ZN(_04280_) );
  AND2_X1 U17845 ( .A1(_02990__PTR11), .A2(P2_P1_InstAddrPointer_PTR10), .ZN(_04281_) );
  AND2_X1 U17846 ( .A1(_02990__PTR13), .A2(P2_P1_InstAddrPointer_PTR12), .ZN(_04282_) );
  AND2_X1 U17847 ( .A1(_02990__PTR15), .A2(P2_P1_InstAddrPointer_PTR14), .ZN(_04283_) );
  AND2_X1 U17848 ( .A1(_02990__PTR17), .A2(P2_P1_InstAddrPointer_PTR16), .ZN(_04284_) );
  AND2_X1 U17849 ( .A1(_02990__PTR19), .A2(P2_P1_InstAddrPointer_PTR18), .ZN(_04285_) );
  AND2_X1 U17850 ( .A1(_02990__PTR21), .A2(P2_P1_InstAddrPointer_PTR20), .ZN(_04286_) );
  AND2_X1 U17851 ( .A1(_02990__PTR23), .A2(P2_P1_InstAddrPointer_PTR22), .ZN(_04287_) );
  AND2_X1 U17852 ( .A1(_02990__PTR25), .A2(P2_P1_InstAddrPointer_PTR24), .ZN(_04288_) );
  AND2_X1 U17853 ( .A1(_02990__PTR27), .A2(P2_P1_InstAddrPointer_PTR26), .ZN(_04289_) );
  AND2_X1 U17854 ( .A1(_02990__PTR29), .A2(P2_P1_InstAddrPointer_PTR28), .ZN(_04290_) );
  AND2_X1 U17855 ( .A1(_02988__PTR31), .A2(P2_P1_InstAddrPointer_PTR30), .ZN(_04291_) );
  AND2_X1 U17856 ( .A1(_04308_), .A2(_04333_), .ZN(_04293_) );
  AND2_X1 U17857 ( .A1(_04310_), .A2(_04335_), .ZN(_04294_) );
  AND2_X1 U17858 ( .A1(_04312_), .A2(_04337_), .ZN(_04295_) );
  AND2_X1 U17859 ( .A1(_04314_), .A2(_04339_), .ZN(_04296_) );
  AND2_X1 U17860 ( .A1(_04316_), .A2(_04341_), .ZN(_04297_) );
  AND2_X1 U17861 ( .A1(_04318_), .A2(_04343_), .ZN(_04298_) );
  AND2_X1 U17862 ( .A1(_04320_), .A2(_04345_), .ZN(_04299_) );
  AND2_X1 U17863 ( .A1(_04321_), .A2(_02989__PTR3), .ZN(_04300_) );
  AND2_X1 U17864 ( .A1(_04323_), .A2(_04347_), .ZN(_04301_) );
  AND2_X1 U17865 ( .A1(_04325_), .A2(_04349_), .ZN(_04302_) );
  AND2_X1 U17866 ( .A1(_04327_), .A2(_04351_), .ZN(_04303_) );
  AND2_X1 U17867 ( .A1(_04328_), .A2(_02989__PTR7), .ZN(_04304_) );
  AND2_X1 U17868 ( .A1(_04330_), .A2(_04354_), .ZN(_04305_) );
  AND2_X1 U17869 ( .A1(_04331_), .A2(_02989__PTR15), .ZN(_04306_) );
  AND2_X1 U17870 ( .A1(_02990__PTR11), .A2(_02990__PTR10), .ZN(_04310_) );
  AND2_X1 U17871 ( .A1(_02990__PTR13), .A2(_02990__PTR12), .ZN(_04311_) );
  AND2_X1 U17872 ( .A1(_04310_), .A2(_04309_), .ZN(_04322_) );
  AND2_X1 U17873 ( .A1(_04327_), .A2(_04326_), .ZN(_04330_) );
  AND2_X1 U17874 ( .A1(_04330_), .A2(_04329_), .ZN(_04331_) );
  OR2_X1 U17875 ( .A1(P2_P1_InstAddrPointer_PTR3), .A2(_04277_), .ZN(_04332_) );
  OR2_X1 U17876 ( .A1(P2_P1_InstAddrPointer_PTR5), .A2(_04278_), .ZN(_04333_) );
  OR2_X1 U17877 ( .A1(P2_P1_InstAddrPointer_PTR7), .A2(_04279_), .ZN(_04334_) );
  OR2_X1 U17878 ( .A1(P2_P1_InstAddrPointer_PTR9), .A2(_04280_), .ZN(_04335_) );
  OR2_X1 U17879 ( .A1(P2_P1_InstAddrPointer_PTR11), .A2(_04281_), .ZN(_04336_) );
  OR2_X1 U17880 ( .A1(P2_P1_InstAddrPointer_PTR13), .A2(_04282_), .ZN(_04337_) );
  OR2_X1 U17881 ( .A1(P2_P1_InstAddrPointer_PTR15), .A2(_04283_), .ZN(_04338_) );
  OR2_X1 U17882 ( .A1(P2_P1_InstAddrPointer_PTR17), .A2(_04284_), .ZN(_04339_) );
  OR2_X1 U17883 ( .A1(P2_P1_InstAddrPointer_PTR19), .A2(_04285_), .ZN(_04340_) );
  OR2_X1 U17884 ( .A1(P2_P1_InstAddrPointer_PTR21), .A2(_04286_), .ZN(_04341_) );
  OR2_X1 U17885 ( .A1(P2_P1_InstAddrPointer_PTR23), .A2(_04287_), .ZN(_04342_) );
  OR2_X1 U17886 ( .A1(P2_P1_InstAddrPointer_PTR25), .A2(_04288_), .ZN(_04343_) );
  OR2_X1 U17887 ( .A1(P2_P1_InstAddrPointer_PTR27), .A2(_04289_), .ZN(_04344_) );
  OR2_X1 U17888 ( .A1(P2_P1_InstAddrPointer_PTR29), .A2(_04290_), .ZN(_04345_) );
  OR2_X1 U17889 ( .A1(_04332_), .A2(_04292_), .ZN(_02989__PTR3) );
  OR2_X1 U17890 ( .A1(_04334_), .A2(_04293_), .ZN(_04346_) );
  OR2_X1 U17891 ( .A1(_04336_), .A2(_04294_), .ZN(_04347_) );
  OR2_X1 U17892 ( .A1(_04338_), .A2(_04295_), .ZN(_04348_) );
  OR2_X1 U17893 ( .A1(_04340_), .A2(_04296_), .ZN(_04349_) );
  OR2_X1 U17894 ( .A1(_04342_), .A2(_04297_), .ZN(_04350_) );
  OR2_X1 U17895 ( .A1(_04344_), .A2(_04298_), .ZN(_04351_) );
  OR2_X1 U17896 ( .A1(_04291_), .A2(_04299_), .ZN(_04352_) );
  OR2_X1 U17897 ( .A1(_04346_), .A2(_04300_), .ZN(_02989__PTR7) );
  OR2_X1 U17898 ( .A1(_04348_), .A2(_04301_), .ZN(_04353_) );
  OR2_X1 U17899 ( .A1(_04350_), .A2(_04302_), .ZN(_04354_) );
  OR2_X1 U17900 ( .A1(_04352_), .A2(_04303_), .ZN(_04355_) );
  OR2_X1 U17901 ( .A1(_04353_), .A2(_04304_), .ZN(_02989__PTR15) );
  OR2_X1 U17902 ( .A1(_04355_), .A2(_04305_), .ZN(_04356_) );
  OR2_X1 U17903 ( .A1(_04356_), .A2(_04306_), .ZN(_02989__PTR31) );
  AND2_X1 U17904 ( .A1(_02224__PTR43), .A2(_02224__PTR42), .ZN(_04735_) );
  AND2_X1 U17905 ( .A1(_03186__PTR4), .A2(_03187__PTR3), .ZN(_02985__PTR5) );
  OR2_X1 U17906 ( .A1(_02986__PTR3), .A2(_04735_), .ZN(_03187__PTR3) );
  AND2_X1 U17907 ( .A1(_02985__PTR5), .A2(_02984__PTR4), .ZN(_04273_) );
  AND2_X1 U17908 ( .A1(_02224__PTR43), .A2(_02984__PTR2), .ZN(_04274_) );
  AND2_X1 U17909 ( .A1(_02985__PTR5), .A2(_02987__PTR4), .ZN(_04275_) );
  AND2_X1 U17910 ( .A1(_04275_), .A2(_02986__PTR3), .ZN(_04276_) );
  OR2_X1 U17911 ( .A1(_02984__PTR3), .A2(_04274_), .ZN(_02986__PTR3) );
  OR2_X1 U17912 ( .A1(_04273_), .A2(_04276_), .ZN(_02986__PTR5) );
  AND2_X1 U17913 ( .A1(_02982__PTR1), .A2(_02981__PTR0), .ZN(_04267_) );
  AND2_X1 U17914 ( .A1(_02982__PTR3), .A2(_02983__PTR2), .ZN(_04268_) );
  AND2_X1 U17915 ( .A1(_04270_), .A2(_02981__PTR1), .ZN(_04269_) );
  AND2_X1 U17916 ( .A1(_02982__PTR3), .A2(_02982__PTR2), .ZN(_04270_) );
  AND2_X1 U17917 ( .A1(_02982__PTR4), .A2(_02981__PTR3), .ZN(_04271_) );
  OR2_X1 U17918 ( .A1(_02983__PTR0), .A2(_02982__PTR0), .ZN(_02981__PTR0) );
  OR2_X1 U17919 ( .A1(_02983__PTR1), .A2(_04267_), .ZN(_02981__PTR1) );
  OR2_X1 U17920 ( .A1(_02983__PTR3), .A2(_04268_), .ZN(_04272_) );
  OR2_X1 U17921 ( .A1(_04272_), .A2(_04269_), .ZN(_02981__PTR3) );
  OR2_X1 U17922 ( .A1(_02983__PTR4), .A2(_04271_), .ZN(_02981__PTR4) );
  AND2_X1 U17923 ( .A1(P2_EBX_PTR1), .A2(P2_EBX_PTR0), .ZN(_03073__PTR1) );
  AND2_X1 U17924 ( .A1(_04603_), .A2(_03073__PTR1), .ZN(_03073__PTR3) );
  AND2_X1 U17925 ( .A1(_04617_), .A2(_03073__PTR3), .ZN(_03073__PTR7) );
  AND2_X1 U17926 ( .A1(_04623_), .A2(_03073__PTR7), .ZN(_03073__PTR15) );
  AND2_X1 U17927 ( .A1(P2_EBX_PTR3), .A2(P2_EBX_PTR2), .ZN(_04603_) );
  AND2_X1 U17928 ( .A1(P2_EBX_PTR5), .A2(P2_EBX_PTR4), .ZN(_04604_) );
  AND2_X1 U17929 ( .A1(P2_EBX_PTR7), .A2(P2_EBX_PTR6), .ZN(_04605_) );
  AND2_X1 U17930 ( .A1(P2_EBX_PTR9), .A2(P2_EBX_PTR8), .ZN(_04606_) );
  AND2_X1 U17931 ( .A1(P2_EBX_PTR11), .A2(P2_EBX_PTR10), .ZN(_04607_) );
  AND2_X1 U17932 ( .A1(P2_EBX_PTR13), .A2(P2_EBX_PTR12), .ZN(_04608_) );
  AND2_X1 U17933 ( .A1(P2_EBX_PTR15), .A2(P2_EBX_PTR14), .ZN(_04609_) );
  AND2_X1 U17934 ( .A1(P2_EBX_PTR17), .A2(P2_EBX_PTR16), .ZN(_04610_) );
  AND2_X1 U17935 ( .A1(P2_EBX_PTR19), .A2(P2_EBX_PTR18), .ZN(_04611_) );
  AND2_X1 U17936 ( .A1(P2_EBX_PTR21), .A2(P2_EBX_PTR20), .ZN(_04612_) );
  AND2_X1 U17937 ( .A1(P2_EBX_PTR23), .A2(P2_EBX_PTR22), .ZN(_04613_) );
  AND2_X1 U17938 ( .A1(P2_EBX_PTR25), .A2(P2_EBX_PTR24), .ZN(_04614_) );
  AND2_X1 U17939 ( .A1(P2_EBX_PTR27), .A2(P2_EBX_PTR26), .ZN(_04615_) );
  AND2_X1 U17940 ( .A1(P2_EBX_PTR29), .A2(P2_EBX_PTR28), .ZN(_04616_) );
  AND2_X1 U17941 ( .A1(_04605_), .A2(_04604_), .ZN(_04617_) );
  AND2_X1 U17942 ( .A1(_04607_), .A2(_04606_), .ZN(_04618_) );
  AND2_X1 U17943 ( .A1(_04609_), .A2(_04608_), .ZN(_04619_) );
  AND2_X1 U17944 ( .A1(_04611_), .A2(_04610_), .ZN(_04620_) );
  AND2_X1 U17945 ( .A1(_04613_), .A2(_04612_), .ZN(_04621_) );
  AND2_X1 U17946 ( .A1(_04615_), .A2(_04614_), .ZN(_04622_) );
  AND2_X1 U17947 ( .A1(_04619_), .A2(_04618_), .ZN(_04623_) );
  AND2_X1 U17948 ( .A1(_04621_), .A2(_04620_), .ZN(_04624_) );
  AND2_X1 U17949 ( .A1(_04624_), .A2(_03073__PTR15), .ZN(_03073__PTR23) );
  AND2_X1 U17950 ( .A1(_04618_), .A2(_03073__PTR7), .ZN(_03073__PTR11) );
  AND2_X1 U17951 ( .A1(_04620_), .A2(_03073__PTR15), .ZN(_03073__PTR19) );
  AND2_X1 U17952 ( .A1(_04622_), .A2(_03073__PTR23), .ZN(_03073__PTR27) );
  AND2_X1 U17953 ( .A1(_04604_), .A2(_03073__PTR3), .ZN(_03073__PTR5) );
  AND2_X1 U17954 ( .A1(_04606_), .A2(_03073__PTR7), .ZN(_03073__PTR9) );
  AND2_X1 U17955 ( .A1(_04608_), .A2(_03073__PTR11), .ZN(_03073__PTR13) );
  AND2_X1 U17956 ( .A1(_04610_), .A2(_03073__PTR15), .ZN(_03073__PTR17) );
  AND2_X1 U17957 ( .A1(_04612_), .A2(_03073__PTR19), .ZN(_03073__PTR21) );
  AND2_X1 U17958 ( .A1(_04614_), .A2(_03073__PTR23), .ZN(_03073__PTR25) );
  AND2_X1 U17959 ( .A1(_04616_), .A2(_03073__PTR27), .ZN(_03073__PTR29) );
  AND2_X1 U17960 ( .A1(P2_EBX_PTR2), .A2(_03073__PTR1), .ZN(_03073__PTR2) );
  AND2_X1 U17961 ( .A1(P2_EBX_PTR4), .A2(_03073__PTR3), .ZN(_03073__PTR4) );
  AND2_X1 U17962 ( .A1(P2_EBX_PTR6), .A2(_03073__PTR5), .ZN(_03073__PTR6) );
  AND2_X1 U17963 ( .A1(P2_EBX_PTR8), .A2(_03073__PTR7), .ZN(_03073__PTR8) );
  AND2_X1 U17964 ( .A1(P2_EBX_PTR10), .A2(_03073__PTR9), .ZN(_03073__PTR10) );
  AND2_X1 U17965 ( .A1(P2_EBX_PTR12), .A2(_03073__PTR11), .ZN(_03073__PTR12) );
  AND2_X1 U17966 ( .A1(P2_EBX_PTR14), .A2(_03073__PTR13), .ZN(_03073__PTR14) );
  AND2_X1 U17967 ( .A1(P2_EBX_PTR16), .A2(_03073__PTR15), .ZN(_03073__PTR16) );
  AND2_X1 U17968 ( .A1(P2_EBX_PTR18), .A2(_03073__PTR17), .ZN(_03073__PTR18) );
  AND2_X1 U17969 ( .A1(P2_EBX_PTR20), .A2(_03073__PTR19), .ZN(_03073__PTR20) );
  AND2_X1 U17970 ( .A1(P2_EBX_PTR22), .A2(_03073__PTR21), .ZN(_03073__PTR22) );
  AND2_X1 U17971 ( .A1(P2_EBX_PTR24), .A2(_03073__PTR23), .ZN(_03073__PTR24) );
  AND2_X1 U17972 ( .A1(P2_EBX_PTR26), .A2(_03073__PTR25), .ZN(_03073__PTR26) );
  AND2_X1 U17973 ( .A1(P2_EBX_PTR28), .A2(_03073__PTR27), .ZN(_03073__PTR28) );
  AND2_X1 U17974 ( .A1(P2_EBX_PTR30), .A2(_03073__PTR29), .ZN(_03073__PTR30) );
  AND2_X1 U17975 ( .A1(P2_EAX_PTR1), .A2(P2_EAX_PTR0), .ZN(_03072__PTR1) );
  AND2_X1 U17976 ( .A1(_04589_), .A2(_03072__PTR1), .ZN(_03072__PTR3) );
  AND2_X1 U17977 ( .A1(_04597_), .A2(_03072__PTR3), .ZN(_03072__PTR7) );
  AND2_X1 U17978 ( .A1(_04601_), .A2(_03072__PTR7), .ZN(_03072__PTR15) );
  AND2_X1 U17979 ( .A1(P2_EAX_PTR3), .A2(P2_EAX_PTR2), .ZN(_04589_) );
  AND2_X1 U17980 ( .A1(P2_EAX_PTR5), .A2(P2_EAX_PTR4), .ZN(_04590_) );
  AND2_X1 U17981 ( .A1(P2_EAX_PTR7), .A2(P2_EAX_PTR6), .ZN(_04591_) );
  AND2_X1 U17982 ( .A1(P2_EAX_PTR9), .A2(P2_EAX_PTR8), .ZN(_04592_) );
  AND2_X1 U17983 ( .A1(P2_EAX_PTR11), .A2(P2_EAX_PTR10), .ZN(_04593_) );
  AND2_X1 U17984 ( .A1(P2_EAX_PTR13), .A2(P2_EAX_PTR12), .ZN(_04594_) );
  AND2_X1 U17985 ( .A1(P2_EAX_PTR15), .A2(P2_EAX_PTR14), .ZN(_04595_) );
  AND2_X1 U17986 ( .A1(P2_EAX_PTR17), .A2(P2_EAX_PTR16), .ZN(_04596_) );
  AND2_X1 U17987 ( .A1(P2_EAX_PTR27), .A2(P2_EAX_PTR26), .ZN(_04585_) );
  AND2_X1 U17988 ( .A1(P2_EAX_PTR29), .A2(P2_EAX_PTR28), .ZN(_04586_) );
  AND2_X1 U17989 ( .A1(_04591_), .A2(_04590_), .ZN(_04597_) );
  AND2_X1 U17990 ( .A1(_04593_), .A2(_04592_), .ZN(_04598_) );
  AND2_X1 U17991 ( .A1(_04595_), .A2(_04594_), .ZN(_04599_) );
  AND2_X1 U17992 ( .A1(_04581_), .A2(_04596_), .ZN(_04600_) );
  AND2_X1 U17993 ( .A1(_04585_), .A2(_04584_), .ZN(_04588_) );
  AND2_X1 U17994 ( .A1(_04599_), .A2(_04598_), .ZN(_04601_) );
  AND2_X1 U17995 ( .A1(_04587_), .A2(_04600_), .ZN(_04602_) );
  AND2_X1 U17996 ( .A1(_04602_), .A2(_03072__PTR15), .ZN(_03072__PTR23) );
  AND2_X1 U17997 ( .A1(_04598_), .A2(_03072__PTR7), .ZN(_03072__PTR11) );
  AND2_X1 U17998 ( .A1(_04600_), .A2(_03072__PTR15), .ZN(_03072__PTR19) );
  AND2_X1 U17999 ( .A1(_04588_), .A2(_03072__PTR23), .ZN(_03072__PTR27) );
  AND2_X1 U18000 ( .A1(_04590_), .A2(_03072__PTR3), .ZN(_03072__PTR5) );
  AND2_X1 U18001 ( .A1(_04592_), .A2(_03072__PTR7), .ZN(_03072__PTR9) );
  AND2_X1 U18002 ( .A1(_04594_), .A2(_03072__PTR11), .ZN(_03072__PTR13) );
  AND2_X1 U18003 ( .A1(_04596_), .A2(_03072__PTR15), .ZN(_03072__PTR17) );
  AND2_X1 U18004 ( .A1(_04582_), .A2(_03072__PTR19), .ZN(_03072__PTR21) );
  AND2_X1 U18005 ( .A1(_04584_), .A2(_03072__PTR23), .ZN(_03072__PTR25) );
  AND2_X1 U18006 ( .A1(_04586_), .A2(_03072__PTR27), .ZN(_03072__PTR29) );
  AND2_X1 U18007 ( .A1(P2_EAX_PTR2), .A2(_03072__PTR1), .ZN(_03072__PTR2) );
  AND2_X1 U18008 ( .A1(P2_EAX_PTR4), .A2(_03072__PTR3), .ZN(_03072__PTR4) );
  AND2_X1 U18009 ( .A1(P2_EAX_PTR6), .A2(_03072__PTR5), .ZN(_03072__PTR6) );
  AND2_X1 U18010 ( .A1(P2_EAX_PTR8), .A2(_03072__PTR7), .ZN(_03072__PTR8) );
  AND2_X1 U18011 ( .A1(P2_EAX_PTR10), .A2(_03072__PTR9), .ZN(_03072__PTR10) );
  AND2_X1 U18012 ( .A1(P2_EAX_PTR12), .A2(_03072__PTR11), .ZN(_03072__PTR12) );
  AND2_X1 U18013 ( .A1(P2_EAX_PTR14), .A2(_03072__PTR13), .ZN(_03072__PTR14) );
  AND2_X1 U18014 ( .A1(P2_EAX_PTR16), .A2(_03072__PTR15), .ZN(_03072__PTR16) );
  AND2_X1 U18015 ( .A1(P2_EAX_PTR18), .A2(_03072__PTR17), .ZN(_03072__PTR18) );
  AND2_X1 U18016 ( .A1(P2_EAX_PTR20), .A2(_03072__PTR19), .ZN(_03072__PTR20) );
  AND2_X1 U18017 ( .A1(P2_EAX_PTR22), .A2(_03072__PTR21), .ZN(_03072__PTR22) );
  AND2_X1 U18018 ( .A1(P2_EAX_PTR24), .A2(_03072__PTR23), .ZN(_03072__PTR24) );
  AND2_X1 U18019 ( .A1(P2_EAX_PTR26), .A2(_03072__PTR25), .ZN(_03072__PTR26) );
  AND2_X1 U18020 ( .A1(P2_EAX_PTR28), .A2(_03072__PTR27), .ZN(_03072__PTR28) );
  AND2_X1 U18021 ( .A1(P2_EAX_PTR30), .A2(_03072__PTR29), .ZN(_03072__PTR30) );
  AND2_X1 U18022 ( .A1(P2_EAX_PTR17), .A2(_03069__PTR0), .ZN(_03069__PTR1) );
  AND2_X1 U18023 ( .A1(_04581_), .A2(_03069__PTR1), .ZN(_03069__PTR3) );
  AND2_X1 U18024 ( .A1(_04587_), .A2(_03069__PTR3), .ZN(_03069__PTR7) );
  AND2_X1 U18025 ( .A1(P2_EAX_PTR19), .A2(P2_EAX_PTR18), .ZN(_04581_) );
  AND2_X1 U18026 ( .A1(P2_EAX_PTR21), .A2(P2_EAX_PTR20), .ZN(_04582_) );
  AND2_X1 U18027 ( .A1(P2_EAX_PTR23), .A2(P2_EAX_PTR22), .ZN(_04583_) );
  AND2_X1 U18028 ( .A1(P2_EAX_PTR25), .A2(P2_EAX_PTR24), .ZN(_04584_) );
  AND2_X1 U18029 ( .A1(_04583_), .A2(_04582_), .ZN(_04587_) );
  AND2_X1 U18030 ( .A1(_04588_), .A2(_03069__PTR7), .ZN(_03069__PTR11) );
  AND2_X1 U18031 ( .A1(_04582_), .A2(_03069__PTR3), .ZN(_03069__PTR5) );
  AND2_X1 U18032 ( .A1(_04584_), .A2(_03069__PTR7), .ZN(_03069__PTR9) );
  AND2_X1 U18033 ( .A1(_04586_), .A2(_03069__PTR11), .ZN(_03069__PTR13) );
  AND2_X1 U18034 ( .A1(P2_EAX_PTR18), .A2(_03069__PTR1), .ZN(_03069__PTR2) );
  AND2_X1 U18035 ( .A1(P2_EAX_PTR20), .A2(_03069__PTR3), .ZN(_03069__PTR4) );
  AND2_X1 U18036 ( .A1(P2_EAX_PTR22), .A2(_03069__PTR5), .ZN(_03069__PTR6) );
  AND2_X1 U18037 ( .A1(P2_EAX_PTR24), .A2(_03069__PTR7), .ZN(_03069__PTR8) );
  AND2_X1 U18038 ( .A1(P2_EAX_PTR26), .A2(_03069__PTR9), .ZN(_03069__PTR10) );
  AND2_X1 U18039 ( .A1(P2_EAX_PTR28), .A2(_03069__PTR11), .ZN(_03069__PTR12) );
  AND2_X1 U18040 ( .A1(P2_rEIP_PTR2), .A2(P2_rEIP_PTR1), .ZN(_03066__PTR1) );
  AND2_X1 U18041 ( .A1(_04364_), .A2(_03066__PTR1), .ZN(_03066__PTR3) );
  AND2_X1 U18042 ( .A1(_04378_), .A2(_03066__PTR3), .ZN(_03066__PTR7) );
  AND2_X1 U18043 ( .A1(_04384_), .A2(_03066__PTR7), .ZN(_03066__PTR15) );
  AND2_X1 U18044 ( .A1(P2_rEIP_PTR4), .A2(P2_rEIP_PTR3), .ZN(_04364_) );
  AND2_X1 U18045 ( .A1(P2_rEIP_PTR6), .A2(P2_rEIP_PTR5), .ZN(_04365_) );
  AND2_X1 U18046 ( .A1(P2_rEIP_PTR10), .A2(P2_rEIP_PTR9), .ZN(_04367_) );
  AND2_X1 U18047 ( .A1(P2_rEIP_PTR12), .A2(P2_rEIP_PTR11), .ZN(_04368_) );
  AND2_X1 U18048 ( .A1(P2_rEIP_PTR14), .A2(P2_rEIP_PTR13), .ZN(_04369_) );
  AND2_X1 U18049 ( .A1(P2_rEIP_PTR18), .A2(P2_rEIP_PTR17), .ZN(_04371_) );
  AND2_X1 U18050 ( .A1(P2_rEIP_PTR22), .A2(P2_rEIP_PTR21), .ZN(_04373_) );
  AND2_X1 U18051 ( .A1(P2_rEIP_PTR24), .A2(P2_rEIP_PTR23), .ZN(_04374_) );
  AND2_X1 U18052 ( .A1(P2_rEIP_PTR26), .A2(P2_rEIP_PTR25), .ZN(_04375_) );
  AND2_X1 U18053 ( .A1(_04366_), .A2(_04365_), .ZN(_04378_) );
  AND2_X1 U18054 ( .A1(_04368_), .A2(_04367_), .ZN(_04379_) );
  AND2_X1 U18055 ( .A1(_04370_), .A2(_04369_), .ZN(_04380_) );
  AND2_X1 U18056 ( .A1(_04372_), .A2(_04371_), .ZN(_04381_) );
  AND2_X1 U18057 ( .A1(_04374_), .A2(_04373_), .ZN(_04382_) );
  AND2_X1 U18058 ( .A1(_04376_), .A2(_04375_), .ZN(_04383_) );
  AND2_X1 U18059 ( .A1(_04380_), .A2(_04379_), .ZN(_04384_) );
  AND2_X1 U18060 ( .A1(_04385_), .A2(_03066__PTR15), .ZN(_03066__PTR23) );
  AND2_X1 U18061 ( .A1(_04379_), .A2(_03066__PTR7), .ZN(_03066__PTR11) );
  AND2_X1 U18062 ( .A1(_04381_), .A2(_03066__PTR15), .ZN(_03066__PTR19) );
  AND2_X1 U18063 ( .A1(_04383_), .A2(_03066__PTR23), .ZN(_03066__PTR27) );
  AND2_X1 U18064 ( .A1(_04365_), .A2(_03066__PTR3), .ZN(_03066__PTR5) );
  AND2_X1 U18065 ( .A1(_04367_), .A2(_03066__PTR7), .ZN(_03066__PTR9) );
  AND2_X1 U18066 ( .A1(_04369_), .A2(_03066__PTR11), .ZN(_03066__PTR13) );
  AND2_X1 U18067 ( .A1(_04371_), .A2(_03066__PTR15), .ZN(_03066__PTR17) );
  AND2_X1 U18068 ( .A1(_04373_), .A2(_03066__PTR19), .ZN(_03066__PTR21) );
  AND2_X1 U18069 ( .A1(_04375_), .A2(_03066__PTR23), .ZN(_03066__PTR25) );
  AND2_X1 U18070 ( .A1(_04377_), .A2(_03066__PTR27), .ZN(_03066__PTR29) );
  AND2_X1 U18071 ( .A1(P2_rEIP_PTR3), .A2(_03066__PTR1), .ZN(_03066__PTR2) );
  AND2_X1 U18072 ( .A1(P2_rEIP_PTR5), .A2(_03066__PTR3), .ZN(_03066__PTR4) );
  AND2_X1 U18073 ( .A1(P2_rEIP_PTR7), .A2(_03066__PTR5), .ZN(_03066__PTR6) );
  AND2_X1 U18074 ( .A1(P2_rEIP_PTR9), .A2(_03066__PTR7), .ZN(_03066__PTR8) );
  AND2_X1 U18075 ( .A1(P2_rEIP_PTR11), .A2(_03066__PTR9), .ZN(_03066__PTR10) );
  AND2_X1 U18076 ( .A1(P2_rEIP_PTR13), .A2(_03066__PTR11), .ZN(_03066__PTR12) );
  AND2_X1 U18077 ( .A1(P2_rEIP_PTR15), .A2(_03066__PTR13), .ZN(_03066__PTR14) );
  AND2_X1 U18078 ( .A1(P2_rEIP_PTR17), .A2(_03066__PTR15), .ZN(_03066__PTR16) );
  AND2_X1 U18079 ( .A1(P2_rEIP_PTR19), .A2(_03066__PTR17), .ZN(_03066__PTR18) );
  AND2_X1 U18080 ( .A1(P2_rEIP_PTR21), .A2(_03066__PTR19), .ZN(_03066__PTR20) );
  AND2_X1 U18081 ( .A1(P2_rEIP_PTR23), .A2(_03066__PTR21), .ZN(_03066__PTR22) );
  AND2_X1 U18082 ( .A1(P2_rEIP_PTR25), .A2(_03066__PTR23), .ZN(_03066__PTR24) );
  AND2_X1 U18083 ( .A1(P2_rEIP_PTR27), .A2(_03066__PTR25), .ZN(_03066__PTR26) );
  AND2_X1 U18084 ( .A1(P2_rEIP_PTR29), .A2(_03066__PTR27), .ZN(_03066__PTR28) );
  AND2_X1 U18085 ( .A1(_02979__PTR1), .A2(_02389__PTR32), .ZN(_03192__PTR1) );
  AND2_X1 U18086 ( .A1(_04202_), .A2(_03192__PTR1), .ZN(_03192__PTR3) );
  AND2_X1 U18087 ( .A1(_04231_), .A2(_03192__PTR3), .ZN(_03192__PTR7) );
  AND2_X1 U18088 ( .A1(_04238_), .A2(_03192__PTR7), .ZN(_03192__PTR15) );
  AND2_X1 U18089 ( .A1(_02979__PTR5), .A2(_02979__PTR4), .ZN(_04217_) );
  AND2_X1 U18090 ( .A1(_02979__PTR15), .A2(_02979__PTR14), .ZN(_04222_) );
  AND2_X1 U18091 ( .A1(_02979__PTR17), .A2(_02979__PTR16), .ZN(_04223_) );
  AND2_X1 U18092 ( .A1(_02979__PTR21), .A2(_02979__PTR20), .ZN(_04225_) );
  AND2_X1 U18093 ( .A1(_04233_), .A2(_04232_), .ZN(_04238_) );
  AND2_X1 U18094 ( .A1(_04235_), .A2(_04234_), .ZN(_04239_) );
  AND2_X1 U18095 ( .A1(_04237_), .A2(_04236_), .ZN(_04240_) );
  AND2_X1 U18096 ( .A1(_04240_), .A2(_04239_), .ZN(_04241_) );
  AND2_X1 U18097 ( .A1(_04239_), .A2(_03192__PTR15), .ZN(_03192__PTR23) );
  AND2_X1 U18098 ( .A1(_04232_), .A2(_03192__PTR7), .ZN(_03192__PTR11) );
  AND2_X1 U18099 ( .A1(_04234_), .A2(_03192__PTR15), .ZN(_03192__PTR19) );
  AND2_X1 U18100 ( .A1(_04236_), .A2(_03192__PTR23), .ZN(_03192__PTR27) );
  AND2_X1 U18101 ( .A1(_04217_), .A2(_03192__PTR3), .ZN(_03192__PTR5) );
  AND2_X1 U18102 ( .A1(_04219_), .A2(_03192__PTR7), .ZN(_03192__PTR9) );
  AND2_X1 U18103 ( .A1(_04221_), .A2(_03192__PTR11), .ZN(_03192__PTR13) );
  AND2_X1 U18104 ( .A1(_04223_), .A2(_03192__PTR15), .ZN(_03192__PTR17) );
  AND2_X1 U18105 ( .A1(_04225_), .A2(_03192__PTR19), .ZN(_03192__PTR21) );
  AND2_X1 U18106 ( .A1(_04227_), .A2(_03192__PTR23), .ZN(_03192__PTR25) );
  AND2_X1 U18107 ( .A1(_04229_), .A2(_03192__PTR27), .ZN(_03192__PTR29) );
  AND2_X1 U18108 ( .A1(_02979__PTR2), .A2(_03192__PTR1), .ZN(_03192__PTR2) );
  AND2_X1 U18109 ( .A1(_02979__PTR4), .A2(_03192__PTR3), .ZN(_03192__PTR4) );
  AND2_X1 U18110 ( .A1(_02979__PTR6), .A2(_03192__PTR5), .ZN(_03192__PTR6) );
  AND2_X1 U18111 ( .A1(_02979__PTR8), .A2(_03192__PTR7), .ZN(_03192__PTR8) );
  AND2_X1 U18112 ( .A1(_02979__PTR10), .A2(_03192__PTR9), .ZN(_03192__PTR10) );
  AND2_X1 U18113 ( .A1(_02979__PTR12), .A2(_03192__PTR11), .ZN(_03192__PTR12) );
  AND2_X1 U18114 ( .A1(_02979__PTR14), .A2(_03192__PTR13), .ZN(_03192__PTR14) );
  AND2_X1 U18115 ( .A1(_02979__PTR16), .A2(_03192__PTR15), .ZN(_03192__PTR16) );
  AND2_X1 U18116 ( .A1(_02979__PTR18), .A2(_03192__PTR17), .ZN(_03192__PTR18) );
  AND2_X1 U18117 ( .A1(_02979__PTR20), .A2(_03192__PTR19), .ZN(_03192__PTR20) );
  AND2_X1 U18118 ( .A1(_02979__PTR22), .A2(_03192__PTR21), .ZN(_03192__PTR22) );
  AND2_X1 U18119 ( .A1(_02979__PTR24), .A2(_03192__PTR23), .ZN(_03192__PTR24) );
  AND2_X1 U18120 ( .A1(_02979__PTR26), .A2(_03192__PTR25), .ZN(_03192__PTR26) );
  AND2_X1 U18121 ( .A1(_02979__PTR28), .A2(_03192__PTR27), .ZN(_03192__PTR28) );
  AND2_X1 U18122 ( .A1(_02979__PTR30), .A2(_03192__PTR29), .ZN(_03192__PTR30) );
  AND2_X1 U18123 ( .A1(_02979__PTR3), .A2(P2_EBX_PTR2), .ZN(_04187_) );
  AND2_X1 U18124 ( .A1(_02979__PTR5), .A2(P2_EBX_PTR4), .ZN(_04188_) );
  AND2_X1 U18125 ( .A1(_02979__PTR7), .A2(P2_EBX_PTR6), .ZN(_04189_) );
  AND2_X1 U18126 ( .A1(_02979__PTR9), .A2(P2_EBX_PTR8), .ZN(_04190_) );
  AND2_X1 U18127 ( .A1(_02979__PTR11), .A2(P2_EBX_PTR10), .ZN(_04191_) );
  AND2_X1 U18128 ( .A1(_02979__PTR13), .A2(P2_EBX_PTR12), .ZN(_04192_) );
  AND2_X1 U18129 ( .A1(_02979__PTR15), .A2(P2_EBX_PTR14), .ZN(_04193_) );
  AND2_X1 U18130 ( .A1(_02979__PTR17), .A2(P2_EBX_PTR16), .ZN(_04194_) );
  AND2_X1 U18131 ( .A1(_02979__PTR19), .A2(P2_EBX_PTR18), .ZN(_04195_) );
  AND2_X1 U18132 ( .A1(_02979__PTR21), .A2(P2_EBX_PTR20), .ZN(_04196_) );
  AND2_X1 U18133 ( .A1(_02979__PTR23), .A2(P2_EBX_PTR22), .ZN(_04197_) );
  AND2_X1 U18134 ( .A1(_02979__PTR25), .A2(P2_EBX_PTR24), .ZN(_04198_) );
  AND2_X1 U18135 ( .A1(_02979__PTR27), .A2(P2_EBX_PTR26), .ZN(_04199_) );
  AND2_X1 U18136 ( .A1(_02979__PTR29), .A2(P2_EBX_PTR28), .ZN(_04200_) );
  AND2_X1 U18137 ( .A1(_02977__PTR31), .A2(P2_EBX_PTR30), .ZN(_04201_) );
  AND2_X1 U18138 ( .A1(_04218_), .A2(_04243_), .ZN(_04203_) );
  AND2_X1 U18139 ( .A1(_04220_), .A2(_04245_), .ZN(_04204_) );
  AND2_X1 U18140 ( .A1(_04222_), .A2(_04247_), .ZN(_04205_) );
  AND2_X1 U18141 ( .A1(_04224_), .A2(_04249_), .ZN(_04206_) );
  AND2_X1 U18142 ( .A1(_04226_), .A2(_04251_), .ZN(_04207_) );
  AND2_X1 U18143 ( .A1(_04228_), .A2(_04253_), .ZN(_04208_) );
  AND2_X1 U18144 ( .A1(_04230_), .A2(_04255_), .ZN(_04209_) );
  AND2_X1 U18145 ( .A1(_04231_), .A2(_02978__PTR3), .ZN(_04210_) );
  AND2_X1 U18146 ( .A1(_04233_), .A2(_04257_), .ZN(_04211_) );
  AND2_X1 U18147 ( .A1(_04235_), .A2(_04259_), .ZN(_04212_) );
  AND2_X1 U18148 ( .A1(_04237_), .A2(_04261_), .ZN(_04213_) );
  AND2_X1 U18149 ( .A1(_04238_), .A2(_02978__PTR7), .ZN(_04214_) );
  AND2_X1 U18150 ( .A1(_04240_), .A2(_04264_), .ZN(_04215_) );
  AND2_X1 U18151 ( .A1(_04241_), .A2(_02978__PTR15), .ZN(_04216_) );
  AND2_X1 U18152 ( .A1(_02979__PTR3), .A2(_02979__PTR2), .ZN(_04202_) );
  AND2_X1 U18153 ( .A1(_02979__PTR7), .A2(_02979__PTR6), .ZN(_04218_) );
  AND2_X1 U18154 ( .A1(_02979__PTR9), .A2(_02979__PTR8), .ZN(_04219_) );
  AND2_X1 U18155 ( .A1(_02979__PTR11), .A2(_02979__PTR10), .ZN(_04220_) );
  AND2_X1 U18156 ( .A1(_02979__PTR13), .A2(_02979__PTR12), .ZN(_04221_) );
  AND2_X1 U18157 ( .A1(_02979__PTR19), .A2(_02979__PTR18), .ZN(_04224_) );
  AND2_X1 U18158 ( .A1(_02979__PTR23), .A2(_02979__PTR22), .ZN(_04226_) );
  AND2_X1 U18159 ( .A1(_02979__PTR25), .A2(_02979__PTR24), .ZN(_04227_) );
  AND2_X1 U18160 ( .A1(_02979__PTR27), .A2(_02979__PTR26), .ZN(_04228_) );
  AND2_X1 U18161 ( .A1(_02979__PTR29), .A2(_02979__PTR28), .ZN(_04229_) );
  AND2_X1 U18162 ( .A1(_02977__PTR31), .A2(_02979__PTR30), .ZN(_04230_) );
  AND2_X1 U18163 ( .A1(_04218_), .A2(_04217_), .ZN(_04231_) );
  AND2_X1 U18164 ( .A1(_04220_), .A2(_04219_), .ZN(_04232_) );
  AND2_X1 U18165 ( .A1(_04222_), .A2(_04221_), .ZN(_04233_) );
  AND2_X1 U18166 ( .A1(_04224_), .A2(_04223_), .ZN(_04234_) );
  AND2_X1 U18167 ( .A1(_04226_), .A2(_04225_), .ZN(_04235_) );
  AND2_X1 U18168 ( .A1(_04228_), .A2(_04227_), .ZN(_04236_) );
  AND2_X1 U18169 ( .A1(_04230_), .A2(_04229_), .ZN(_04237_) );
  OR2_X1 U18170 ( .A1(P2_EBX_PTR3), .A2(_04187_), .ZN(_04242_) );
  OR2_X1 U18171 ( .A1(P2_EBX_PTR5), .A2(_04188_), .ZN(_04243_) );
  OR2_X1 U18172 ( .A1(P2_EBX_PTR7), .A2(_04189_), .ZN(_04244_) );
  OR2_X1 U18173 ( .A1(P2_EBX_PTR9), .A2(_04190_), .ZN(_04245_) );
  OR2_X1 U18174 ( .A1(P2_EBX_PTR11), .A2(_04191_), .ZN(_04246_) );
  OR2_X1 U18175 ( .A1(P2_EBX_PTR13), .A2(_04192_), .ZN(_04247_) );
  OR2_X1 U18176 ( .A1(P2_EBX_PTR15), .A2(_04193_), .ZN(_04248_) );
  OR2_X1 U18177 ( .A1(P2_EBX_PTR17), .A2(_04194_), .ZN(_04249_) );
  OR2_X1 U18178 ( .A1(P2_EBX_PTR19), .A2(_04195_), .ZN(_04250_) );
  OR2_X1 U18179 ( .A1(P2_EBX_PTR21), .A2(_04196_), .ZN(_04251_) );
  OR2_X1 U18180 ( .A1(P2_EBX_PTR23), .A2(_04197_), .ZN(_04252_) );
  OR2_X1 U18181 ( .A1(P2_EBX_PTR25), .A2(_04198_), .ZN(_04253_) );
  OR2_X1 U18182 ( .A1(P2_EBX_PTR27), .A2(_04199_), .ZN(_04254_) );
  OR2_X1 U18183 ( .A1(P2_EBX_PTR29), .A2(_04200_), .ZN(_04255_) );
  OR2_X1 U18184 ( .A1(_04242_), .A2(_04202_), .ZN(_02978__PTR3) );
  OR2_X1 U18185 ( .A1(_04244_), .A2(_04203_), .ZN(_04256_) );
  OR2_X1 U18186 ( .A1(_04246_), .A2(_04204_), .ZN(_04257_) );
  OR2_X1 U18187 ( .A1(_04248_), .A2(_04205_), .ZN(_04258_) );
  OR2_X1 U18188 ( .A1(_04250_), .A2(_04206_), .ZN(_04259_) );
  OR2_X1 U18189 ( .A1(_04252_), .A2(_04207_), .ZN(_04260_) );
  OR2_X1 U18190 ( .A1(_04254_), .A2(_04208_), .ZN(_04261_) );
  OR2_X1 U18191 ( .A1(_04201_), .A2(_04209_), .ZN(_04262_) );
  OR2_X1 U18192 ( .A1(_04256_), .A2(_04210_), .ZN(_02978__PTR7) );
  OR2_X1 U18193 ( .A1(_04258_), .A2(_04211_), .ZN(_04263_) );
  OR2_X1 U18194 ( .A1(_04260_), .A2(_04212_), .ZN(_04264_) );
  OR2_X1 U18195 ( .A1(_04262_), .A2(_04213_), .ZN(_04265_) );
  OR2_X1 U18196 ( .A1(_04263_), .A2(_04214_), .ZN(_02978__PTR15) );
  OR2_X1 U18197 ( .A1(_04265_), .A2(_04215_), .ZN(_04266_) );
  OR2_X1 U18198 ( .A1(_04266_), .A2(_04216_), .ZN(_02978__PTR31) );
  AND2_X1 U18199 ( .A1(_03177__PTR1), .A2(_03176__PTR0), .ZN(_04625_) );
  AND2_X1 U18200 ( .A1(_03177__PTR3), .A2(_03178__PTR2), .ZN(_04626_) );
  AND2_X1 U18201 ( .A1(_04628_), .A2(_03176__PTR1), .ZN(_04627_) );
  AND2_X1 U18202 ( .A1(_03177__PTR3), .A2(_03177__PTR2), .ZN(_04628_) );
  AND2_X1 U18203 ( .A1(_03177__PTR4), .A2(_03176__PTR3), .ZN(_04629_) );
  AND2_X1 U18204 ( .A1(_03177__PTR2), .A2(_03176__PTR1), .ZN(_04630_) );
  OR2_X1 U18205 ( .A1(_03178__PTR0), .A2(_02963__PTR0), .ZN(_03176__PTR0) );
  OR2_X1 U18206 ( .A1(_03178__PTR1), .A2(_04625_), .ZN(_03176__PTR1) );
  OR2_X1 U18207 ( .A1(_03178__PTR3), .A2(_04626_), .ZN(_04631_) );
  OR2_X1 U18208 ( .A1(_04631_), .A2(_04627_), .ZN(_03176__PTR3) );
  OR2_X1 U18209 ( .A1(_03178__PTR4), .A2(_04629_), .ZN(_02965__PTR5) );
  OR2_X1 U18210 ( .A1(_03178__PTR2), .A2(_04630_), .ZN(_03176__PTR2) );
  AND2_X1 U18211 ( .A1(_02962__PTR1), .A2(_02963__PTR0), .ZN(_00942__PTR0) );
  AND2_X1 U18212 ( .A1(_02964__PTR3), .A2(_02974__PTR1), .ZN(_02974__PTR3) );
  AND2_X1 U18213 ( .A1(_02965__PTR5), .A2(_02963__PTR4), .ZN(_00942__PTR2) );
  AND2_X1 U18214 ( .A1(_00942__PTR2), .A2(_02974__PTR3), .ZN(_04186_) );
  OR2_X1 U18215 ( .A1(_02963__PTR1), .A2(_00942__PTR0), .ZN(_02974__PTR1) );
  OR2_X1 U18216 ( .A1(_02961__PTR5), .A2(_04186_), .ZN(_02974__PTR5) );
  AND2_X1 U18217 ( .A1(P2_P1_InstQueueRd_Addr_PTR1), .A2(P2_P1_InstQueueRd_Addr_PTR0), .ZN(_02995__PTR1) );
  AND2_X1 U18218 ( .A1(_02178__PTR5), .A2(_02995__PTR1), .ZN(_04580_) );
  OR2_X1 U18219 ( .A1(P2_P1_InstQueueRd_Addr_PTR2), .A2(_04580_), .ZN(_03064__PTR2) );
  AND2_X1 U18220 ( .A1(P2_P1_InstQueueRd_Addr_PTR2), .A2(P2_P1_InstQueueRd_Addr_PTR1), .ZN(_03062__PTR1) );
  AND2_X1 U18221 ( .A1(P2_P1_InstQueueRd_Addr_PTR3), .A2(_03062__PTR1), .ZN(_03062__PTR2) );
  AND2_X1 U18222 ( .A1(_02179__PTR1), .A2(_03059__PTR0), .ZN(_03059__PTR1) );
  AND2_X1 U18223 ( .A1(_04576_), .A2(_03059__PTR1), .ZN(_03059__PTR3) );
  AND2_X1 U18224 ( .A1(_04579_), .A2(_03059__PTR3), .ZN(_03059__PTR7) );
  AND2_X1 U18225 ( .A1(_02179__PTR3), .A2(_02179__PTR2), .ZN(_04576_) );
  AND2_X1 U18226 ( .A1(_02179__PTR5), .A2(_02179__PTR4), .ZN(_04577_) );
  AND2_X1 U18227 ( .A1(_02179__PTR7), .A2(_02179__PTR6), .ZN(_04578_) );
  AND2_X1 U18228 ( .A1(_04578_), .A2(_04577_), .ZN(_04579_) );
  AND2_X1 U18229 ( .A1(_04577_), .A2(_03059__PTR3), .ZN(_03059__PTR5) );
  AND2_X1 U18230 ( .A1(_02179__PTR2), .A2(_03059__PTR1), .ZN(_03059__PTR2) );
  AND2_X1 U18231 ( .A1(_02179__PTR4), .A2(_03059__PTR3), .ZN(_03059__PTR4) );
  AND2_X1 U18232 ( .A1(_02179__PTR6), .A2(_03059__PTR5), .ZN(_03059__PTR6) );
  AND2_X1 U18233 ( .A1(_02182__PTR4), .A2(P2_P1_InstQueueRd_Addr_PTR0), .ZN(_04575_) );
  AND2_X1 U18234 ( .A1(P2_P1_InstQueueRd_Addr_PTR2), .A2(_03058__PTR1), .ZN(_03058__PTR2) );
  OR2_X1 U18235 ( .A1(P2_P1_InstQueueRd_Addr_PTR1), .A2(_04575_), .ZN(_03058__PTR1) );
  AND2_X1 U18236 ( .A1(P2_P1_InstAddrPointer_PTR3), .A2(P2_P1_InstAddrPointer_PTR2), .ZN(_04454_) );
  AND2_X1 U18237 ( .A1(_04536_), .A2(_03043__PTR1), .ZN(_04535_) );
  AND2_X1 U18238 ( .A1(_04468_), .A2(_03051__PTR3), .ZN(_03051__PTR7) );
  AND2_X1 U18239 ( .A1(_04474_), .A2(_03051__PTR7), .ZN(_03051__PTR15) );
  AND2_X1 U18240 ( .A1(P2_P1_InstAddrPointer_PTR3), .A2(_02990__PTR2), .ZN(_04536_) );
  AND2_X1 U18241 ( .A1(P2_P1_InstAddrPointer_PTR5), .A2(P2_P1_InstAddrPointer_PTR4), .ZN(_04455_) );
  AND2_X1 U18242 ( .A1(P2_P1_InstAddrPointer_PTR7), .A2(P2_P1_InstAddrPointer_PTR6), .ZN(_04456_) );
  AND2_X1 U18243 ( .A1(P2_P1_InstAddrPointer_PTR9), .A2(P2_P1_InstAddrPointer_PTR8), .ZN(_04457_) );
  AND2_X1 U18244 ( .A1(P2_P1_InstAddrPointer_PTR11), .A2(P2_P1_InstAddrPointer_PTR10), .ZN(_04458_) );
  AND2_X1 U18245 ( .A1(P2_P1_InstAddrPointer_PTR13), .A2(P2_P1_InstAddrPointer_PTR12), .ZN(_04459_) );
  AND2_X1 U18246 ( .A1(P2_P1_InstAddrPointer_PTR15), .A2(P2_P1_InstAddrPointer_PTR14), .ZN(_04460_) );
  AND2_X1 U18247 ( .A1(P2_P1_InstAddrPointer_PTR19), .A2(P2_P1_InstAddrPointer_PTR18), .ZN(_04462_) );
  AND2_X1 U18248 ( .A1(P2_P1_InstAddrPointer_PTR21), .A2(P2_P1_InstAddrPointer_PTR20), .ZN(_04463_) );
  AND2_X1 U18249 ( .A1(P2_P1_InstAddrPointer_PTR23), .A2(P2_P1_InstAddrPointer_PTR22), .ZN(_04464_) );
  AND2_X1 U18250 ( .A1(P2_P1_InstAddrPointer_PTR25), .A2(P2_P1_InstAddrPointer_PTR24), .ZN(_04465_) );
  AND2_X1 U18251 ( .A1(P2_P1_InstAddrPointer_PTR27), .A2(P2_P1_InstAddrPointer_PTR26), .ZN(_04466_) );
  AND2_X1 U18252 ( .A1(P2_P1_InstAddrPointer_PTR29), .A2(P2_P1_InstAddrPointer_PTR28), .ZN(_04467_) );
  AND2_X1 U18253 ( .A1(_04456_), .A2(_04455_), .ZN(_04468_) );
  AND2_X1 U18254 ( .A1(_04458_), .A2(_04457_), .ZN(_04469_) );
  AND2_X1 U18255 ( .A1(_04460_), .A2(_04459_), .ZN(_04470_) );
  AND2_X1 U18256 ( .A1(_04462_), .A2(_04461_), .ZN(_04471_) );
  AND2_X1 U18257 ( .A1(_04466_), .A2(_04465_), .ZN(_04473_) );
  AND2_X1 U18258 ( .A1(_04472_), .A2(_04471_), .ZN(_04475_) );
  AND2_X1 U18259 ( .A1(_04475_), .A2(_03051__PTR15), .ZN(_03051__PTR23) );
  AND2_X1 U18260 ( .A1(_04469_), .A2(_03051__PTR7), .ZN(_03051__PTR11) );
  AND2_X1 U18261 ( .A1(_04471_), .A2(_03051__PTR15), .ZN(_03051__PTR19) );
  AND2_X1 U18262 ( .A1(_04473_), .A2(_03051__PTR23), .ZN(_03051__PTR27) );
  AND2_X1 U18263 ( .A1(_04455_), .A2(_03051__PTR3), .ZN(_03051__PTR5) );
  AND2_X1 U18264 ( .A1(_04457_), .A2(_03051__PTR7), .ZN(_03051__PTR9) );
  AND2_X1 U18265 ( .A1(_04459_), .A2(_03051__PTR11), .ZN(_03051__PTR13) );
  AND2_X1 U18266 ( .A1(_04461_), .A2(_03051__PTR15), .ZN(_03051__PTR17) );
  AND2_X1 U18267 ( .A1(_04463_), .A2(_03051__PTR19), .ZN(_03051__PTR21) );
  AND2_X1 U18268 ( .A1(_04465_), .A2(_03051__PTR23), .ZN(_03051__PTR25) );
  AND2_X1 U18269 ( .A1(_04467_), .A2(_03051__PTR27), .ZN(_03051__PTR29) );
  AND2_X1 U18270 ( .A1(_02990__PTR2), .A2(_03043__PTR1), .ZN(_04537_) );
  AND2_X1 U18271 ( .A1(P2_P1_InstAddrPointer_PTR4), .A2(_03051__PTR3), .ZN(_03051__PTR4) );
  AND2_X1 U18272 ( .A1(P2_P1_InstAddrPointer_PTR6), .A2(_03051__PTR5), .ZN(_03051__PTR6) );
  AND2_X1 U18273 ( .A1(P2_P1_InstAddrPointer_PTR8), .A2(_03051__PTR7), .ZN(_03051__PTR8) );
  AND2_X1 U18274 ( .A1(P2_P1_InstAddrPointer_PTR10), .A2(_03051__PTR9), .ZN(_03051__PTR10) );
  AND2_X1 U18275 ( .A1(P2_P1_InstAddrPointer_PTR12), .A2(_03051__PTR11), .ZN(_03051__PTR12) );
  AND2_X1 U18276 ( .A1(P2_P1_InstAddrPointer_PTR14), .A2(_03051__PTR13), .ZN(_03051__PTR14) );
  AND2_X1 U18277 ( .A1(P2_P1_InstAddrPointer_PTR16), .A2(_03051__PTR15), .ZN(_03051__PTR16) );
  AND2_X1 U18278 ( .A1(P2_P1_InstAddrPointer_PTR18), .A2(_03051__PTR17), .ZN(_03051__PTR18) );
  AND2_X1 U18279 ( .A1(P2_P1_InstAddrPointer_PTR20), .A2(_03051__PTR19), .ZN(_03051__PTR20) );
  AND2_X1 U18280 ( .A1(P2_P1_InstAddrPointer_PTR22), .A2(_03051__PTR21), .ZN(_03051__PTR22) );
  AND2_X1 U18281 ( .A1(P2_P1_InstAddrPointer_PTR24), .A2(_03051__PTR23), .ZN(_03051__PTR24) );
  AND2_X1 U18282 ( .A1(P2_P1_InstAddrPointer_PTR26), .A2(_03051__PTR25), .ZN(_03051__PTR26) );
  AND2_X1 U18283 ( .A1(P2_P1_InstAddrPointer_PTR28), .A2(_03051__PTR27), .ZN(_03051__PTR28) );
  AND2_X1 U18284 ( .A1(P2_P1_InstAddrPointer_PTR30), .A2(_03051__PTR29), .ZN(_03051__PTR30) );
  OR2_X1 U18285 ( .A1(_04454_), .A2(_04535_), .ZN(_03051__PTR3) );
  OR2_X1 U18286 ( .A1(P2_P1_InstAddrPointer_PTR2), .A2(_04537_), .ZN(_03051__PTR2) );
  AND2_X1 U18287 ( .A1(_03054__PTR1), .A2(_03053__PTR0), .ZN(_04538_) );
  AND2_X1 U18288 ( .A1(_03054__PTR3), .A2(_03056__PTR2), .ZN(_04539_) );
  AND2_X1 U18289 ( .A1(_03054__PTR5), .A2(_03056__PTR4), .ZN(_04540_) );
  AND2_X1 U18290 ( .A1(_03054__PTR7), .A2(_03056__PTR6), .ZN(_04541_) );
  AND2_X1 U18291 ( .A1(_04545_), .A2(_03053__PTR1), .ZN(_04542_) );
  AND2_X1 U18292 ( .A1(_04547_), .A2(_04572_), .ZN(_04543_) );
  AND2_X1 U18293 ( .A1(_04559_), .A2(_03053__PTR3), .ZN(_04544_) );
  AND2_X1 U18294 ( .A1(_04565_), .A2(_03053__PTR7), .ZN(_03053__PTR15) );
  AND2_X1 U18295 ( .A1(_03054__PTR3), .A2(_03054__PTR2), .ZN(_04545_) );
  AND2_X1 U18296 ( .A1(_03054__PTR5), .A2(_03054__PTR4), .ZN(_04546_) );
  AND2_X1 U18297 ( .A1(_03054__PTR7), .A2(_03054__PTR6), .ZN(_04547_) );
  AND2_X1 U18298 ( .A1(_03052__PTR9), .A2(_03052__PTR8), .ZN(_04548_) );
  AND2_X1 U18299 ( .A1(_03052__PTR11), .A2(_03052__PTR10), .ZN(_04549_) );
  AND2_X1 U18300 ( .A1(_03052__PTR13), .A2(_03052__PTR12), .ZN(_04550_) );
  AND2_X1 U18301 ( .A1(_03052__PTR15), .A2(_03052__PTR14), .ZN(_04551_) );
  AND2_X1 U18302 ( .A1(_03052__PTR17), .A2(_03052__PTR16), .ZN(_04552_) );
  AND2_X1 U18303 ( .A1(_03052__PTR19), .A2(_03052__PTR18), .ZN(_04553_) );
  AND2_X1 U18304 ( .A1(_03052__PTR21), .A2(_03052__PTR20), .ZN(_04554_) );
  AND2_X1 U18305 ( .A1(_03052__PTR23), .A2(_03052__PTR22), .ZN(_04555_) );
  AND2_X1 U18306 ( .A1(_03052__PTR25), .A2(_03052__PTR24), .ZN(_04556_) );
  AND2_X1 U18307 ( .A1(_03052__PTR27), .A2(_03052__PTR26), .ZN(_04557_) );
  AND2_X1 U18308 ( .A1(_03052__PTR29), .A2(_03052__PTR28), .ZN(_04558_) );
  AND2_X1 U18309 ( .A1(_04547_), .A2(_04546_), .ZN(_04559_) );
  AND2_X1 U18310 ( .A1(_04549_), .A2(_04548_), .ZN(_04560_) );
  AND2_X1 U18311 ( .A1(_04551_), .A2(_04550_), .ZN(_04561_) );
  AND2_X1 U18312 ( .A1(_04553_), .A2(_04552_), .ZN(_04562_) );
  AND2_X1 U18313 ( .A1(_04555_), .A2(_04554_), .ZN(_04563_) );
  AND2_X1 U18314 ( .A1(_04557_), .A2(_04556_), .ZN(_04564_) );
  AND2_X1 U18315 ( .A1(_04561_), .A2(_04560_), .ZN(_04565_) );
  AND2_X1 U18316 ( .A1(_04563_), .A2(_04562_), .ZN(_04566_) );
  AND2_X1 U18317 ( .A1(_04566_), .A2(_03053__PTR15), .ZN(_03053__PTR23) );
  AND2_X1 U18318 ( .A1(_04560_), .A2(_03053__PTR7), .ZN(_03053__PTR11) );
  AND2_X1 U18319 ( .A1(_04562_), .A2(_03053__PTR15), .ZN(_03053__PTR19) );
  AND2_X1 U18320 ( .A1(_04564_), .A2(_03053__PTR23), .ZN(_03053__PTR27) );
  AND2_X1 U18321 ( .A1(_04546_), .A2(_03053__PTR3), .ZN(_04567_) );
  AND2_X1 U18322 ( .A1(_04548_), .A2(_03053__PTR7), .ZN(_03053__PTR9) );
  AND2_X1 U18323 ( .A1(_04550_), .A2(_03053__PTR11), .ZN(_03053__PTR13) );
  AND2_X1 U18324 ( .A1(_04552_), .A2(_03053__PTR15), .ZN(_03053__PTR17) );
  AND2_X1 U18325 ( .A1(_04554_), .A2(_03053__PTR19), .ZN(_03053__PTR21) );
  AND2_X1 U18326 ( .A1(_04556_), .A2(_03053__PTR23), .ZN(_03053__PTR25) );
  AND2_X1 U18327 ( .A1(_04558_), .A2(_03053__PTR27), .ZN(_03053__PTR29) );
  AND2_X1 U18328 ( .A1(_03054__PTR2), .A2(_03053__PTR1), .ZN(_04568_) );
  AND2_X1 U18329 ( .A1(_03054__PTR4), .A2(_03053__PTR3), .ZN(_04569_) );
  AND2_X1 U18330 ( .A1(_03054__PTR6), .A2(_03053__PTR5), .ZN(_04570_) );
  AND2_X1 U18331 ( .A1(_03052__PTR8), .A2(_03053__PTR7), .ZN(_03053__PTR8) );
  AND2_X1 U18332 ( .A1(_03052__PTR10), .A2(_03053__PTR9), .ZN(_03053__PTR10) );
  AND2_X1 U18333 ( .A1(_03052__PTR12), .A2(_03053__PTR11), .ZN(_03053__PTR12) );
  AND2_X1 U18334 ( .A1(_03052__PTR14), .A2(_03053__PTR13), .ZN(_03053__PTR14) );
  AND2_X1 U18335 ( .A1(_03052__PTR16), .A2(_03053__PTR15), .ZN(_03053__PTR16) );
  AND2_X1 U18336 ( .A1(_03052__PTR18), .A2(_03053__PTR17), .ZN(_03053__PTR18) );
  AND2_X1 U18337 ( .A1(_03052__PTR20), .A2(_03053__PTR19), .ZN(_03053__PTR20) );
  AND2_X1 U18338 ( .A1(_03052__PTR22), .A2(_03053__PTR21), .ZN(_03053__PTR22) );
  AND2_X1 U18339 ( .A1(_03052__PTR24), .A2(_03053__PTR23), .ZN(_03053__PTR24) );
  AND2_X1 U18340 ( .A1(_03052__PTR26), .A2(_03053__PTR25), .ZN(_03053__PTR26) );
  AND2_X1 U18341 ( .A1(_03052__PTR28), .A2(_03053__PTR27), .ZN(_03053__PTR28) );
  AND2_X1 U18342 ( .A1(_03052__PTR30), .A2(_03053__PTR29), .ZN(_03053__PTR30) );
  OR2_X1 U18343 ( .A1(_03056__PTR1), .A2(_04538_), .ZN(_03053__PTR1) );
  OR2_X1 U18344 ( .A1(_03056__PTR3), .A2(_04539_), .ZN(_04571_) );
  OR2_X1 U18345 ( .A1(_03056__PTR5), .A2(_04540_), .ZN(_04572_) );
  OR2_X1 U18346 ( .A1(_03056__PTR7), .A2(_04541_), .ZN(_04573_) );
  OR2_X1 U18347 ( .A1(_04571_), .A2(_04542_), .ZN(_03053__PTR3) );
  OR2_X1 U18348 ( .A1(_04573_), .A2(_04543_), .ZN(_04574_) );
  OR2_X1 U18349 ( .A1(_04574_), .A2(_04544_), .ZN(_03053__PTR7) );
  OR2_X1 U18350 ( .A1(_04572_), .A2(_04567_), .ZN(_03053__PTR5) );
  OR2_X1 U18351 ( .A1(_03056__PTR2), .A2(_04568_), .ZN(_03053__PTR2) );
  OR2_X1 U18352 ( .A1(_03056__PTR4), .A2(_04569_), .ZN(_03053__PTR4) );
  OR2_X1 U18353 ( .A1(_03056__PTR6), .A2(_04570_), .ZN(_03053__PTR6) );
  AND2_X1 U18354 ( .A1(_00944__PTR1), .A2(_02963__PTR1), .ZN(_04184_) );
  AND2_X1 U18355 ( .A1(_02963__PTR3), .A2(_02962__PTR2), .ZN(_00944__PTR1) );
  AND2_X1 U18356 ( .A1(_00942__PTR2), .A2(_02971__PTR3), .ZN(_04185_) );
  OR2_X1 U18357 ( .A1(_02964__PTR3), .A2(_04184_), .ZN(_02971__PTR3) );
  OR2_X1 U18358 ( .A1(_02961__PTR5), .A2(_04185_), .ZN(_02971__PTR5) );
  AND2_X1 U18359 ( .A1(P2_P1_InstAddrPointer_PTR2), .A2(P2_P1_InstAddrPointer_PTR1), .ZN(_03046__PTR1) );
  AND2_X1 U18360 ( .A1(_04476_), .A2(_03046__PTR1), .ZN(_03046__PTR3) );
  AND2_X1 U18361 ( .A1(_04490_), .A2(_03046__PTR3), .ZN(_03046__PTR7) );
  AND2_X1 U18362 ( .A1(_04496_), .A2(_03046__PTR7), .ZN(_03046__PTR15) );
  AND2_X1 U18363 ( .A1(P2_P1_InstAddrPointer_PTR4), .A2(P2_P1_InstAddrPointer_PTR3), .ZN(_04476_) );
  AND2_X1 U18364 ( .A1(P2_P1_InstAddrPointer_PTR6), .A2(P2_P1_InstAddrPointer_PTR5), .ZN(_04477_) );
  AND2_X1 U18365 ( .A1(P2_P1_InstAddrPointer_PTR8), .A2(P2_P1_InstAddrPointer_PTR7), .ZN(_04478_) );
  AND2_X1 U18366 ( .A1(P2_P1_InstAddrPointer_PTR10), .A2(P2_P1_InstAddrPointer_PTR9), .ZN(_04479_) );
  AND2_X1 U18367 ( .A1(P2_P1_InstAddrPointer_PTR12), .A2(P2_P1_InstAddrPointer_PTR11), .ZN(_04480_) );
  AND2_X1 U18368 ( .A1(P2_P1_InstAddrPointer_PTR14), .A2(P2_P1_InstAddrPointer_PTR13), .ZN(_04481_) );
  AND2_X1 U18369 ( .A1(P2_P1_InstAddrPointer_PTR16), .A2(P2_P1_InstAddrPointer_PTR15), .ZN(_04482_) );
  AND2_X1 U18370 ( .A1(P2_P1_InstAddrPointer_PTR18), .A2(P2_P1_InstAddrPointer_PTR17), .ZN(_04483_) );
  AND2_X1 U18371 ( .A1(P2_P1_InstAddrPointer_PTR20), .A2(P2_P1_InstAddrPointer_PTR19), .ZN(_04484_) );
  AND2_X1 U18372 ( .A1(P2_P1_InstAddrPointer_PTR22), .A2(P2_P1_InstAddrPointer_PTR21), .ZN(_04485_) );
  AND2_X1 U18373 ( .A1(P2_P1_InstAddrPointer_PTR24), .A2(P2_P1_InstAddrPointer_PTR23), .ZN(_04486_) );
  AND2_X1 U18374 ( .A1(P2_P1_InstAddrPointer_PTR26), .A2(P2_P1_InstAddrPointer_PTR25), .ZN(_04487_) );
  AND2_X1 U18375 ( .A1(P2_P1_InstAddrPointer_PTR28), .A2(P2_P1_InstAddrPointer_PTR27), .ZN(_04488_) );
  AND2_X1 U18376 ( .A1(P2_P1_InstAddrPointer_PTR30), .A2(P2_P1_InstAddrPointer_PTR29), .ZN(_04489_) );
  AND2_X1 U18377 ( .A1(_04478_), .A2(_04477_), .ZN(_04490_) );
  AND2_X1 U18378 ( .A1(_04480_), .A2(_04479_), .ZN(_04491_) );
  AND2_X1 U18379 ( .A1(_04482_), .A2(_04481_), .ZN(_04492_) );
  AND2_X1 U18380 ( .A1(_04484_), .A2(_04483_), .ZN(_04493_) );
  AND2_X1 U18381 ( .A1(_04486_), .A2(_04485_), .ZN(_04494_) );
  AND2_X1 U18382 ( .A1(_04488_), .A2(_04487_), .ZN(_04495_) );
  AND2_X1 U18383 ( .A1(_04492_), .A2(_04491_), .ZN(_04496_) );
  AND2_X1 U18384 ( .A1(_04494_), .A2(_04493_), .ZN(_04497_) );
  AND2_X1 U18385 ( .A1(_04497_), .A2(_03046__PTR15), .ZN(_03046__PTR23) );
  AND2_X1 U18386 ( .A1(_04491_), .A2(_03046__PTR7), .ZN(_03046__PTR11) );
  AND2_X1 U18387 ( .A1(_04493_), .A2(_03046__PTR15), .ZN(_03046__PTR19) );
  AND2_X1 U18388 ( .A1(_04495_), .A2(_03046__PTR23), .ZN(_03046__PTR27) );
  AND2_X1 U18389 ( .A1(_04477_), .A2(_03046__PTR3), .ZN(_03046__PTR5) );
  AND2_X1 U18390 ( .A1(_04479_), .A2(_03046__PTR7), .ZN(_03046__PTR9) );
  AND2_X1 U18391 ( .A1(_04481_), .A2(_03046__PTR11), .ZN(_03046__PTR13) );
  AND2_X1 U18392 ( .A1(_04483_), .A2(_03046__PTR15), .ZN(_03046__PTR17) );
  AND2_X1 U18393 ( .A1(_04485_), .A2(_03046__PTR19), .ZN(_03046__PTR21) );
  AND2_X1 U18394 ( .A1(_04487_), .A2(_03046__PTR23), .ZN(_03046__PTR25) );
  AND2_X1 U18395 ( .A1(_04489_), .A2(_03046__PTR27), .ZN(_03046__PTR29) );
  AND2_X1 U18396 ( .A1(P2_P1_InstAddrPointer_PTR3), .A2(_03046__PTR1), .ZN(_03046__PTR2) );
  AND2_X1 U18397 ( .A1(P2_P1_InstAddrPointer_PTR5), .A2(_03046__PTR3), .ZN(_03046__PTR4) );
  AND2_X1 U18398 ( .A1(P2_P1_InstAddrPointer_PTR7), .A2(_03046__PTR5), .ZN(_03046__PTR6) );
  AND2_X1 U18399 ( .A1(P2_P1_InstAddrPointer_PTR9), .A2(_03046__PTR7), .ZN(_03046__PTR8) );
  AND2_X1 U18400 ( .A1(P2_P1_InstAddrPointer_PTR11), .A2(_03046__PTR9), .ZN(_03046__PTR10) );
  AND2_X1 U18401 ( .A1(P2_P1_InstAddrPointer_PTR13), .A2(_03046__PTR11), .ZN(_03046__PTR12) );
  AND2_X1 U18402 ( .A1(P2_P1_InstAddrPointer_PTR15), .A2(_03046__PTR13), .ZN(_03046__PTR14) );
  AND2_X1 U18403 ( .A1(P2_P1_InstAddrPointer_PTR17), .A2(_03046__PTR15), .ZN(_03046__PTR16) );
  AND2_X1 U18404 ( .A1(P2_P1_InstAddrPointer_PTR19), .A2(_03046__PTR17), .ZN(_03046__PTR18) );
  AND2_X1 U18405 ( .A1(P2_P1_InstAddrPointer_PTR21), .A2(_03046__PTR19), .ZN(_03046__PTR20) );
  AND2_X1 U18406 ( .A1(P2_P1_InstAddrPointer_PTR23), .A2(_03046__PTR21), .ZN(_03046__PTR22) );
  AND2_X1 U18407 ( .A1(P2_P1_InstAddrPointer_PTR25), .A2(_03046__PTR23), .ZN(_03046__PTR24) );
  AND2_X1 U18408 ( .A1(P2_P1_InstAddrPointer_PTR27), .A2(_03046__PTR25), .ZN(_03046__PTR26) );
  AND2_X1 U18409 ( .A1(P2_P1_InstAddrPointer_PTR29), .A2(_03046__PTR27), .ZN(_03046__PTR28) );
  AND2_X1 U18410 ( .A1(_03048__PTR1), .A2(_03047__PTR0), .ZN(_04498_) );
  AND2_X1 U18411 ( .A1(_03048__PTR3), .A2(_03050__PTR2), .ZN(_04499_) );
  AND2_X1 U18412 ( .A1(_03048__PTR5), .A2(_03050__PTR4), .ZN(_04500_) );
  AND2_X1 U18413 ( .A1(_03048__PTR7), .A2(_03050__PTR6), .ZN(_04501_) );
  AND2_X1 U18414 ( .A1(_04505_), .A2(_03047__PTR1), .ZN(_04502_) );
  AND2_X1 U18415 ( .A1(_04507_), .A2(_04532_), .ZN(_04503_) );
  AND2_X1 U18416 ( .A1(_04519_), .A2(_03047__PTR3), .ZN(_04504_) );
  AND2_X1 U18417 ( .A1(_04525_), .A2(_03047__PTR7), .ZN(_03047__PTR15) );
  AND2_X1 U18418 ( .A1(_03048__PTR3), .A2(_03048__PTR2), .ZN(_04505_) );
  AND2_X1 U18419 ( .A1(_03048__PTR5), .A2(_03048__PTR4), .ZN(_04506_) );
  AND2_X1 U18420 ( .A1(_03048__PTR7), .A2(_03048__PTR6), .ZN(_04507_) );
  AND2_X1 U18421 ( .A1(_02373__PTR41), .A2(_02373__PTR40), .ZN(_04508_) );
  AND2_X1 U18422 ( .A1(_02373__PTR43), .A2(_02373__PTR42), .ZN(_04509_) );
  AND2_X1 U18423 ( .A1(_02373__PTR45), .A2(_02373__PTR44), .ZN(_04510_) );
  AND2_X1 U18424 ( .A1(_02373__PTR47), .A2(_02373__PTR46), .ZN(_04511_) );
  AND2_X1 U18425 ( .A1(_02373__PTR49), .A2(_02373__PTR48), .ZN(_04512_) );
  AND2_X1 U18426 ( .A1(_02373__PTR51), .A2(_02373__PTR50), .ZN(_04513_) );
  AND2_X1 U18427 ( .A1(_02373__PTR53), .A2(_02373__PTR52), .ZN(_04514_) );
  AND2_X1 U18428 ( .A1(_02373__PTR55), .A2(_02373__PTR54), .ZN(_04515_) );
  AND2_X1 U18429 ( .A1(_02373__PTR57), .A2(_02373__PTR56), .ZN(_04516_) );
  AND2_X1 U18430 ( .A1(_02373__PTR59), .A2(_02373__PTR58), .ZN(_04517_) );
  AND2_X1 U18431 ( .A1(_02373__PTR61), .A2(_02373__PTR60), .ZN(_04518_) );
  AND2_X1 U18432 ( .A1(_04507_), .A2(_04506_), .ZN(_04519_) );
  AND2_X1 U18433 ( .A1(_04509_), .A2(_04508_), .ZN(_04520_) );
  AND2_X1 U18434 ( .A1(_04511_), .A2(_04510_), .ZN(_04521_) );
  AND2_X1 U18435 ( .A1(_04513_), .A2(_04512_), .ZN(_04522_) );
  AND2_X1 U18436 ( .A1(_04515_), .A2(_04514_), .ZN(_04523_) );
  AND2_X1 U18437 ( .A1(_04517_), .A2(_04516_), .ZN(_04524_) );
  AND2_X1 U18438 ( .A1(_04521_), .A2(_04520_), .ZN(_04525_) );
  AND2_X1 U18439 ( .A1(_04523_), .A2(_04522_), .ZN(_04526_) );
  AND2_X1 U18440 ( .A1(_04526_), .A2(_03047__PTR15), .ZN(_03047__PTR23) );
  AND2_X1 U18441 ( .A1(_04520_), .A2(_03047__PTR7), .ZN(_03047__PTR11) );
  AND2_X1 U18442 ( .A1(_04522_), .A2(_03047__PTR15), .ZN(_03047__PTR19) );
  AND2_X1 U18443 ( .A1(_04524_), .A2(_03047__PTR23), .ZN(_03047__PTR27) );
  AND2_X1 U18444 ( .A1(_04506_), .A2(_03047__PTR3), .ZN(_04527_) );
  AND2_X1 U18445 ( .A1(_04508_), .A2(_03047__PTR7), .ZN(_03047__PTR9) );
  AND2_X1 U18446 ( .A1(_04510_), .A2(_03047__PTR11), .ZN(_03047__PTR13) );
  AND2_X1 U18447 ( .A1(_04512_), .A2(_03047__PTR15), .ZN(_03047__PTR17) );
  AND2_X1 U18448 ( .A1(_04514_), .A2(_03047__PTR19), .ZN(_03047__PTR21) );
  AND2_X1 U18449 ( .A1(_04516_), .A2(_03047__PTR23), .ZN(_03047__PTR25) );
  AND2_X1 U18450 ( .A1(_04518_), .A2(_03047__PTR27), .ZN(_03047__PTR29) );
  AND2_X1 U18451 ( .A1(_03048__PTR2), .A2(_03047__PTR1), .ZN(_04528_) );
  AND2_X1 U18452 ( .A1(_03048__PTR4), .A2(_03047__PTR3), .ZN(_04529_) );
  AND2_X1 U18453 ( .A1(_03048__PTR6), .A2(_03047__PTR5), .ZN(_04530_) );
  AND2_X1 U18454 ( .A1(_02373__PTR40), .A2(_03047__PTR7), .ZN(_03047__PTR8) );
  AND2_X1 U18455 ( .A1(_02373__PTR42), .A2(_03047__PTR9), .ZN(_03047__PTR10) );
  AND2_X1 U18456 ( .A1(_02373__PTR44), .A2(_03047__PTR11), .ZN(_03047__PTR12) );
  AND2_X1 U18457 ( .A1(_02373__PTR46), .A2(_03047__PTR13), .ZN(_03047__PTR14) );
  AND2_X1 U18458 ( .A1(_02373__PTR48), .A2(_03047__PTR15), .ZN(_03047__PTR16) );
  AND2_X1 U18459 ( .A1(_02373__PTR50), .A2(_03047__PTR17), .ZN(_03047__PTR18) );
  AND2_X1 U18460 ( .A1(_02373__PTR52), .A2(_03047__PTR19), .ZN(_03047__PTR20) );
  AND2_X1 U18461 ( .A1(_02373__PTR54), .A2(_03047__PTR21), .ZN(_03047__PTR22) );
  AND2_X1 U18462 ( .A1(_02373__PTR56), .A2(_03047__PTR23), .ZN(_03047__PTR24) );
  AND2_X1 U18463 ( .A1(_02373__PTR58), .A2(_03047__PTR25), .ZN(_03047__PTR26) );
  AND2_X1 U18464 ( .A1(_02373__PTR60), .A2(_03047__PTR27), .ZN(_03047__PTR28) );
  AND2_X1 U18465 ( .A1(_02373__PTR62), .A2(_03047__PTR29), .ZN(_03047__PTR30) );
  OR2_X1 U18466 ( .A1(_03050__PTR1), .A2(_04498_), .ZN(_03047__PTR1) );
  OR2_X1 U18467 ( .A1(_03050__PTR3), .A2(_04499_), .ZN(_04531_) );
  OR2_X1 U18468 ( .A1(_03050__PTR5), .A2(_04500_), .ZN(_04532_) );
  OR2_X1 U18469 ( .A1(_03050__PTR7), .A2(_04501_), .ZN(_04533_) );
  OR2_X1 U18470 ( .A1(_04531_), .A2(_04502_), .ZN(_03047__PTR3) );
  OR2_X1 U18471 ( .A1(_04533_), .A2(_04503_), .ZN(_04534_) );
  OR2_X1 U18472 ( .A1(_04534_), .A2(_04504_), .ZN(_03047__PTR7) );
  OR2_X1 U18473 ( .A1(_04532_), .A2(_04527_), .ZN(_03047__PTR5) );
  OR2_X1 U18474 ( .A1(_03050__PTR2), .A2(_04528_), .ZN(_03047__PTR2) );
  OR2_X1 U18475 ( .A1(_03050__PTR4), .A2(_04529_), .ZN(_03047__PTR4) );
  OR2_X1 U18476 ( .A1(_03050__PTR6), .A2(_04530_), .ZN(_03047__PTR6) );
  AND2_X1 U18477 ( .A1(_02177__PTR3), .A2(_02968__PTR2), .ZN(_04169_) );
  AND2_X1 U18478 ( .A1(_02177__PTR5), .A2(_02968__PTR4), .ZN(_04170_) );
  AND2_X1 U18479 ( .A1(_02177__PTR7), .A2(_02968__PTR6), .ZN(_04632_) );
  AND2_X1 U18480 ( .A1(_04635_), .A2(_04182_), .ZN(_04633_) );
  AND2_X1 U18481 ( .A1(_04636_), .A2(_02969__PTR3), .ZN(_04634_) );
  AND2_X1 U18482 ( .A1(_02177__PTR7), .A2(_02177__PTR6), .ZN(_04635_) );
  AND2_X1 U18483 ( .A1(_04635_), .A2(_04175_), .ZN(_04636_) );
  AND2_X1 U18484 ( .A1(_02177__PTR4), .A2(_02969__PTR3), .ZN(_04179_) );
  OR2_X1 U18485 ( .A1(_02968__PTR3), .A2(_04169_), .ZN(_04181_) );
  OR2_X1 U18486 ( .A1(_02968__PTR7), .A2(_04632_), .ZN(_04637_) );
  OR2_X1 U18487 ( .A1(_04637_), .A2(_04633_), .ZN(_04638_) );
  OR2_X1 U18488 ( .A1(_04638_), .A2(_04634_), .ZN(_03179__PTR8) );
  OR2_X1 U18489 ( .A1(_04182_), .A2(_04178_), .ZN(_02969__PTR5) );
  AND2_X1 U18490 ( .A1(P2_P1_InstAddrPointer_PTR1), .A2(P2_P1_InstAddrPointer_PTR0), .ZN(_03043__PTR1) );
  AND2_X1 U18491 ( .A1(_04454_), .A2(_03043__PTR1), .ZN(_03043__PTR3) );
  AND2_X1 U18492 ( .A1(_04468_), .A2(_03043__PTR3), .ZN(_03043__PTR7) );
  AND2_X1 U18493 ( .A1(_04474_), .A2(_03043__PTR7), .ZN(_03043__PTR15) );
  AND2_X1 U18494 ( .A1(P2_P1_InstAddrPointer_PTR17), .A2(P2_P1_InstAddrPointer_PTR16), .ZN(_04461_) );
  AND2_X1 U18495 ( .A1(_04464_), .A2(_04463_), .ZN(_04472_) );
  AND2_X1 U18496 ( .A1(_04470_), .A2(_04469_), .ZN(_04474_) );
  AND2_X1 U18497 ( .A1(_04475_), .A2(_03043__PTR15), .ZN(_03043__PTR23) );
  AND2_X1 U18498 ( .A1(_04469_), .A2(_03043__PTR7), .ZN(_03043__PTR11) );
  AND2_X1 U18499 ( .A1(_04471_), .A2(_03043__PTR15), .ZN(_03043__PTR19) );
  AND2_X1 U18500 ( .A1(_04473_), .A2(_03043__PTR23), .ZN(_03043__PTR27) );
  AND2_X1 U18501 ( .A1(_04455_), .A2(_03043__PTR3), .ZN(_03043__PTR5) );
  AND2_X1 U18502 ( .A1(_04457_), .A2(_03043__PTR7), .ZN(_03043__PTR9) );
  AND2_X1 U18503 ( .A1(_04459_), .A2(_03043__PTR11), .ZN(_03043__PTR13) );
  AND2_X1 U18504 ( .A1(_04461_), .A2(_03043__PTR15), .ZN(_03043__PTR17) );
  AND2_X1 U18505 ( .A1(_04463_), .A2(_03043__PTR19), .ZN(_03043__PTR21) );
  AND2_X1 U18506 ( .A1(_04465_), .A2(_03043__PTR23), .ZN(_03043__PTR25) );
  AND2_X1 U18507 ( .A1(_04467_), .A2(_03043__PTR27), .ZN(_03043__PTR29) );
  AND2_X1 U18508 ( .A1(P2_P1_InstAddrPointer_PTR2), .A2(_03043__PTR1), .ZN(_03043__PTR2) );
  AND2_X1 U18509 ( .A1(P2_P1_InstAddrPointer_PTR4), .A2(_03043__PTR3), .ZN(_03043__PTR4) );
  AND2_X1 U18510 ( .A1(P2_P1_InstAddrPointer_PTR6), .A2(_03043__PTR5), .ZN(_03043__PTR6) );
  AND2_X1 U18511 ( .A1(P2_P1_InstAddrPointer_PTR8), .A2(_03043__PTR7), .ZN(_03043__PTR8) );
  AND2_X1 U18512 ( .A1(P2_P1_InstAddrPointer_PTR10), .A2(_03043__PTR9), .ZN(_03043__PTR10) );
  AND2_X1 U18513 ( .A1(P2_P1_InstAddrPointer_PTR12), .A2(_03043__PTR11), .ZN(_03043__PTR12) );
  AND2_X1 U18514 ( .A1(P2_P1_InstAddrPointer_PTR14), .A2(_03043__PTR13), .ZN(_03043__PTR14) );
  AND2_X1 U18515 ( .A1(P2_P1_InstAddrPointer_PTR16), .A2(_03043__PTR15), .ZN(_03043__PTR16) );
  AND2_X1 U18516 ( .A1(P2_P1_InstAddrPointer_PTR18), .A2(_03043__PTR17), .ZN(_03043__PTR18) );
  AND2_X1 U18517 ( .A1(P2_P1_InstAddrPointer_PTR20), .A2(_03043__PTR19), .ZN(_03043__PTR20) );
  AND2_X1 U18518 ( .A1(P2_P1_InstAddrPointer_PTR22), .A2(_03043__PTR21), .ZN(_03043__PTR22) );
  AND2_X1 U18519 ( .A1(P2_P1_InstAddrPointer_PTR24), .A2(_03043__PTR23), .ZN(_03043__PTR24) );
  AND2_X1 U18520 ( .A1(P2_P1_InstAddrPointer_PTR26), .A2(_03043__PTR25), .ZN(_03043__PTR26) );
  AND2_X1 U18521 ( .A1(P2_P1_InstAddrPointer_PTR28), .A2(_03043__PTR27), .ZN(_03043__PTR28) );
  AND2_X1 U18522 ( .A1(P2_P1_InstAddrPointer_PTR30), .A2(_03043__PTR29), .ZN(_03043__PTR30) );
  AND2_X1 U18523 ( .A1(_03054__PTR1), .A2(_03182__PTR0), .ZN(_04639_) );
  AND2_X1 U18524 ( .A1(_03183__PTR3), .A2(_03185__PTR2), .ZN(_04640_) );
  AND2_X1 U18525 ( .A1(_03183__PTR5), .A2(_03185__PTR4), .ZN(_04641_) );
  AND2_X1 U18526 ( .A1(_03183__PTR7), .A2(_03185__PTR6), .ZN(_04642_) );
  AND2_X1 U18527 ( .A1(_03183__PTR9), .A2(_03185__PTR8), .ZN(_04643_) );
  AND2_X1 U18528 ( .A1(_03183__PTR11), .A2(_03185__PTR10), .ZN(_04644_) );
  AND2_X1 U18529 ( .A1(_03183__PTR13), .A2(_03185__PTR12), .ZN(_04645_) );
  AND2_X1 U18530 ( .A1(_03183__PTR15), .A2(_03185__PTR14), .ZN(_04646_) );
  AND2_X1 U18531 ( .A1(_03183__PTR17), .A2(_03185__PTR16), .ZN(_04647_) );
  AND2_X1 U18532 ( .A1(_03183__PTR19), .A2(_03185__PTR18), .ZN(_04648_) );
  AND2_X1 U18533 ( .A1(_03183__PTR21), .A2(_03185__PTR20), .ZN(_04649_) );
  AND2_X1 U18534 ( .A1(_03183__PTR23), .A2(_03185__PTR22), .ZN(_04650_) );
  AND2_X1 U18535 ( .A1(_03183__PTR25), .A2(_03185__PTR24), .ZN(_04651_) );
  AND2_X1 U18536 ( .A1(_03183__PTR27), .A2(_03185__PTR26), .ZN(_04652_) );
  AND2_X1 U18537 ( .A1(_03183__PTR29), .A2(_03185__PTR28), .ZN(_04653_) );
  AND2_X1 U18538 ( .A1(_04665_), .A2(_03182__PTR1), .ZN(_04654_) );
  AND2_X1 U18539 ( .A1(_04667_), .A2(_04714_), .ZN(_04655_) );
  AND2_X1 U18540 ( .A1(_04669_), .A2(_04716_), .ZN(_04656_) );
  AND2_X1 U18541 ( .A1(_04671_), .A2(_04718_), .ZN(_04657_) );
  AND2_X1 U18542 ( .A1(_04673_), .A2(_04720_), .ZN(_04658_) );
  AND2_X1 U18543 ( .A1(_04675_), .A2(_04722_), .ZN(_04659_) );
  AND2_X1 U18544 ( .A1(_04677_), .A2(_04724_), .ZN(_04660_) );
  AND2_X1 U18545 ( .A1(_04679_), .A2(_03182__PTR3), .ZN(_04661_) );
  AND2_X1 U18546 ( .A1(_04681_), .A2(_04728_), .ZN(_04662_) );
  AND2_X1 U18547 ( .A1(_04683_), .A2(_04730_), .ZN(_04663_) );
  AND2_X1 U18548 ( .A1(_04685_), .A2(_03182__PTR7), .ZN(_04664_) );
  AND2_X1 U18549 ( .A1(_03183__PTR3), .A2(_03183__PTR2), .ZN(_04665_) );
  AND2_X1 U18550 ( .A1(_03183__PTR5), .A2(_03183__PTR4), .ZN(_04666_) );
  AND2_X1 U18551 ( .A1(_03183__PTR7), .A2(_03183__PTR6), .ZN(_04667_) );
  AND2_X1 U18552 ( .A1(_03183__PTR9), .A2(_03183__PTR8), .ZN(_04668_) );
  AND2_X1 U18553 ( .A1(_03183__PTR11), .A2(_03183__PTR10), .ZN(_04669_) );
  AND2_X1 U18554 ( .A1(_03183__PTR13), .A2(_03183__PTR12), .ZN(_04670_) );
  AND2_X1 U18555 ( .A1(_03183__PTR15), .A2(_03183__PTR14), .ZN(_04671_) );
  AND2_X1 U18556 ( .A1(_03183__PTR17), .A2(_03183__PTR16), .ZN(_04672_) );
  AND2_X1 U18557 ( .A1(_03183__PTR19), .A2(_03183__PTR18), .ZN(_04673_) );
  AND2_X1 U18558 ( .A1(_03183__PTR21), .A2(_03183__PTR20), .ZN(_04674_) );
  AND2_X1 U18559 ( .A1(_03183__PTR23), .A2(_03183__PTR22), .ZN(_04675_) );
  AND2_X1 U18560 ( .A1(_03183__PTR25), .A2(_03183__PTR24), .ZN(_04676_) );
  AND2_X1 U18561 ( .A1(_03183__PTR27), .A2(_03183__PTR26), .ZN(_04677_) );
  AND2_X1 U18562 ( .A1(_03183__PTR29), .A2(_03183__PTR28), .ZN(_04678_) );
  AND2_X1 U18563 ( .A1(_04667_), .A2(_04666_), .ZN(_04679_) );
  AND2_X1 U18564 ( .A1(_04669_), .A2(_04668_), .ZN(_04680_) );
  AND2_X1 U18565 ( .A1(_04671_), .A2(_04670_), .ZN(_04681_) );
  AND2_X1 U18566 ( .A1(_04673_), .A2(_04672_), .ZN(_04682_) );
  AND2_X1 U18567 ( .A1(_04675_), .A2(_04674_), .ZN(_04683_) );
  AND2_X1 U18568 ( .A1(_04677_), .A2(_04676_), .ZN(_04684_) );
  AND2_X1 U18569 ( .A1(_04681_), .A2(_04680_), .ZN(_04685_) );
  AND2_X1 U18570 ( .A1(_04683_), .A2(_04682_), .ZN(_04686_) );
  AND2_X1 U18571 ( .A1(_04686_), .A2(_03182__PTR15), .ZN(_04687_) );
  AND2_X1 U18572 ( .A1(_04680_), .A2(_03182__PTR7), .ZN(_04688_) );
  AND2_X1 U18573 ( .A1(_04682_), .A2(_03182__PTR15), .ZN(_04689_) );
  AND2_X1 U18574 ( .A1(_04684_), .A2(_03182__PTR23), .ZN(_04690_) );
  AND2_X1 U18575 ( .A1(_04666_), .A2(_03182__PTR3), .ZN(_04691_) );
  AND2_X1 U18576 ( .A1(_04668_), .A2(_03182__PTR7), .ZN(_04692_) );
  AND2_X1 U18577 ( .A1(_04670_), .A2(_03182__PTR11), .ZN(_04693_) );
  AND2_X1 U18578 ( .A1(_04672_), .A2(_03182__PTR15), .ZN(_04694_) );
  AND2_X1 U18579 ( .A1(_04674_), .A2(_03182__PTR19), .ZN(_04695_) );
  AND2_X1 U18580 ( .A1(_04676_), .A2(_03182__PTR23), .ZN(_04696_) );
  AND2_X1 U18581 ( .A1(_04678_), .A2(_03182__PTR27), .ZN(_04697_) );
  AND2_X1 U18582 ( .A1(_03183__PTR2), .A2(_03182__PTR1), .ZN(_04698_) );
  AND2_X1 U18583 ( .A1(_03183__PTR4), .A2(_03182__PTR3), .ZN(_04699_) );
  AND2_X1 U18584 ( .A1(_03183__PTR6), .A2(_03182__PTR5), .ZN(_04700_) );
  AND2_X1 U18585 ( .A1(_03183__PTR8), .A2(_03182__PTR7), .ZN(_04701_) );
  AND2_X1 U18586 ( .A1(_03183__PTR10), .A2(_03182__PTR9), .ZN(_04702_) );
  AND2_X1 U18587 ( .A1(_03183__PTR12), .A2(_03182__PTR11), .ZN(_04703_) );
  AND2_X1 U18588 ( .A1(_03183__PTR14), .A2(_03182__PTR13), .ZN(_04704_) );
  AND2_X1 U18589 ( .A1(_03183__PTR16), .A2(_03182__PTR15), .ZN(_04705_) );
  AND2_X1 U18590 ( .A1(_03183__PTR18), .A2(_03182__PTR17), .ZN(_04706_) );
  AND2_X1 U18591 ( .A1(_03183__PTR20), .A2(_03182__PTR19), .ZN(_04707_) );
  AND2_X1 U18592 ( .A1(_03183__PTR22), .A2(_03182__PTR21), .ZN(_04708_) );
  AND2_X1 U18593 ( .A1(_03183__PTR24), .A2(_03182__PTR23), .ZN(_04709_) );
  AND2_X1 U18594 ( .A1(_03183__PTR26), .A2(_03182__PTR25), .ZN(_04710_) );
  AND2_X1 U18595 ( .A1(_03183__PTR28), .A2(_03182__PTR27), .ZN(_04711_) );
  AND2_X1 U18596 ( .A1(_03183__PTR30), .A2(_03182__PTR29), .ZN(_04712_) );
  OR2_X1 U18597 ( .A1(_03053__PTR0), .A2(_03054__PTR0), .ZN(_03182__PTR0) );
  OR2_X1 U18598 ( .A1(_03056__PTR1), .A2(_04639_), .ZN(_03182__PTR1) );
  OR2_X1 U18599 ( .A1(_03185__PTR3), .A2(_04640_), .ZN(_04713_) );
  OR2_X1 U18600 ( .A1(_03185__PTR5), .A2(_04641_), .ZN(_04714_) );
  OR2_X1 U18601 ( .A1(_03185__PTR7), .A2(_04642_), .ZN(_04715_) );
  OR2_X1 U18602 ( .A1(_03185__PTR9), .A2(_04643_), .ZN(_04716_) );
  OR2_X1 U18603 ( .A1(_03185__PTR11), .A2(_04644_), .ZN(_04717_) );
  OR2_X1 U18604 ( .A1(_03185__PTR13), .A2(_04645_), .ZN(_04718_) );
  OR2_X1 U18605 ( .A1(_03185__PTR15), .A2(_04646_), .ZN(_04719_) );
  OR2_X1 U18606 ( .A1(_03185__PTR17), .A2(_04647_), .ZN(_04720_) );
  OR2_X1 U18607 ( .A1(_03185__PTR19), .A2(_04648_), .ZN(_04721_) );
  OR2_X1 U18608 ( .A1(_03185__PTR21), .A2(_04649_), .ZN(_04722_) );
  OR2_X1 U18609 ( .A1(_03185__PTR23), .A2(_04650_), .ZN(_04723_) );
  OR2_X1 U18610 ( .A1(_03185__PTR25), .A2(_04651_), .ZN(_04724_) );
  OR2_X1 U18611 ( .A1(_03185__PTR27), .A2(_04652_), .ZN(_04725_) );
  OR2_X1 U18612 ( .A1(_03185__PTR29), .A2(_04653_), .ZN(_04726_) );
  OR2_X1 U18613 ( .A1(_04713_), .A2(_04654_), .ZN(_03182__PTR3) );
  OR2_X1 U18614 ( .A1(_04715_), .A2(_04655_), .ZN(_04727_) );
  OR2_X1 U18615 ( .A1(_04717_), .A2(_04656_), .ZN(_04728_) );
  OR2_X1 U18616 ( .A1(_04719_), .A2(_04657_), .ZN(_04729_) );
  OR2_X1 U18617 ( .A1(_04721_), .A2(_04658_), .ZN(_04730_) );
  OR2_X1 U18618 ( .A1(_04723_), .A2(_04659_), .ZN(_04731_) );
  OR2_X1 U18619 ( .A1(_04725_), .A2(_04660_), .ZN(_04732_) );
  OR2_X1 U18620 ( .A1(_04727_), .A2(_04661_), .ZN(_03182__PTR7) );
  OR2_X1 U18621 ( .A1(_04729_), .A2(_04662_), .ZN(_04733_) );
  OR2_X1 U18622 ( .A1(_04731_), .A2(_04663_), .ZN(_04734_) );
  OR2_X1 U18623 ( .A1(_04733_), .A2(_04664_), .ZN(_03182__PTR15) );
  OR2_X1 U18624 ( .A1(_04734_), .A2(_04687_), .ZN(_03182__PTR23) );
  OR2_X1 U18625 ( .A1(_04728_), .A2(_04688_), .ZN(_03182__PTR11) );
  OR2_X1 U18626 ( .A1(_04730_), .A2(_04689_), .ZN(_03182__PTR19) );
  OR2_X1 U18627 ( .A1(_04732_), .A2(_04690_), .ZN(_03182__PTR27) );
  OR2_X1 U18628 ( .A1(_04714_), .A2(_04691_), .ZN(_03182__PTR5) );
  OR2_X1 U18629 ( .A1(_04716_), .A2(_04692_), .ZN(_03182__PTR9) );
  OR2_X1 U18630 ( .A1(_04718_), .A2(_04693_), .ZN(_03182__PTR13) );
  OR2_X1 U18631 ( .A1(_04720_), .A2(_04694_), .ZN(_03182__PTR17) );
  OR2_X1 U18632 ( .A1(_04722_), .A2(_04695_), .ZN(_03182__PTR21) );
  OR2_X1 U18633 ( .A1(_04724_), .A2(_04696_), .ZN(_03182__PTR25) );
  OR2_X1 U18634 ( .A1(_04726_), .A2(_04697_), .ZN(_03182__PTR29) );
  OR2_X1 U18635 ( .A1(_03185__PTR2), .A2(_04698_), .ZN(_03182__PTR2) );
  OR2_X1 U18636 ( .A1(_03185__PTR4), .A2(_04699_), .ZN(_03182__PTR4) );
  OR2_X1 U18637 ( .A1(_03185__PTR6), .A2(_04700_), .ZN(_03182__PTR6) );
  OR2_X1 U18638 ( .A1(_03185__PTR8), .A2(_04701_), .ZN(_03182__PTR8) );
  OR2_X1 U18639 ( .A1(_03185__PTR10), .A2(_04702_), .ZN(_03182__PTR10) );
  OR2_X1 U18640 ( .A1(_03185__PTR12), .A2(_04703_), .ZN(_03182__PTR12) );
  OR2_X1 U18641 ( .A1(_03185__PTR14), .A2(_04704_), .ZN(_03182__PTR14) );
  OR2_X1 U18642 ( .A1(_03185__PTR16), .A2(_04705_), .ZN(_03182__PTR16) );
  OR2_X1 U18643 ( .A1(_03185__PTR18), .A2(_04706_), .ZN(_03182__PTR18) );
  OR2_X1 U18644 ( .A1(_03185__PTR20), .A2(_04707_), .ZN(_03182__PTR20) );
  OR2_X1 U18645 ( .A1(_03185__PTR22), .A2(_04708_), .ZN(_03182__PTR22) );
  OR2_X1 U18646 ( .A1(_03185__PTR24), .A2(_04709_), .ZN(_03182__PTR24) );
  OR2_X1 U18647 ( .A1(_03185__PTR26), .A2(_04710_), .ZN(_03182__PTR26) );
  OR2_X1 U18648 ( .A1(_03185__PTR28), .A2(_04711_), .ZN(_03182__PTR28) );
  OR2_X1 U18649 ( .A1(_03185__PTR30), .A2(_04712_), .ZN(_03182__PTR30) );
  AND2_X1 U18650 ( .A1(_02968__PTR7), .A2(_02968__PTR6), .ZN(_04171_) );
  AND2_X1 U18651 ( .A1(_04176_), .A2(_04182_), .ZN(_04173_) );
  AND2_X1 U18652 ( .A1(_04177_), .A2(_02969__PTR3), .ZN(_04174_) );
  AND2_X1 U18653 ( .A1(_02177__PTR3), .A2(_02177__PTR2), .ZN(_04172_) );
  AND2_X1 U18654 ( .A1(_02177__PTR5), .A2(_02177__PTR4), .ZN(_04175_) );
  AND2_X1 U18655 ( .A1(_02968__PTR7), .A2(_02177__PTR6), .ZN(_04176_) );
  AND2_X1 U18656 ( .A1(_04176_), .A2(_04175_), .ZN(_04177_) );
  AND2_X1 U18657 ( .A1(_04175_), .A2(_02969__PTR3), .ZN(_04178_) );
  AND2_X1 U18658 ( .A1(_02177__PTR6), .A2(_02969__PTR5), .ZN(_04180_) );
  OR2_X1 U18659 ( .A1(_02968__PTR5), .A2(_04170_), .ZN(_04182_) );
  OR2_X1 U18660 ( .A1(_04181_), .A2(_04172_), .ZN(_02969__PTR3) );
  OR2_X1 U18661 ( .A1(_04171_), .A2(_04173_), .ZN(_04183_) );
  OR2_X1 U18662 ( .A1(_04183_), .A2(_04174_), .ZN(_02969__PTR7) );
  OR2_X1 U18663 ( .A1(_02968__PTR4), .A2(_04179_), .ZN(_02969__PTR4) );
  OR2_X1 U18664 ( .A1(_02968__PTR6), .A2(_04180_), .ZN(_02969__PTR6) );
  AND2_X1 U18665 ( .A1(_02963__PTR3), .A2(_02963__PTR2), .ZN(_02964__PTR3) );
  AND2_X1 U18666 ( .A1(_00942__PTR2), .A2(_02964__PTR3), .ZN(_04168_) );
  OR2_X1 U18667 ( .A1(_02961__PTR5), .A2(_04168_), .ZN(_02964__PTR5) );
  AND2_X1 U18668 ( .A1(_03057__PTR1), .A2(_02995__PTR1), .ZN(_02995__PTR3) );
  AND2_X1 U18669 ( .A1(P2_P1_InstQueueRd_Addr_PTR3), .A2(P2_P1_InstQueueRd_Addr_PTR2), .ZN(_03057__PTR1) );
  AND2_X1 U18670 ( .A1(P2_P1_InstQueueRd_Addr_PTR2), .A2(_02995__PTR1), .ZN(_02995__PTR2) );
  AND2_X1 U18671 ( .A1(P2_P1_InstQueueRd_Addr_PTR4), .A2(_02995__PTR3), .ZN(_03044__PTR4) );
  AND2_X1 U18672 ( .A1(P2_P1_PhyAddrPointer_PTR2), .A2(P2_P1_PhyAddrPointer_PTR1), .ZN(_03042__PTR1) );
  AND2_X1 U18673 ( .A1(_04432_), .A2(_03042__PTR1), .ZN(_03042__PTR3) );
  AND2_X1 U18674 ( .A1(_04446_), .A2(_03042__PTR3), .ZN(_03042__PTR7) );
  AND2_X1 U18675 ( .A1(_04452_), .A2(_03042__PTR7), .ZN(_03042__PTR15) );
  AND2_X1 U18676 ( .A1(P2_P1_PhyAddrPointer_PTR4), .A2(P2_P1_PhyAddrPointer_PTR3), .ZN(_04432_) );
  AND2_X1 U18677 ( .A1(P2_P1_PhyAddrPointer_PTR6), .A2(P2_P1_PhyAddrPointer_PTR5), .ZN(_04433_) );
  AND2_X1 U18678 ( .A1(P2_P1_PhyAddrPointer_PTR8), .A2(P2_P1_PhyAddrPointer_PTR7), .ZN(_04434_) );
  AND2_X1 U18679 ( .A1(P2_P1_PhyAddrPointer_PTR10), .A2(P2_P1_PhyAddrPointer_PTR9), .ZN(_04435_) );
  AND2_X1 U18680 ( .A1(P2_P1_PhyAddrPointer_PTR12), .A2(P2_P1_PhyAddrPointer_PTR11), .ZN(_04436_) );
  AND2_X1 U18681 ( .A1(P2_P1_PhyAddrPointer_PTR14), .A2(P2_P1_PhyAddrPointer_PTR13), .ZN(_04437_) );
  AND2_X1 U18682 ( .A1(P2_P1_PhyAddrPointer_PTR16), .A2(P2_P1_PhyAddrPointer_PTR15), .ZN(_04438_) );
  AND2_X1 U18683 ( .A1(P2_P1_PhyAddrPointer_PTR18), .A2(P2_P1_PhyAddrPointer_PTR17), .ZN(_04439_) );
  AND2_X1 U18684 ( .A1(P2_P1_PhyAddrPointer_PTR20), .A2(P2_P1_PhyAddrPointer_PTR19), .ZN(_04440_) );
  AND2_X1 U18685 ( .A1(P2_P1_PhyAddrPointer_PTR22), .A2(P2_P1_PhyAddrPointer_PTR21), .ZN(_04441_) );
  AND2_X1 U18686 ( .A1(P2_P1_PhyAddrPointer_PTR24), .A2(P2_P1_PhyAddrPointer_PTR23), .ZN(_04442_) );
  AND2_X1 U18687 ( .A1(P2_P1_PhyAddrPointer_PTR26), .A2(P2_P1_PhyAddrPointer_PTR25), .ZN(_04443_) );
  AND2_X1 U18688 ( .A1(P2_P1_PhyAddrPointer_PTR28), .A2(P2_P1_PhyAddrPointer_PTR27), .ZN(_04444_) );
  AND2_X1 U18689 ( .A1(P2_P1_PhyAddrPointer_PTR30), .A2(P2_P1_PhyAddrPointer_PTR29), .ZN(_04445_) );
  AND2_X1 U18690 ( .A1(_04434_), .A2(_04433_), .ZN(_04446_) );
  AND2_X1 U18691 ( .A1(_04436_), .A2(_04435_), .ZN(_04447_) );
  AND2_X1 U18692 ( .A1(_04438_), .A2(_04437_), .ZN(_04448_) );
  AND2_X1 U18693 ( .A1(_04440_), .A2(_04439_), .ZN(_04449_) );
  AND2_X1 U18694 ( .A1(_04442_), .A2(_04441_), .ZN(_04450_) );
  AND2_X1 U18695 ( .A1(_04444_), .A2(_04443_), .ZN(_04451_) );
  AND2_X1 U18696 ( .A1(_04448_), .A2(_04447_), .ZN(_04452_) );
  AND2_X1 U18697 ( .A1(_04450_), .A2(_04449_), .ZN(_04453_) );
  AND2_X1 U18698 ( .A1(_04453_), .A2(_03042__PTR15), .ZN(_03042__PTR23) );
  AND2_X1 U18699 ( .A1(_04447_), .A2(_03042__PTR7), .ZN(_03042__PTR11) );
  AND2_X1 U18700 ( .A1(_04449_), .A2(_03042__PTR15), .ZN(_03042__PTR19) );
  AND2_X1 U18701 ( .A1(_04451_), .A2(_03042__PTR23), .ZN(_03042__PTR27) );
  AND2_X1 U18702 ( .A1(_04433_), .A2(_03042__PTR3), .ZN(_03042__PTR5) );
  AND2_X1 U18703 ( .A1(_04435_), .A2(_03042__PTR7), .ZN(_03042__PTR9) );
  AND2_X1 U18704 ( .A1(_04437_), .A2(_03042__PTR11), .ZN(_03042__PTR13) );
  AND2_X1 U18705 ( .A1(_04439_), .A2(_03042__PTR15), .ZN(_03042__PTR17) );
  AND2_X1 U18706 ( .A1(_04441_), .A2(_03042__PTR19), .ZN(_03042__PTR21) );
  AND2_X1 U18707 ( .A1(_04443_), .A2(_03042__PTR23), .ZN(_03042__PTR25) );
  AND2_X1 U18708 ( .A1(_04445_), .A2(_03042__PTR27), .ZN(_03042__PTR29) );
  AND2_X1 U18709 ( .A1(P2_P1_PhyAddrPointer_PTR3), .A2(_03042__PTR1), .ZN(_03042__PTR2) );
  AND2_X1 U18710 ( .A1(P2_P1_PhyAddrPointer_PTR5), .A2(_03042__PTR3), .ZN(_03042__PTR4) );
  AND2_X1 U18711 ( .A1(P2_P1_PhyAddrPointer_PTR7), .A2(_03042__PTR5), .ZN(_03042__PTR6) );
  AND2_X1 U18712 ( .A1(P2_P1_PhyAddrPointer_PTR9), .A2(_03042__PTR7), .ZN(_03042__PTR8) );
  AND2_X1 U18713 ( .A1(P2_P1_PhyAddrPointer_PTR11), .A2(_03042__PTR9), .ZN(_03042__PTR10) );
  AND2_X1 U18714 ( .A1(P2_P1_PhyAddrPointer_PTR13), .A2(_03042__PTR11), .ZN(_03042__PTR12) );
  AND2_X1 U18715 ( .A1(P2_P1_PhyAddrPointer_PTR15), .A2(_03042__PTR13), .ZN(_03042__PTR14) );
  AND2_X1 U18716 ( .A1(P2_P1_PhyAddrPointer_PTR17), .A2(_03042__PTR15), .ZN(_03042__PTR16) );
  AND2_X1 U18717 ( .A1(P2_P1_PhyAddrPointer_PTR19), .A2(_03042__PTR17), .ZN(_03042__PTR18) );
  AND2_X1 U18718 ( .A1(P2_P1_PhyAddrPointer_PTR21), .A2(_03042__PTR19), .ZN(_03042__PTR20) );
  AND2_X1 U18719 ( .A1(P2_P1_PhyAddrPointer_PTR23), .A2(_03042__PTR21), .ZN(_03042__PTR22) );
  AND2_X1 U18720 ( .A1(P2_P1_PhyAddrPointer_PTR25), .A2(_03042__PTR23), .ZN(_03042__PTR24) );
  AND2_X1 U18721 ( .A1(P2_P1_PhyAddrPointer_PTR27), .A2(_03042__PTR25), .ZN(_03042__PTR26) );
  AND2_X1 U18722 ( .A1(P2_P1_PhyAddrPointer_PTR29), .A2(_03042__PTR27), .ZN(_03042__PTR28) );
  AND2_X1 U18723 ( .A1(P2_P1_PhyAddrPointer_PTR1), .A2(_02960__PTR0), .ZN(_03190__PTR1) );
  AND2_X1 U18724 ( .A1(_04103_), .A2(_03190__PTR1), .ZN(_03190__PTR3) );
  AND2_X1 U18725 ( .A1(_04132_), .A2(_03190__PTR3), .ZN(_03190__PTR7) );
  AND2_X1 U18726 ( .A1(_04139_), .A2(_03190__PTR7), .ZN(_03190__PTR15) );
  AND2_X1 U18727 ( .A1(_02960__PTR3), .A2(_02960__PTR2), .ZN(_04103_) );
  AND2_X1 U18728 ( .A1(_02960__PTR5), .A2(_02960__PTR4), .ZN(_04118_) );
  AND2_X1 U18729 ( .A1(_02960__PTR7), .A2(_02960__PTR6), .ZN(_04119_) );
  AND2_X1 U18730 ( .A1(_02960__PTR11), .A2(_02960__PTR10), .ZN(_04121_) );
  AND2_X1 U18731 ( .A1(_02960__PTR19), .A2(_02960__PTR18), .ZN(_04125_) );
  AND2_X1 U18732 ( .A1(_02960__PTR21), .A2(_02960__PTR20), .ZN(_04126_) );
  AND2_X1 U18733 ( .A1(_02960__PTR27), .A2(_02960__PTR26), .ZN(_04129_) );
  AND2_X1 U18734 ( .A1(_02958__PTR31), .A2(_02960__PTR30), .ZN(_04131_) );
  AND2_X1 U18735 ( .A1(_04119_), .A2(_04118_), .ZN(_04132_) );
  AND2_X1 U18736 ( .A1(_04121_), .A2(_04120_), .ZN(_04133_) );
  AND2_X1 U18737 ( .A1(_04123_), .A2(_04122_), .ZN(_04134_) );
  AND2_X1 U18738 ( .A1(_04125_), .A2(_04124_), .ZN(_04135_) );
  AND2_X1 U18739 ( .A1(_04129_), .A2(_04128_), .ZN(_04137_) );
  AND2_X1 U18740 ( .A1(_04136_), .A2(_04135_), .ZN(_04140_) );
  AND2_X1 U18741 ( .A1(_04141_), .A2(_04140_), .ZN(_04142_) );
  AND2_X1 U18742 ( .A1(_04140_), .A2(_03190__PTR15), .ZN(_03190__PTR23) );
  AND2_X1 U18743 ( .A1(_04133_), .A2(_03190__PTR7), .ZN(_03190__PTR11) );
  AND2_X1 U18744 ( .A1(_04135_), .A2(_03190__PTR15), .ZN(_03190__PTR19) );
  AND2_X1 U18745 ( .A1(_04137_), .A2(_03190__PTR23), .ZN(_03190__PTR27) );
  AND2_X1 U18746 ( .A1(_04118_), .A2(_03190__PTR3), .ZN(_03190__PTR5) );
  AND2_X1 U18747 ( .A1(_04120_), .A2(_03190__PTR7), .ZN(_03190__PTR9) );
  AND2_X1 U18748 ( .A1(_04122_), .A2(_03190__PTR11), .ZN(_03190__PTR13) );
  AND2_X1 U18749 ( .A1(_04124_), .A2(_03190__PTR15), .ZN(_03190__PTR17) );
  AND2_X1 U18750 ( .A1(_04126_), .A2(_03190__PTR19), .ZN(_03190__PTR21) );
  AND2_X1 U18751 ( .A1(_04128_), .A2(_03190__PTR23), .ZN(_03190__PTR25) );
  AND2_X1 U18752 ( .A1(_04130_), .A2(_03190__PTR27), .ZN(_03190__PTR29) );
  AND2_X1 U18753 ( .A1(_02960__PTR2), .A2(_03190__PTR1), .ZN(_03190__PTR2) );
  AND2_X1 U18754 ( .A1(_02960__PTR4), .A2(_03190__PTR3), .ZN(_03190__PTR4) );
  AND2_X1 U18755 ( .A1(_02960__PTR6), .A2(_03190__PTR5), .ZN(_03190__PTR6) );
  AND2_X1 U18756 ( .A1(_02960__PTR8), .A2(_03190__PTR7), .ZN(_03190__PTR8) );
  AND2_X1 U18757 ( .A1(_02960__PTR10), .A2(_03190__PTR9), .ZN(_03190__PTR10) );
  AND2_X1 U18758 ( .A1(_02960__PTR12), .A2(_03190__PTR11), .ZN(_03190__PTR12) );
  AND2_X1 U18759 ( .A1(_02960__PTR14), .A2(_03190__PTR13), .ZN(_03190__PTR14) );
  AND2_X1 U18760 ( .A1(_02960__PTR16), .A2(_03190__PTR15), .ZN(_03190__PTR16) );
  AND2_X1 U18761 ( .A1(_02960__PTR18), .A2(_03190__PTR17), .ZN(_03190__PTR18) );
  AND2_X1 U18762 ( .A1(_02960__PTR20), .A2(_03190__PTR19), .ZN(_03190__PTR20) );
  AND2_X1 U18763 ( .A1(_02960__PTR22), .A2(_03190__PTR21), .ZN(_03190__PTR22) );
  AND2_X1 U18764 ( .A1(_02960__PTR24), .A2(_03190__PTR23), .ZN(_03190__PTR24) );
  AND2_X1 U18765 ( .A1(_02960__PTR26), .A2(_03190__PTR25), .ZN(_03190__PTR26) );
  AND2_X1 U18766 ( .A1(_02960__PTR28), .A2(_03190__PTR27), .ZN(_03190__PTR28) );
  AND2_X1 U18767 ( .A1(_02960__PTR30), .A2(_03190__PTR29), .ZN(_03190__PTR30) );
  AND2_X1 U18768 ( .A1(_02960__PTR3), .A2(_02184__PTR130), .ZN(_04088_) );
  AND2_X1 U18769 ( .A1(_02960__PTR5), .A2(_02184__PTR132), .ZN(_04089_) );
  AND2_X1 U18770 ( .A1(_02960__PTR7), .A2(_02184__PTR134), .ZN(_04090_) );
  AND2_X1 U18771 ( .A1(_02960__PTR9), .A2(_02184__PTR136), .ZN(_04091_) );
  AND2_X1 U18772 ( .A1(_02960__PTR11), .A2(_02184__PTR138), .ZN(_04092_) );
  AND2_X1 U18773 ( .A1(_02960__PTR13), .A2(_02184__PTR140), .ZN(_04093_) );
  AND2_X1 U18774 ( .A1(_02960__PTR15), .A2(_02184__PTR142), .ZN(_04094_) );
  AND2_X1 U18775 ( .A1(_02960__PTR17), .A2(_02184__PTR144), .ZN(_04095_) );
  AND2_X1 U18776 ( .A1(_02960__PTR19), .A2(_02184__PTR146), .ZN(_04096_) );
  AND2_X1 U18777 ( .A1(_02960__PTR21), .A2(_02184__PTR148), .ZN(_04097_) );
  AND2_X1 U18778 ( .A1(_02960__PTR23), .A2(_02184__PTR150), .ZN(_04098_) );
  AND2_X1 U18779 ( .A1(_02960__PTR25), .A2(_02184__PTR152), .ZN(_04099_) );
  AND2_X1 U18780 ( .A1(_02960__PTR27), .A2(_02184__PTR154), .ZN(_04100_) );
  AND2_X1 U18781 ( .A1(_02960__PTR29), .A2(_02184__PTR156), .ZN(_04101_) );
  AND2_X1 U18782 ( .A1(_02958__PTR31), .A2(_02184__PTR158), .ZN(_04102_) );
  AND2_X1 U18783 ( .A1(_04119_), .A2(_04144_), .ZN(_04104_) );
  AND2_X1 U18784 ( .A1(_04121_), .A2(_04146_), .ZN(_04105_) );
  AND2_X1 U18785 ( .A1(_04123_), .A2(_04148_), .ZN(_04106_) );
  AND2_X1 U18786 ( .A1(_04125_), .A2(_04150_), .ZN(_04107_) );
  AND2_X1 U18787 ( .A1(_04127_), .A2(_04152_), .ZN(_04108_) );
  AND2_X1 U18788 ( .A1(_04129_), .A2(_04154_), .ZN(_04109_) );
  AND2_X1 U18789 ( .A1(_04131_), .A2(_04156_), .ZN(_04110_) );
  AND2_X1 U18790 ( .A1(_04132_), .A2(_02959__PTR3), .ZN(_04111_) );
  AND2_X1 U18791 ( .A1(_04134_), .A2(_04158_), .ZN(_04112_) );
  AND2_X1 U18792 ( .A1(_04136_), .A2(_04160_), .ZN(_04113_) );
  AND2_X1 U18793 ( .A1(_04138_), .A2(_04162_), .ZN(_04114_) );
  AND2_X1 U18794 ( .A1(_04139_), .A2(_02959__PTR7), .ZN(_04115_) );
  AND2_X1 U18795 ( .A1(_04141_), .A2(_04165_), .ZN(_04116_) );
  AND2_X1 U18796 ( .A1(_04142_), .A2(_02959__PTR15), .ZN(_04117_) );
  AND2_X1 U18797 ( .A1(_02960__PTR9), .A2(_02960__PTR8), .ZN(_04120_) );
  AND2_X1 U18798 ( .A1(_02960__PTR13), .A2(_02960__PTR12), .ZN(_04122_) );
  AND2_X1 U18799 ( .A1(_02960__PTR15), .A2(_02960__PTR14), .ZN(_04123_) );
  AND2_X1 U18800 ( .A1(_02960__PTR17), .A2(_02960__PTR16), .ZN(_04124_) );
  AND2_X1 U18801 ( .A1(_02960__PTR23), .A2(_02960__PTR22), .ZN(_04127_) );
  AND2_X1 U18802 ( .A1(_02960__PTR25), .A2(_02960__PTR24), .ZN(_04128_) );
  AND2_X1 U18803 ( .A1(_02960__PTR29), .A2(_02960__PTR28), .ZN(_04130_) );
  AND2_X1 U18804 ( .A1(_04127_), .A2(_04126_), .ZN(_04136_) );
  AND2_X1 U18805 ( .A1(_04131_), .A2(_04130_), .ZN(_04138_) );
  AND2_X1 U18806 ( .A1(_04134_), .A2(_04133_), .ZN(_04139_) );
  AND2_X1 U18807 ( .A1(_04138_), .A2(_04137_), .ZN(_04141_) );
  OR2_X1 U18808 ( .A1(_02184__PTR131), .A2(_04088_), .ZN(_04143_) );
  OR2_X1 U18809 ( .A1(_02184__PTR133), .A2(_04089_), .ZN(_04144_) );
  OR2_X1 U18810 ( .A1(_02184__PTR135), .A2(_04090_), .ZN(_04145_) );
  OR2_X1 U18811 ( .A1(_02184__PTR137), .A2(_04091_), .ZN(_04146_) );
  OR2_X1 U18812 ( .A1(_02184__PTR139), .A2(_04092_), .ZN(_04147_) );
  OR2_X1 U18813 ( .A1(_02184__PTR141), .A2(_04093_), .ZN(_04148_) );
  OR2_X1 U18814 ( .A1(_02184__PTR143), .A2(_04094_), .ZN(_04149_) );
  OR2_X1 U18815 ( .A1(_02184__PTR145), .A2(_04095_), .ZN(_04150_) );
  OR2_X1 U18816 ( .A1(_02184__PTR147), .A2(_04096_), .ZN(_04151_) );
  OR2_X1 U18817 ( .A1(_02184__PTR149), .A2(_04097_), .ZN(_04152_) );
  OR2_X1 U18818 ( .A1(_02184__PTR151), .A2(_04098_), .ZN(_04153_) );
  OR2_X1 U18819 ( .A1(_02184__PTR153), .A2(_04099_), .ZN(_04154_) );
  OR2_X1 U18820 ( .A1(_02184__PTR155), .A2(_04100_), .ZN(_04155_) );
  OR2_X1 U18821 ( .A1(_02184__PTR157), .A2(_04101_), .ZN(_04156_) );
  OR2_X1 U18822 ( .A1(_04143_), .A2(_04103_), .ZN(_02959__PTR3) );
  OR2_X1 U18823 ( .A1(_04145_), .A2(_04104_), .ZN(_04157_) );
  OR2_X1 U18824 ( .A1(_04147_), .A2(_04105_), .ZN(_04158_) );
  OR2_X1 U18825 ( .A1(_04149_), .A2(_04106_), .ZN(_04159_) );
  OR2_X1 U18826 ( .A1(_04151_), .A2(_04107_), .ZN(_04160_) );
  OR2_X1 U18827 ( .A1(_04153_), .A2(_04108_), .ZN(_04161_) );
  OR2_X1 U18828 ( .A1(_04155_), .A2(_04109_), .ZN(_04162_) );
  OR2_X1 U18829 ( .A1(_04102_), .A2(_04110_), .ZN(_04163_) );
  OR2_X1 U18830 ( .A1(_04157_), .A2(_04111_), .ZN(_02959__PTR7) );
  OR2_X1 U18831 ( .A1(_04159_), .A2(_04112_), .ZN(_04164_) );
  OR2_X1 U18832 ( .A1(_04161_), .A2(_04113_), .ZN(_04165_) );
  OR2_X1 U18833 ( .A1(_04163_), .A2(_04114_), .ZN(_04166_) );
  OR2_X1 U18834 ( .A1(_04164_), .A2(_04115_), .ZN(_02959__PTR15) );
  OR2_X1 U18835 ( .A1(_04166_), .A2(_04116_), .ZN(_04167_) );
  OR2_X1 U18836 ( .A1(_04167_), .A2(_04117_), .ZN(_02959__PTR31) );
  AND2_X1 U18837 ( .A1(P2_P1_PhyAddrPointer_PTR3), .A2(P2_P1_PhyAddrPointer_PTR2), .ZN(_03039__PTR1) );
  AND2_X1 U18838 ( .A1(_04411_), .A2(_03039__PTR1), .ZN(_03039__PTR3) );
  AND2_X1 U18839 ( .A1(_04424_), .A2(_03039__PTR3), .ZN(_03039__PTR7) );
  AND2_X1 U18840 ( .A1(_04430_), .A2(_03039__PTR7), .ZN(_03039__PTR15) );
  AND2_X1 U18841 ( .A1(P2_P1_PhyAddrPointer_PTR5), .A2(P2_P1_PhyAddrPointer_PTR4), .ZN(_04411_) );
  AND2_X1 U18842 ( .A1(P2_P1_PhyAddrPointer_PTR7), .A2(P2_P1_PhyAddrPointer_PTR6), .ZN(_04412_) );
  AND2_X1 U18843 ( .A1(P2_P1_PhyAddrPointer_PTR9), .A2(P2_P1_PhyAddrPointer_PTR8), .ZN(_04413_) );
  AND2_X1 U18844 ( .A1(P2_P1_PhyAddrPointer_PTR11), .A2(P2_P1_PhyAddrPointer_PTR10), .ZN(_04414_) );
  AND2_X1 U18845 ( .A1(P2_P1_PhyAddrPointer_PTR13), .A2(P2_P1_PhyAddrPointer_PTR12), .ZN(_04415_) );
  AND2_X1 U18846 ( .A1(P2_P1_PhyAddrPointer_PTR15), .A2(P2_P1_PhyAddrPointer_PTR14), .ZN(_04416_) );
  AND2_X1 U18847 ( .A1(P2_P1_PhyAddrPointer_PTR17), .A2(P2_P1_PhyAddrPointer_PTR16), .ZN(_04417_) );
  AND2_X1 U18848 ( .A1(P2_P1_PhyAddrPointer_PTR19), .A2(P2_P1_PhyAddrPointer_PTR18), .ZN(_04418_) );
  AND2_X1 U18849 ( .A1(P2_P1_PhyAddrPointer_PTR21), .A2(P2_P1_PhyAddrPointer_PTR20), .ZN(_04419_) );
  AND2_X1 U18850 ( .A1(P2_P1_PhyAddrPointer_PTR23), .A2(P2_P1_PhyAddrPointer_PTR22), .ZN(_04420_) );
  AND2_X1 U18851 ( .A1(P2_P1_PhyAddrPointer_PTR25), .A2(P2_P1_PhyAddrPointer_PTR24), .ZN(_04421_) );
  AND2_X1 U18852 ( .A1(P2_P1_PhyAddrPointer_PTR27), .A2(P2_P1_PhyAddrPointer_PTR26), .ZN(_04422_) );
  AND2_X1 U18853 ( .A1(P2_P1_PhyAddrPointer_PTR29), .A2(P2_P1_PhyAddrPointer_PTR28), .ZN(_04423_) );
  AND2_X1 U18854 ( .A1(_04413_), .A2(_04412_), .ZN(_04424_) );
  AND2_X1 U18855 ( .A1(_04415_), .A2(_04414_), .ZN(_04425_) );
  AND2_X1 U18856 ( .A1(_04417_), .A2(_04416_), .ZN(_04426_) );
  AND2_X1 U18857 ( .A1(_04419_), .A2(_04418_), .ZN(_04427_) );
  AND2_X1 U18858 ( .A1(_04421_), .A2(_04420_), .ZN(_04428_) );
  AND2_X1 U18859 ( .A1(_04423_), .A2(_04422_), .ZN(_04429_) );
  AND2_X1 U18860 ( .A1(_04426_), .A2(_04425_), .ZN(_04430_) );
  AND2_X1 U18861 ( .A1(_04428_), .A2(_04427_), .ZN(_04431_) );
  AND2_X1 U18862 ( .A1(_04431_), .A2(_03039__PTR15), .ZN(_03039__PTR23) );
  AND2_X1 U18863 ( .A1(_04425_), .A2(_03039__PTR7), .ZN(_03039__PTR11) );
  AND2_X1 U18864 ( .A1(_04427_), .A2(_03039__PTR15), .ZN(_03039__PTR19) );
  AND2_X1 U18865 ( .A1(_04429_), .A2(_03039__PTR23), .ZN(_03039__PTR27) );
  AND2_X1 U18866 ( .A1(_04412_), .A2(_03039__PTR3), .ZN(_03039__PTR5) );
  AND2_X1 U18867 ( .A1(_04414_), .A2(_03039__PTR7), .ZN(_03039__PTR9) );
  AND2_X1 U18868 ( .A1(_04416_), .A2(_03039__PTR11), .ZN(_03039__PTR13) );
  AND2_X1 U18869 ( .A1(_04418_), .A2(_03039__PTR15), .ZN(_03039__PTR17) );
  AND2_X1 U18870 ( .A1(_04420_), .A2(_03039__PTR19), .ZN(_03039__PTR21) );
  AND2_X1 U18871 ( .A1(_04422_), .A2(_03039__PTR23), .ZN(_03039__PTR25) );
  AND2_X1 U18872 ( .A1(P2_P1_PhyAddrPointer_PTR4), .A2(_03039__PTR1), .ZN(_03039__PTR2) );
  AND2_X1 U18873 ( .A1(P2_P1_PhyAddrPointer_PTR6), .A2(_03039__PTR3), .ZN(_03039__PTR4) );
  AND2_X1 U18874 ( .A1(P2_P1_PhyAddrPointer_PTR8), .A2(_03039__PTR5), .ZN(_03039__PTR6) );
  AND2_X1 U18875 ( .A1(P2_P1_PhyAddrPointer_PTR10), .A2(_03039__PTR7), .ZN(_03039__PTR8) );
  AND2_X1 U18876 ( .A1(P2_P1_PhyAddrPointer_PTR12), .A2(_03039__PTR9), .ZN(_03039__PTR10) );
  AND2_X1 U18877 ( .A1(P2_P1_PhyAddrPointer_PTR14), .A2(_03039__PTR11), .ZN(_03039__PTR12) );
  AND2_X1 U18878 ( .A1(P2_P1_PhyAddrPointer_PTR16), .A2(_03039__PTR13), .ZN(_03039__PTR14) );
  AND2_X1 U18879 ( .A1(P2_P1_PhyAddrPointer_PTR18), .A2(_03039__PTR15), .ZN(_03039__PTR16) );
  AND2_X1 U18880 ( .A1(P2_P1_PhyAddrPointer_PTR20), .A2(_03039__PTR17), .ZN(_03039__PTR18) );
  AND2_X1 U18881 ( .A1(P2_P1_PhyAddrPointer_PTR22), .A2(_03039__PTR19), .ZN(_03039__PTR20) );
  AND2_X1 U18882 ( .A1(P2_P1_PhyAddrPointer_PTR24), .A2(_03039__PTR21), .ZN(_03039__PTR22) );
  AND2_X1 U18883 ( .A1(P2_P1_PhyAddrPointer_PTR26), .A2(_03039__PTR23), .ZN(_03039__PTR24) );
  AND2_X1 U18884 ( .A1(P2_P1_PhyAddrPointer_PTR28), .A2(_03039__PTR25), .ZN(_03039__PTR26) );
  AND2_X1 U18885 ( .A1(P2_P1_PhyAddrPointer_PTR30), .A2(_03039__PTR27), .ZN(_03039__PTR28) );
  AND2_X1 U18886 ( .A1(P2_P1_InstQueueWr_Addr_PTR1), .A2(P2_P1_InstQueueWr_Addr_PTR0), .ZN(_03024__PTR1) );
  AND2_X1 U18887 ( .A1(P2_P1_InstQueueWr_Addr_PTR2), .A2(_03024__PTR1), .ZN(_03024__PTR2) );
  AND2_X1 U18888 ( .A1(_02129__PTR1), .A2(_02129__PTR0), .ZN(_03025__PTR1) );
  AND2_X1 U18889 ( .A1(_02129__PTR2), .A2(_03025__PTR1), .ZN(_03025__PTR2) );
  AND2_X1 U18890 ( .A1(_02131__PTR1), .A2(P2_P1_InstQueueWr_Addr_PTR0), .ZN(_03030__PTR1) );
  AND2_X1 U18891 ( .A1(_02131__PTR2), .A2(_03030__PTR1), .ZN(_03030__PTR2) );
  AND2_X1 U18892 ( .A1(_02133__PTR1), .A2(_02129__PTR0), .ZN(_03035__PTR1) );
  AND2_X1 U18893 ( .A1(_02133__PTR2), .A2(_03035__PTR1), .ZN(_03035__PTR2) );
  AND2_X1 U18894 ( .A1(di2_PTR25), .A2(_03032__PTR0), .ZN(_03032__PTR1) );
  AND2_X1 U18895 ( .A1(_04388_), .A2(_03032__PTR1), .ZN(_03032__PTR3) );
  AND2_X1 U18896 ( .A1(di2_PTR27), .A2(di2_PTR26), .ZN(_04388_) );
  AND2_X1 U18897 ( .A1(di2_PTR29), .A2(di2_PTR28), .ZN(_04389_) );
  AND2_X1 U18898 ( .A1(_04389_), .A2(_03032__PTR3), .ZN(_03032__PTR5) );
  AND2_X1 U18899 ( .A1(di2_PTR26), .A2(_03032__PTR1), .ZN(_03032__PTR2) );
  AND2_X1 U18900 ( .A1(di2_PTR28), .A2(_03032__PTR3), .ZN(_03032__PTR4) );
  AND2_X1 U18901 ( .A1(di2_PTR30), .A2(_03032__PTR5), .ZN(_03032__PTR6) );
  AND2_X1 U18902 ( .A1(di2_PTR17), .A2(_03027__PTR0), .ZN(_03027__PTR1) );
  AND2_X1 U18903 ( .A1(_04386_), .A2(_03027__PTR1), .ZN(_03027__PTR3) );
  AND2_X1 U18904 ( .A1(di2_PTR19), .A2(di2_PTR18), .ZN(_04386_) );
  AND2_X1 U18905 ( .A1(di2_PTR21), .A2(di2_PTR20), .ZN(_04387_) );
  AND2_X1 U18906 ( .A1(_04387_), .A2(_03027__PTR3), .ZN(_03027__PTR5) );
  AND2_X1 U18907 ( .A1(di2_PTR18), .A2(_03027__PTR1), .ZN(_03027__PTR2) );
  AND2_X1 U18908 ( .A1(di2_PTR20), .A2(_03027__PTR3), .ZN(_03027__PTR4) );
  AND2_X1 U18909 ( .A1(di2_PTR22), .A2(_03027__PTR5), .ZN(_03027__PTR6) );
  AND2_X1 U18910 ( .A1(P2_rEIP_PTR2), .A2(_03023__PTR0), .ZN(_03023__PTR1) );
  AND2_X1 U18911 ( .A1(_04364_), .A2(_03023__PTR1), .ZN(_03023__PTR3) );
  AND2_X1 U18912 ( .A1(_04378_), .A2(_03023__PTR3), .ZN(_03023__PTR7) );
  AND2_X1 U18913 ( .A1(_04384_), .A2(_03023__PTR7), .ZN(_03023__PTR15) );
  AND2_X1 U18914 ( .A1(P2_rEIP_PTR8), .A2(P2_rEIP_PTR7), .ZN(_04366_) );
  AND2_X1 U18915 ( .A1(P2_rEIP_PTR16), .A2(P2_rEIP_PTR15), .ZN(_04370_) );
  AND2_X1 U18916 ( .A1(P2_rEIP_PTR20), .A2(P2_rEIP_PTR19), .ZN(_04372_) );
  AND2_X1 U18917 ( .A1(P2_rEIP_PTR28), .A2(P2_rEIP_PTR27), .ZN(_04376_) );
  AND2_X1 U18918 ( .A1(P2_rEIP_PTR30), .A2(P2_rEIP_PTR29), .ZN(_04377_) );
  AND2_X1 U18919 ( .A1(_04382_), .A2(_04381_), .ZN(_04385_) );
  AND2_X1 U18920 ( .A1(_04385_), .A2(_03023__PTR15), .ZN(_03023__PTR23) );
  AND2_X1 U18921 ( .A1(_04379_), .A2(_03023__PTR7), .ZN(_03023__PTR11) );
  AND2_X1 U18922 ( .A1(_04381_), .A2(_03023__PTR15), .ZN(_03023__PTR19) );
  AND2_X1 U18923 ( .A1(_04383_), .A2(_03023__PTR23), .ZN(_03023__PTR27) );
  AND2_X1 U18924 ( .A1(_04365_), .A2(_03023__PTR3), .ZN(_03023__PTR5) );
  AND2_X1 U18925 ( .A1(_04367_), .A2(_03023__PTR7), .ZN(_03023__PTR9) );
  AND2_X1 U18926 ( .A1(_04369_), .A2(_03023__PTR11), .ZN(_03023__PTR13) );
  AND2_X1 U18927 ( .A1(_04371_), .A2(_03023__PTR15), .ZN(_03023__PTR17) );
  AND2_X1 U18928 ( .A1(_04373_), .A2(_03023__PTR19), .ZN(_03023__PTR21) );
  AND2_X1 U18929 ( .A1(_04375_), .A2(_03023__PTR23), .ZN(_03023__PTR25) );
  AND2_X1 U18930 ( .A1(P2_rEIP_PTR3), .A2(_03023__PTR1), .ZN(_03023__PTR2) );
  AND2_X1 U18931 ( .A1(P2_rEIP_PTR5), .A2(_03023__PTR3), .ZN(_03023__PTR4) );
  AND2_X1 U18932 ( .A1(P2_rEIP_PTR7), .A2(_03023__PTR5), .ZN(_03023__PTR6) );
  AND2_X1 U18933 ( .A1(P2_rEIP_PTR9), .A2(_03023__PTR7), .ZN(_03023__PTR8) );
  AND2_X1 U18934 ( .A1(P2_rEIP_PTR11), .A2(_03023__PTR9), .ZN(_03023__PTR10) );
  AND2_X1 U18935 ( .A1(P2_rEIP_PTR13), .A2(_03023__PTR11), .ZN(_03023__PTR12) );
  AND2_X1 U18936 ( .A1(P2_rEIP_PTR15), .A2(_03023__PTR13), .ZN(_03023__PTR14) );
  AND2_X1 U18937 ( .A1(P2_rEIP_PTR17), .A2(_03023__PTR15), .ZN(_03023__PTR16) );
  AND2_X1 U18938 ( .A1(P2_rEIP_PTR19), .A2(_03023__PTR17), .ZN(_03023__PTR18) );
  AND2_X1 U18939 ( .A1(P2_rEIP_PTR21), .A2(_03023__PTR19), .ZN(_03023__PTR20) );
  AND2_X1 U18940 ( .A1(P2_rEIP_PTR23), .A2(_03023__PTR21), .ZN(_03023__PTR22) );
  AND2_X1 U18941 ( .A1(P2_rEIP_PTR25), .A2(_03023__PTR23), .ZN(_03023__PTR24) );
  AND2_X1 U18942 ( .A1(P2_rEIP_PTR27), .A2(_03023__PTR25), .ZN(_03023__PTR26) );
  AND2_X1 U18943 ( .A1(P2_rEIP_PTR29), .A2(_03023__PTR27), .ZN(_03023__PTR28) );
  AND2_X1 U18944 ( .A1(P2_rEIP_PTR3), .A2(_03038__PTR0), .ZN(_03038__PTR1) );
  AND2_X1 U18945 ( .A1(_04390_), .A2(_03038__PTR1), .ZN(_03038__PTR3) );
  AND2_X1 U18946 ( .A1(_04403_), .A2(_03038__PTR3), .ZN(_03038__PTR7) );
  AND2_X1 U18947 ( .A1(_04409_), .A2(_03038__PTR7), .ZN(_03038__PTR15) );
  AND2_X1 U18948 ( .A1(P2_rEIP_PTR5), .A2(P2_rEIP_PTR4), .ZN(_04390_) );
  AND2_X1 U18949 ( .A1(P2_rEIP_PTR7), .A2(P2_rEIP_PTR6), .ZN(_04391_) );
  AND2_X1 U18950 ( .A1(P2_rEIP_PTR9), .A2(P2_rEIP_PTR8), .ZN(_04392_) );
  AND2_X1 U18951 ( .A1(P2_rEIP_PTR11), .A2(P2_rEIP_PTR10), .ZN(_04393_) );
  AND2_X1 U18952 ( .A1(P2_rEIP_PTR13), .A2(P2_rEIP_PTR12), .ZN(_04394_) );
  AND2_X1 U18953 ( .A1(P2_rEIP_PTR15), .A2(P2_rEIP_PTR14), .ZN(_04395_) );
  AND2_X1 U18954 ( .A1(P2_rEIP_PTR17), .A2(P2_rEIP_PTR16), .ZN(_04396_) );
  AND2_X1 U18955 ( .A1(P2_rEIP_PTR19), .A2(P2_rEIP_PTR18), .ZN(_04397_) );
  AND2_X1 U18956 ( .A1(P2_rEIP_PTR21), .A2(P2_rEIP_PTR20), .ZN(_04398_) );
  AND2_X1 U18957 ( .A1(P2_rEIP_PTR23), .A2(P2_rEIP_PTR22), .ZN(_04399_) );
  AND2_X1 U18958 ( .A1(P2_rEIP_PTR25), .A2(P2_rEIP_PTR24), .ZN(_04400_) );
  AND2_X1 U18959 ( .A1(P2_rEIP_PTR27), .A2(P2_rEIP_PTR26), .ZN(_04401_) );
  AND2_X1 U18960 ( .A1(P2_rEIP_PTR29), .A2(P2_rEIP_PTR28), .ZN(_04402_) );
  AND2_X1 U18961 ( .A1(_04392_), .A2(_04391_), .ZN(_04403_) );
  AND2_X1 U18962 ( .A1(_04394_), .A2(_04393_), .ZN(_04404_) );
  AND2_X1 U18963 ( .A1(_04396_), .A2(_04395_), .ZN(_04405_) );
  AND2_X1 U18964 ( .A1(_04398_), .A2(_04397_), .ZN(_04406_) );
  AND2_X1 U18965 ( .A1(_04400_), .A2(_04399_), .ZN(_04407_) );
  AND2_X1 U18966 ( .A1(_04402_), .A2(_04401_), .ZN(_04408_) );
  AND2_X1 U18967 ( .A1(_04405_), .A2(_04404_), .ZN(_04409_) );
  AND2_X1 U18968 ( .A1(_04407_), .A2(_04406_), .ZN(_04410_) );
  AND2_X1 U18969 ( .A1(_04410_), .A2(_03038__PTR15), .ZN(_03038__PTR23) );
  AND2_X1 U18970 ( .A1(_04404_), .A2(_03038__PTR7), .ZN(_03038__PTR11) );
  AND2_X1 U18971 ( .A1(_04406_), .A2(_03038__PTR15), .ZN(_03038__PTR19) );
  AND2_X1 U18972 ( .A1(_04408_), .A2(_03038__PTR23), .ZN(_03038__PTR27) );
  AND2_X1 U18973 ( .A1(_04391_), .A2(_03038__PTR3), .ZN(_03038__PTR5) );
  AND2_X1 U18974 ( .A1(_04393_), .A2(_03038__PTR7), .ZN(_03038__PTR9) );
  AND2_X1 U18975 ( .A1(_04395_), .A2(_03038__PTR11), .ZN(_03038__PTR13) );
  AND2_X1 U18976 ( .A1(_04397_), .A2(_03038__PTR15), .ZN(_03038__PTR17) );
  AND2_X1 U18977 ( .A1(_04399_), .A2(_03038__PTR19), .ZN(_03038__PTR21) );
  AND2_X1 U18978 ( .A1(_04401_), .A2(_03038__PTR23), .ZN(_03038__PTR25) );
  AND2_X1 U18979 ( .A1(P2_rEIP_PTR4), .A2(_03038__PTR1), .ZN(_03038__PTR2) );
  AND2_X1 U18980 ( .A1(P2_rEIP_PTR6), .A2(_03038__PTR3), .ZN(_03038__PTR4) );
  AND2_X1 U18981 ( .A1(P2_rEIP_PTR8), .A2(_03038__PTR5), .ZN(_03038__PTR6) );
  AND2_X1 U18982 ( .A1(P2_rEIP_PTR10), .A2(_03038__PTR7), .ZN(_03038__PTR8) );
  AND2_X1 U18983 ( .A1(P2_rEIP_PTR12), .A2(_03038__PTR9), .ZN(_03038__PTR10) );
  AND2_X1 U18984 ( .A1(P2_rEIP_PTR14), .A2(_03038__PTR11), .ZN(_03038__PTR12) );
  AND2_X1 U18985 ( .A1(P2_rEIP_PTR16), .A2(_03038__PTR13), .ZN(_03038__PTR14) );
  AND2_X1 U18986 ( .A1(P2_rEIP_PTR18), .A2(_03038__PTR15), .ZN(_03038__PTR16) );
  AND2_X1 U18987 ( .A1(P2_rEIP_PTR20), .A2(_03038__PTR17), .ZN(_03038__PTR18) );
  AND2_X1 U18988 ( .A1(P2_rEIP_PTR22), .A2(_03038__PTR19), .ZN(_03038__PTR20) );
  AND2_X1 U18989 ( .A1(P2_rEIP_PTR24), .A2(_03038__PTR21), .ZN(_03038__PTR22) );
  AND2_X1 U18990 ( .A1(P2_rEIP_PTR26), .A2(_03038__PTR23), .ZN(_03038__PTR24) );
  AND2_X1 U18991 ( .A1(P2_rEIP_PTR28), .A2(_03038__PTR25), .ZN(_03038__PTR26) );
  AND2_X1 U18992 ( .A1(P2_rEIP_PTR30), .A2(_03038__PTR27), .ZN(_03038__PTR28) );
  AND2_X1 U18993 ( .A1(_03241__PTR4), .A2(_03240__PTR3), .ZN(_03243_) );
  OR2_X1 U18994 ( .A1(P3_P1_InstQueueRd_Addr_PTR4), .A2(_03243_), .ZN(_03240__PTR4) );
  AND2_X1 U18995 ( .A1(_02513__PTR59), .A2(_03236__PTR2), .ZN(_05005_) );
  AND2_X1 U18996 ( .A1(_03433__PTR4), .A2(_03434__PTR3), .ZN(_03237__PTR5) );
  OR2_X1 U18997 ( .A1(_05011_), .A2(_05008_), .ZN(_03434__PTR3) );
  AND2_X1 U18998 ( .A1(_03236__PTR1), .A2(_03236__PTR0), .ZN(_03238__PTR1) );
  AND2_X1 U18999 ( .A1(_03237__PTR5), .A2(_03236__PTR4), .ZN(_05006_) );
  AND2_X1 U19000 ( .A1(_05008_), .A2(_03238__PTR1), .ZN(_05007_) );
  AND2_X1 U19001 ( .A1(_02513__PTR59), .A2(_02513__PTR58), .ZN(_05008_) );
  AND2_X1 U19002 ( .A1(_03237__PTR5), .A2(_03239__PTR4), .ZN(_05009_) );
  AND2_X1 U19003 ( .A1(_05009_), .A2(_03238__PTR3), .ZN(_05010_) );
  OR2_X1 U19004 ( .A1(_03236__PTR3), .A2(_05005_), .ZN(_05011_) );
  OR2_X1 U19005 ( .A1(_05011_), .A2(_05007_), .ZN(_03238__PTR3) );
  OR2_X1 U19006 ( .A1(_05006_), .A2(_05010_), .ZN(_02475__PTR28) );
  AND2_X1 U19007 ( .A1(_03319__PTR1), .A2(P3_P1_InstAddrPointer_PTR0), .ZN(_03320__PTR1) );
  AND2_X1 U19008 ( .A1(_03235__PTR9), .A2(_03235__PTR8), .ZN(_04957_) );
  AND2_X1 U19009 ( .A1(_03235__PTR19), .A2(_03235__PTR18), .ZN(_04962_) );
  AND2_X1 U19010 ( .A1(_04973_), .A2(_04972_), .ZN(_04977_) );
  AND2_X1 U19011 ( .A1(_04975_), .A2(_04974_), .ZN(_04978_) );
  AND2_X1 U19012 ( .A1(_03235__PTR3), .A2(P3_P1_InstAddrPointer_PTR2), .ZN(_04925_) );
  AND2_X1 U19013 ( .A1(_03235__PTR5), .A2(P3_P1_InstAddrPointer_PTR4), .ZN(_04926_) );
  AND2_X1 U19014 ( .A1(_03235__PTR7), .A2(P3_P1_InstAddrPointer_PTR6), .ZN(_04927_) );
  AND2_X1 U19015 ( .A1(_03235__PTR9), .A2(P3_P1_InstAddrPointer_PTR8), .ZN(_04928_) );
  AND2_X1 U19016 ( .A1(_03235__PTR11), .A2(P3_P1_InstAddrPointer_PTR10), .ZN(_04929_) );
  AND2_X1 U19017 ( .A1(_03235__PTR13), .A2(P3_P1_InstAddrPointer_PTR12), .ZN(_04930_) );
  AND2_X1 U19018 ( .A1(_03235__PTR15), .A2(P3_P1_InstAddrPointer_PTR14), .ZN(_04931_) );
  AND2_X1 U19019 ( .A1(_03235__PTR17), .A2(P3_P1_InstAddrPointer_PTR16), .ZN(_04932_) );
  AND2_X1 U19020 ( .A1(_03235__PTR19), .A2(P3_P1_InstAddrPointer_PTR18), .ZN(_04933_) );
  AND2_X1 U19021 ( .A1(_03235__PTR21), .A2(P3_P1_InstAddrPointer_PTR20), .ZN(_04934_) );
  AND2_X1 U19022 ( .A1(_03235__PTR23), .A2(P3_P1_InstAddrPointer_PTR22), .ZN(_04935_) );
  AND2_X1 U19023 ( .A1(_03235__PTR25), .A2(P3_P1_InstAddrPointer_PTR24), .ZN(_04936_) );
  AND2_X1 U19024 ( .A1(_03235__PTR27), .A2(P3_P1_InstAddrPointer_PTR26), .ZN(_04937_) );
  AND2_X1 U19025 ( .A1(_03235__PTR29), .A2(P3_P1_InstAddrPointer_PTR28), .ZN(_04938_) );
  AND2_X1 U19026 ( .A1(_03233__PTR31), .A2(P3_P1_InstAddrPointer_PTR30), .ZN(_04939_) );
  AND2_X1 U19027 ( .A1(_04956_), .A2(_04981_), .ZN(_04941_) );
  AND2_X1 U19028 ( .A1(_04958_), .A2(_04983_), .ZN(_04942_) );
  AND2_X1 U19029 ( .A1(_04960_), .A2(_04985_), .ZN(_04943_) );
  AND2_X1 U19030 ( .A1(_04962_), .A2(_04987_), .ZN(_04944_) );
  AND2_X1 U19031 ( .A1(_04964_), .A2(_04989_), .ZN(_04945_) );
  AND2_X1 U19032 ( .A1(_04966_), .A2(_04991_), .ZN(_04946_) );
  AND2_X1 U19033 ( .A1(_04968_), .A2(_04993_), .ZN(_04947_) );
  AND2_X1 U19034 ( .A1(_04969_), .A2(_03234__PTR3), .ZN(_04948_) );
  AND2_X1 U19035 ( .A1(_04971_), .A2(_04995_), .ZN(_04949_) );
  AND2_X1 U19036 ( .A1(_04973_), .A2(_04997_), .ZN(_04950_) );
  AND2_X1 U19037 ( .A1(_04975_), .A2(_04999_), .ZN(_04951_) );
  AND2_X1 U19038 ( .A1(_04976_), .A2(_03234__PTR7), .ZN(_04952_) );
  AND2_X1 U19039 ( .A1(_04978_), .A2(_05002_), .ZN(_04953_) );
  AND2_X1 U19040 ( .A1(_04979_), .A2(_03234__PTR15), .ZN(_04954_) );
  AND2_X1 U19041 ( .A1(_03235__PTR3), .A2(_03235__PTR2), .ZN(_04940_) );
  AND2_X1 U19042 ( .A1(_03235__PTR5), .A2(_03235__PTR4), .ZN(_04955_) );
  AND2_X1 U19043 ( .A1(_03235__PTR7), .A2(_03235__PTR6), .ZN(_04956_) );
  AND2_X1 U19044 ( .A1(_03235__PTR11), .A2(_03235__PTR10), .ZN(_04958_) );
  AND2_X1 U19045 ( .A1(_03235__PTR13), .A2(_03235__PTR12), .ZN(_04959_) );
  AND2_X1 U19046 ( .A1(_03235__PTR15), .A2(_03235__PTR14), .ZN(_04960_) );
  AND2_X1 U19047 ( .A1(_03235__PTR17), .A2(_03235__PTR16), .ZN(_04961_) );
  AND2_X1 U19048 ( .A1(_03235__PTR21), .A2(_03235__PTR20), .ZN(_04963_) );
  AND2_X1 U19049 ( .A1(_03235__PTR23), .A2(_03235__PTR22), .ZN(_04964_) );
  AND2_X1 U19050 ( .A1(_03235__PTR25), .A2(_03235__PTR24), .ZN(_04965_) );
  AND2_X1 U19051 ( .A1(_03235__PTR27), .A2(_03235__PTR26), .ZN(_04966_) );
  AND2_X1 U19052 ( .A1(_03235__PTR29), .A2(_03235__PTR28), .ZN(_04967_) );
  AND2_X1 U19053 ( .A1(_03233__PTR31), .A2(_03235__PTR30), .ZN(_04968_) );
  AND2_X1 U19054 ( .A1(_04956_), .A2(_04955_), .ZN(_04969_) );
  AND2_X1 U19055 ( .A1(_04958_), .A2(_04957_), .ZN(_04970_) );
  AND2_X1 U19056 ( .A1(_04960_), .A2(_04959_), .ZN(_04971_) );
  AND2_X1 U19057 ( .A1(_04962_), .A2(_04961_), .ZN(_04972_) );
  AND2_X1 U19058 ( .A1(_04964_), .A2(_04963_), .ZN(_04973_) );
  AND2_X1 U19059 ( .A1(_04966_), .A2(_04965_), .ZN(_04974_) );
  AND2_X1 U19060 ( .A1(_04968_), .A2(_04967_), .ZN(_04975_) );
  AND2_X1 U19061 ( .A1(_04971_), .A2(_04970_), .ZN(_04976_) );
  AND2_X1 U19062 ( .A1(_04978_), .A2(_04977_), .ZN(_04979_) );
  OR2_X1 U19063 ( .A1(P3_P1_InstAddrPointer_PTR3), .A2(_04925_), .ZN(_04980_) );
  OR2_X1 U19064 ( .A1(P3_P1_InstAddrPointer_PTR5), .A2(_04926_), .ZN(_04981_) );
  OR2_X1 U19065 ( .A1(P3_P1_InstAddrPointer_PTR7), .A2(_04927_), .ZN(_04982_) );
  OR2_X1 U19066 ( .A1(P3_P1_InstAddrPointer_PTR9), .A2(_04928_), .ZN(_04983_) );
  OR2_X1 U19067 ( .A1(P3_P1_InstAddrPointer_PTR11), .A2(_04929_), .ZN(_04984_) );
  OR2_X1 U19068 ( .A1(P3_P1_InstAddrPointer_PTR13), .A2(_04930_), .ZN(_04985_) );
  OR2_X1 U19069 ( .A1(P3_P1_InstAddrPointer_PTR15), .A2(_04931_), .ZN(_04986_) );
  OR2_X1 U19070 ( .A1(P3_P1_InstAddrPointer_PTR17), .A2(_04932_), .ZN(_04987_) );
  OR2_X1 U19071 ( .A1(P3_P1_InstAddrPointer_PTR19), .A2(_04933_), .ZN(_04988_) );
  OR2_X1 U19072 ( .A1(P3_P1_InstAddrPointer_PTR21), .A2(_04934_), .ZN(_04989_) );
  OR2_X1 U19073 ( .A1(P3_P1_InstAddrPointer_PTR23), .A2(_04935_), .ZN(_04990_) );
  OR2_X1 U19074 ( .A1(P3_P1_InstAddrPointer_PTR25), .A2(_04936_), .ZN(_04991_) );
  OR2_X1 U19075 ( .A1(P3_P1_InstAddrPointer_PTR27), .A2(_04937_), .ZN(_04992_) );
  OR2_X1 U19076 ( .A1(P3_P1_InstAddrPointer_PTR29), .A2(_04938_), .ZN(_04993_) );
  OR2_X1 U19077 ( .A1(_04980_), .A2(_04940_), .ZN(_03234__PTR3) );
  OR2_X1 U19078 ( .A1(_04982_), .A2(_04941_), .ZN(_04994_) );
  OR2_X1 U19079 ( .A1(_04984_), .A2(_04942_), .ZN(_04995_) );
  OR2_X1 U19080 ( .A1(_04986_), .A2(_04943_), .ZN(_04996_) );
  OR2_X1 U19081 ( .A1(_04988_), .A2(_04944_), .ZN(_04997_) );
  OR2_X1 U19082 ( .A1(_04990_), .A2(_04945_), .ZN(_04998_) );
  OR2_X1 U19083 ( .A1(_04992_), .A2(_04946_), .ZN(_04999_) );
  OR2_X1 U19084 ( .A1(_04939_), .A2(_04947_), .ZN(_05000_) );
  OR2_X1 U19085 ( .A1(_04994_), .A2(_04948_), .ZN(_03234__PTR7) );
  OR2_X1 U19086 ( .A1(_04996_), .A2(_04949_), .ZN(_05001_) );
  OR2_X1 U19087 ( .A1(_04998_), .A2(_04950_), .ZN(_05002_) );
  OR2_X1 U19088 ( .A1(_05000_), .A2(_04951_), .ZN(_05003_) );
  OR2_X1 U19089 ( .A1(_05001_), .A2(_04952_), .ZN(_03234__PTR15) );
  OR2_X1 U19090 ( .A1(_05003_), .A2(_04953_), .ZN(_05004_) );
  OR2_X1 U19091 ( .A1(_05004_), .A2(_04954_), .ZN(_03234__PTR31) );
  AND2_X1 U19092 ( .A1(_02513__PTR43), .A2(_02513__PTR42), .ZN(_05383_) );
  AND2_X1 U19093 ( .A1(_03431__PTR4), .A2(_03432__PTR3), .ZN(_03230__PTR5) );
  OR2_X1 U19094 ( .A1(_03231__PTR3), .A2(_05383_), .ZN(_03432__PTR3) );
  AND2_X1 U19095 ( .A1(_03230__PTR5), .A2(_03229__PTR4), .ZN(_04921_) );
  AND2_X1 U19096 ( .A1(_02513__PTR43), .A2(_03229__PTR2), .ZN(_04922_) );
  AND2_X1 U19097 ( .A1(_03230__PTR5), .A2(_03232__PTR4), .ZN(_04923_) );
  AND2_X1 U19098 ( .A1(_04923_), .A2(_03231__PTR3), .ZN(_04924_) );
  OR2_X1 U19099 ( .A1(_03229__PTR3), .A2(_04922_), .ZN(_03231__PTR3) );
  OR2_X1 U19100 ( .A1(_04921_), .A2(_04924_), .ZN(_03231__PTR5) );
  AND2_X1 U19101 ( .A1(_03227__PTR1), .A2(_03226__PTR0), .ZN(_04915_) );
  AND2_X1 U19102 ( .A1(_03227__PTR3), .A2(_03228__PTR2), .ZN(_04916_) );
  AND2_X1 U19103 ( .A1(_04918_), .A2(_03226__PTR1), .ZN(_04917_) );
  AND2_X1 U19104 ( .A1(_03227__PTR3), .A2(_03227__PTR2), .ZN(_04918_) );
  AND2_X1 U19105 ( .A1(_03227__PTR4), .A2(_03226__PTR3), .ZN(_04919_) );
  OR2_X1 U19106 ( .A1(_03228__PTR0), .A2(_03227__PTR0), .ZN(_03226__PTR0) );
  OR2_X1 U19107 ( .A1(_03228__PTR1), .A2(_04915_), .ZN(_03226__PTR1) );
  OR2_X1 U19108 ( .A1(_03228__PTR3), .A2(_04916_), .ZN(_04920_) );
  OR2_X1 U19109 ( .A1(_04920_), .A2(_04917_), .ZN(_03226__PTR3) );
  OR2_X1 U19110 ( .A1(_03228__PTR4), .A2(_04919_), .ZN(_03226__PTR4) );
  AND2_X1 U19111 ( .A1(P3_EBX_PTR1), .A2(P3_EBX_PTR0), .ZN(_03318__PTR1) );
  AND2_X1 U19112 ( .A1(_05251_), .A2(_03318__PTR1), .ZN(_03318__PTR3) );
  AND2_X1 U19113 ( .A1(_05265_), .A2(_03318__PTR3), .ZN(_03318__PTR7) );
  AND2_X1 U19114 ( .A1(_05271_), .A2(_03318__PTR7), .ZN(_03318__PTR15) );
  AND2_X1 U19115 ( .A1(P3_EBX_PTR3), .A2(P3_EBX_PTR2), .ZN(_05251_) );
  AND2_X1 U19116 ( .A1(P3_EBX_PTR5), .A2(P3_EBX_PTR4), .ZN(_05252_) );
  AND2_X1 U19117 ( .A1(P3_EBX_PTR7), .A2(P3_EBX_PTR6), .ZN(_05253_) );
  AND2_X1 U19118 ( .A1(P3_EBX_PTR9), .A2(P3_EBX_PTR8), .ZN(_05254_) );
  AND2_X1 U19119 ( .A1(P3_EBX_PTR11), .A2(P3_EBX_PTR10), .ZN(_05255_) );
  AND2_X1 U19120 ( .A1(P3_EBX_PTR13), .A2(P3_EBX_PTR12), .ZN(_05256_) );
  AND2_X1 U19121 ( .A1(P3_EBX_PTR15), .A2(P3_EBX_PTR14), .ZN(_05257_) );
  AND2_X1 U19122 ( .A1(P3_EBX_PTR17), .A2(P3_EBX_PTR16), .ZN(_05258_) );
  AND2_X1 U19123 ( .A1(P3_EBX_PTR19), .A2(P3_EBX_PTR18), .ZN(_05259_) );
  AND2_X1 U19124 ( .A1(P3_EBX_PTR21), .A2(P3_EBX_PTR20), .ZN(_05260_) );
  AND2_X1 U19125 ( .A1(P3_EBX_PTR23), .A2(P3_EBX_PTR22), .ZN(_05261_) );
  AND2_X1 U19126 ( .A1(P3_EBX_PTR25), .A2(P3_EBX_PTR24), .ZN(_05262_) );
  AND2_X1 U19127 ( .A1(P3_EBX_PTR27), .A2(P3_EBX_PTR26), .ZN(_05263_) );
  AND2_X1 U19128 ( .A1(P3_EBX_PTR29), .A2(P3_EBX_PTR28), .ZN(_05264_) );
  AND2_X1 U19129 ( .A1(_05253_), .A2(_05252_), .ZN(_05265_) );
  AND2_X1 U19130 ( .A1(_05255_), .A2(_05254_), .ZN(_05266_) );
  AND2_X1 U19131 ( .A1(_05257_), .A2(_05256_), .ZN(_05267_) );
  AND2_X1 U19132 ( .A1(_05259_), .A2(_05258_), .ZN(_05268_) );
  AND2_X1 U19133 ( .A1(_05261_), .A2(_05260_), .ZN(_05269_) );
  AND2_X1 U19134 ( .A1(_05263_), .A2(_05262_), .ZN(_05270_) );
  AND2_X1 U19135 ( .A1(_05267_), .A2(_05266_), .ZN(_05271_) );
  AND2_X1 U19136 ( .A1(_05269_), .A2(_05268_), .ZN(_05272_) );
  AND2_X1 U19137 ( .A1(_05272_), .A2(_03318__PTR15), .ZN(_03318__PTR23) );
  AND2_X1 U19138 ( .A1(_05266_), .A2(_03318__PTR7), .ZN(_03318__PTR11) );
  AND2_X1 U19139 ( .A1(_05268_), .A2(_03318__PTR15), .ZN(_03318__PTR19) );
  AND2_X1 U19140 ( .A1(_05270_), .A2(_03318__PTR23), .ZN(_03318__PTR27) );
  AND2_X1 U19141 ( .A1(_05252_), .A2(_03318__PTR3), .ZN(_03318__PTR5) );
  AND2_X1 U19142 ( .A1(_05254_), .A2(_03318__PTR7), .ZN(_03318__PTR9) );
  AND2_X1 U19143 ( .A1(_05256_), .A2(_03318__PTR11), .ZN(_03318__PTR13) );
  AND2_X1 U19144 ( .A1(_05258_), .A2(_03318__PTR15), .ZN(_03318__PTR17) );
  AND2_X1 U19145 ( .A1(_05260_), .A2(_03318__PTR19), .ZN(_03318__PTR21) );
  AND2_X1 U19146 ( .A1(_05262_), .A2(_03318__PTR23), .ZN(_03318__PTR25) );
  AND2_X1 U19147 ( .A1(_05264_), .A2(_03318__PTR27), .ZN(_03318__PTR29) );
  AND2_X1 U19148 ( .A1(P3_EBX_PTR2), .A2(_03318__PTR1), .ZN(_03318__PTR2) );
  AND2_X1 U19149 ( .A1(P3_EBX_PTR4), .A2(_03318__PTR3), .ZN(_03318__PTR4) );
  AND2_X1 U19150 ( .A1(P3_EBX_PTR6), .A2(_03318__PTR5), .ZN(_03318__PTR6) );
  AND2_X1 U19151 ( .A1(P3_EBX_PTR8), .A2(_03318__PTR7), .ZN(_03318__PTR8) );
  AND2_X1 U19152 ( .A1(P3_EBX_PTR10), .A2(_03318__PTR9), .ZN(_03318__PTR10) );
  AND2_X1 U19153 ( .A1(P3_EBX_PTR12), .A2(_03318__PTR11), .ZN(_03318__PTR12) );
  AND2_X1 U19154 ( .A1(P3_EBX_PTR14), .A2(_03318__PTR13), .ZN(_03318__PTR14) );
  AND2_X1 U19155 ( .A1(P3_EBX_PTR16), .A2(_03318__PTR15), .ZN(_03318__PTR16) );
  AND2_X1 U19156 ( .A1(P3_EBX_PTR18), .A2(_03318__PTR17), .ZN(_03318__PTR18) );
  AND2_X1 U19157 ( .A1(P3_EBX_PTR20), .A2(_03318__PTR19), .ZN(_03318__PTR20) );
  AND2_X1 U19158 ( .A1(P3_EBX_PTR22), .A2(_03318__PTR21), .ZN(_03318__PTR22) );
  AND2_X1 U19159 ( .A1(P3_EBX_PTR24), .A2(_03318__PTR23), .ZN(_03318__PTR24) );
  AND2_X1 U19160 ( .A1(P3_EBX_PTR26), .A2(_03318__PTR25), .ZN(_03318__PTR26) );
  AND2_X1 U19161 ( .A1(P3_EBX_PTR28), .A2(_03318__PTR27), .ZN(_03318__PTR28) );
  AND2_X1 U19162 ( .A1(P3_EBX_PTR30), .A2(_03318__PTR29), .ZN(_03318__PTR30) );
  AND2_X1 U19163 ( .A1(P3_EAX_PTR1), .A2(P3_EAX_PTR0), .ZN(_03317__PTR1) );
  AND2_X1 U19164 ( .A1(_05237_), .A2(_03317__PTR1), .ZN(_03317__PTR3) );
  AND2_X1 U19165 ( .A1(_05245_), .A2(_03317__PTR3), .ZN(_03317__PTR7) );
  AND2_X1 U19166 ( .A1(_05249_), .A2(_03317__PTR7), .ZN(_03317__PTR15) );
  AND2_X1 U19167 ( .A1(P3_EAX_PTR3), .A2(P3_EAX_PTR2), .ZN(_05237_) );
  AND2_X1 U19168 ( .A1(P3_EAX_PTR5), .A2(P3_EAX_PTR4), .ZN(_05238_) );
  AND2_X1 U19169 ( .A1(P3_EAX_PTR7), .A2(P3_EAX_PTR6), .ZN(_05239_) );
  AND2_X1 U19170 ( .A1(P3_EAX_PTR9), .A2(P3_EAX_PTR8), .ZN(_05240_) );
  AND2_X1 U19171 ( .A1(P3_EAX_PTR11), .A2(P3_EAX_PTR10), .ZN(_05241_) );
  AND2_X1 U19172 ( .A1(P3_EAX_PTR13), .A2(P3_EAX_PTR12), .ZN(_05242_) );
  AND2_X1 U19173 ( .A1(P3_EAX_PTR15), .A2(P3_EAX_PTR14), .ZN(_05243_) );
  AND2_X1 U19174 ( .A1(P3_EAX_PTR17), .A2(P3_EAX_PTR16), .ZN(_05244_) );
  AND2_X1 U19175 ( .A1(P3_EAX_PTR23), .A2(P3_EAX_PTR22), .ZN(_05231_) );
  AND2_X1 U19176 ( .A1(P3_EAX_PTR25), .A2(P3_EAX_PTR24), .ZN(_05232_) );
  AND2_X1 U19177 ( .A1(P3_EAX_PTR27), .A2(P3_EAX_PTR26), .ZN(_05233_) );
  AND2_X1 U19178 ( .A1(P3_EAX_PTR29), .A2(P3_EAX_PTR28), .ZN(_05234_) );
  AND2_X1 U19179 ( .A1(_05239_), .A2(_05238_), .ZN(_05245_) );
  AND2_X1 U19180 ( .A1(_05241_), .A2(_05240_), .ZN(_05246_) );
  AND2_X1 U19181 ( .A1(_05243_), .A2(_05242_), .ZN(_05247_) );
  AND2_X1 U19182 ( .A1(_05229_), .A2(_05244_), .ZN(_05248_) );
  AND2_X1 U19183 ( .A1(_05231_), .A2(_05230_), .ZN(_05235_) );
  AND2_X1 U19184 ( .A1(_05233_), .A2(_05232_), .ZN(_05236_) );
  AND2_X1 U19185 ( .A1(_05247_), .A2(_05246_), .ZN(_05249_) );
  AND2_X1 U19186 ( .A1(_05235_), .A2(_05248_), .ZN(_05250_) );
  AND2_X1 U19187 ( .A1(_05250_), .A2(_03317__PTR15), .ZN(_03317__PTR23) );
  AND2_X1 U19188 ( .A1(_05246_), .A2(_03317__PTR7), .ZN(_03317__PTR11) );
  AND2_X1 U19189 ( .A1(_05248_), .A2(_03317__PTR15), .ZN(_03317__PTR19) );
  AND2_X1 U19190 ( .A1(_05236_), .A2(_03317__PTR23), .ZN(_03317__PTR27) );
  AND2_X1 U19191 ( .A1(_05238_), .A2(_03317__PTR3), .ZN(_03317__PTR5) );
  AND2_X1 U19192 ( .A1(_05240_), .A2(_03317__PTR7), .ZN(_03317__PTR9) );
  AND2_X1 U19193 ( .A1(_05242_), .A2(_03317__PTR11), .ZN(_03317__PTR13) );
  AND2_X1 U19194 ( .A1(_05244_), .A2(_03317__PTR15), .ZN(_03317__PTR17) );
  AND2_X1 U19195 ( .A1(_05230_), .A2(_03317__PTR19), .ZN(_03317__PTR21) );
  AND2_X1 U19196 ( .A1(_05232_), .A2(_03317__PTR23), .ZN(_03317__PTR25) );
  AND2_X1 U19197 ( .A1(_05234_), .A2(_03317__PTR27), .ZN(_03317__PTR29) );
  AND2_X1 U19198 ( .A1(P3_EAX_PTR2), .A2(_03317__PTR1), .ZN(_03317__PTR2) );
  AND2_X1 U19199 ( .A1(P3_EAX_PTR4), .A2(_03317__PTR3), .ZN(_03317__PTR4) );
  AND2_X1 U19200 ( .A1(P3_EAX_PTR6), .A2(_03317__PTR5), .ZN(_03317__PTR6) );
  AND2_X1 U19201 ( .A1(P3_EAX_PTR8), .A2(_03317__PTR7), .ZN(_03317__PTR8) );
  AND2_X1 U19202 ( .A1(P3_EAX_PTR10), .A2(_03317__PTR9), .ZN(_03317__PTR10) );
  AND2_X1 U19203 ( .A1(P3_EAX_PTR12), .A2(_03317__PTR11), .ZN(_03317__PTR12) );
  AND2_X1 U19204 ( .A1(P3_EAX_PTR14), .A2(_03317__PTR13), .ZN(_03317__PTR14) );
  AND2_X1 U19205 ( .A1(P3_EAX_PTR16), .A2(_03317__PTR15), .ZN(_03317__PTR16) );
  AND2_X1 U19206 ( .A1(P3_EAX_PTR18), .A2(_03317__PTR17), .ZN(_03317__PTR18) );
  AND2_X1 U19207 ( .A1(P3_EAX_PTR20), .A2(_03317__PTR19), .ZN(_03317__PTR20) );
  AND2_X1 U19208 ( .A1(P3_EAX_PTR22), .A2(_03317__PTR21), .ZN(_03317__PTR22) );
  AND2_X1 U19209 ( .A1(P3_EAX_PTR24), .A2(_03317__PTR23), .ZN(_03317__PTR24) );
  AND2_X1 U19210 ( .A1(P3_EAX_PTR26), .A2(_03317__PTR25), .ZN(_03317__PTR26) );
  AND2_X1 U19211 ( .A1(P3_EAX_PTR28), .A2(_03317__PTR27), .ZN(_03317__PTR28) );
  AND2_X1 U19212 ( .A1(P3_EAX_PTR30), .A2(_03317__PTR29), .ZN(_03317__PTR30) );
  AND2_X1 U19213 ( .A1(P3_EAX_PTR17), .A2(_03314__PTR0), .ZN(_03314__PTR1) );
  AND2_X1 U19214 ( .A1(_05229_), .A2(_03314__PTR1), .ZN(_03314__PTR3) );
  AND2_X1 U19215 ( .A1(_05235_), .A2(_03314__PTR3), .ZN(_03314__PTR7) );
  AND2_X1 U19216 ( .A1(P3_EAX_PTR19), .A2(P3_EAX_PTR18), .ZN(_05229_) );
  AND2_X1 U19217 ( .A1(P3_EAX_PTR21), .A2(P3_EAX_PTR20), .ZN(_05230_) );
  AND2_X1 U19218 ( .A1(_05236_), .A2(_03314__PTR7), .ZN(_03314__PTR11) );
  AND2_X1 U19219 ( .A1(_05230_), .A2(_03314__PTR3), .ZN(_03314__PTR5) );
  AND2_X1 U19220 ( .A1(_05232_), .A2(_03314__PTR7), .ZN(_03314__PTR9) );
  AND2_X1 U19221 ( .A1(_05234_), .A2(_03314__PTR11), .ZN(_03314__PTR13) );
  AND2_X1 U19222 ( .A1(P3_EAX_PTR18), .A2(_03314__PTR1), .ZN(_03314__PTR2) );
  AND2_X1 U19223 ( .A1(P3_EAX_PTR20), .A2(_03314__PTR3), .ZN(_03314__PTR4) );
  AND2_X1 U19224 ( .A1(P3_EAX_PTR22), .A2(_03314__PTR5), .ZN(_03314__PTR6) );
  AND2_X1 U19225 ( .A1(P3_EAX_PTR24), .A2(_03314__PTR7), .ZN(_03314__PTR8) );
  AND2_X1 U19226 ( .A1(P3_EAX_PTR26), .A2(_03314__PTR9), .ZN(_03314__PTR10) );
  AND2_X1 U19227 ( .A1(P3_EAX_PTR28), .A2(_03314__PTR11), .ZN(_03314__PTR12) );
  AND2_X1 U19228 ( .A1(P3_rEIP_PTR2), .A2(P3_rEIP_PTR1), .ZN(_03311__PTR1) );
  AND2_X1 U19229 ( .A1(_05012_), .A2(_03311__PTR1), .ZN(_03311__PTR3) );
  AND2_X1 U19230 ( .A1(_05026_), .A2(_03311__PTR3), .ZN(_03311__PTR7) );
  AND2_X1 U19231 ( .A1(_05032_), .A2(_03311__PTR7), .ZN(_03311__PTR15) );
  AND2_X1 U19232 ( .A1(P3_rEIP_PTR4), .A2(P3_rEIP_PTR3), .ZN(_05012_) );
  AND2_X1 U19233 ( .A1(P3_rEIP_PTR6), .A2(P3_rEIP_PTR5), .ZN(_05013_) );
  AND2_X1 U19234 ( .A1(P3_rEIP_PTR8), .A2(P3_rEIP_PTR7), .ZN(_05014_) );
  AND2_X1 U19235 ( .A1(P3_rEIP_PTR10), .A2(P3_rEIP_PTR9), .ZN(_05015_) );
  AND2_X1 U19236 ( .A1(P3_rEIP_PTR12), .A2(P3_rEIP_PTR11), .ZN(_05016_) );
  AND2_X1 U19237 ( .A1(P3_rEIP_PTR14), .A2(P3_rEIP_PTR13), .ZN(_05017_) );
  AND2_X1 U19238 ( .A1(P3_rEIP_PTR16), .A2(P3_rEIP_PTR15), .ZN(_05018_) );
  AND2_X1 U19239 ( .A1(P3_rEIP_PTR18), .A2(P3_rEIP_PTR17), .ZN(_05019_) );
  AND2_X1 U19240 ( .A1(P3_rEIP_PTR20), .A2(P3_rEIP_PTR19), .ZN(_05020_) );
  AND2_X1 U19241 ( .A1(P3_rEIP_PTR22), .A2(P3_rEIP_PTR21), .ZN(_05021_) );
  AND2_X1 U19242 ( .A1(P3_rEIP_PTR24), .A2(P3_rEIP_PTR23), .ZN(_05022_) );
  AND2_X1 U19243 ( .A1(P3_rEIP_PTR26), .A2(P3_rEIP_PTR25), .ZN(_05023_) );
  AND2_X1 U19244 ( .A1(P3_rEIP_PTR28), .A2(P3_rEIP_PTR27), .ZN(_05024_) );
  AND2_X1 U19245 ( .A1(P3_rEIP_PTR30), .A2(P3_rEIP_PTR29), .ZN(_05025_) );
  AND2_X1 U19246 ( .A1(_05014_), .A2(_05013_), .ZN(_05026_) );
  AND2_X1 U19247 ( .A1(_05016_), .A2(_05015_), .ZN(_05027_) );
  AND2_X1 U19248 ( .A1(_05018_), .A2(_05017_), .ZN(_05028_) );
  AND2_X1 U19249 ( .A1(_05020_), .A2(_05019_), .ZN(_05029_) );
  AND2_X1 U19250 ( .A1(_05022_), .A2(_05021_), .ZN(_05030_) );
  AND2_X1 U19251 ( .A1(_05024_), .A2(_05023_), .ZN(_05031_) );
  AND2_X1 U19252 ( .A1(_05028_), .A2(_05027_), .ZN(_05032_) );
  AND2_X1 U19253 ( .A1(_05030_), .A2(_05029_), .ZN(_05033_) );
  AND2_X1 U19254 ( .A1(_05033_), .A2(_03311__PTR15), .ZN(_03311__PTR23) );
  AND2_X1 U19255 ( .A1(_05027_), .A2(_03311__PTR7), .ZN(_03311__PTR11) );
  AND2_X1 U19256 ( .A1(_05029_), .A2(_03311__PTR15), .ZN(_03311__PTR19) );
  AND2_X1 U19257 ( .A1(_05031_), .A2(_03311__PTR23), .ZN(_03311__PTR27) );
  AND2_X1 U19258 ( .A1(_05013_), .A2(_03311__PTR3), .ZN(_03311__PTR5) );
  AND2_X1 U19259 ( .A1(_05015_), .A2(_03311__PTR7), .ZN(_03311__PTR9) );
  AND2_X1 U19260 ( .A1(_05017_), .A2(_03311__PTR11), .ZN(_03311__PTR13) );
  AND2_X1 U19261 ( .A1(_05019_), .A2(_03311__PTR15), .ZN(_03311__PTR17) );
  AND2_X1 U19262 ( .A1(_05021_), .A2(_03311__PTR19), .ZN(_03311__PTR21) );
  AND2_X1 U19263 ( .A1(_05023_), .A2(_03311__PTR23), .ZN(_03311__PTR25) );
  AND2_X1 U19264 ( .A1(_05025_), .A2(_03311__PTR27), .ZN(_03311__PTR29) );
  AND2_X1 U19265 ( .A1(P3_rEIP_PTR3), .A2(_03311__PTR1), .ZN(_03311__PTR2) );
  AND2_X1 U19266 ( .A1(P3_rEIP_PTR5), .A2(_03311__PTR3), .ZN(_03311__PTR4) );
  AND2_X1 U19267 ( .A1(P3_rEIP_PTR7), .A2(_03311__PTR5), .ZN(_03311__PTR6) );
  AND2_X1 U19268 ( .A1(P3_rEIP_PTR9), .A2(_03311__PTR7), .ZN(_03311__PTR8) );
  AND2_X1 U19269 ( .A1(P3_rEIP_PTR11), .A2(_03311__PTR9), .ZN(_03311__PTR10) );
  AND2_X1 U19270 ( .A1(P3_rEIP_PTR13), .A2(_03311__PTR11), .ZN(_03311__PTR12) );
  AND2_X1 U19271 ( .A1(P3_rEIP_PTR15), .A2(_03311__PTR13), .ZN(_03311__PTR14) );
  AND2_X1 U19272 ( .A1(P3_rEIP_PTR17), .A2(_03311__PTR15), .ZN(_03311__PTR16) );
  AND2_X1 U19273 ( .A1(P3_rEIP_PTR19), .A2(_03311__PTR17), .ZN(_03311__PTR18) );
  AND2_X1 U19274 ( .A1(P3_rEIP_PTR21), .A2(_03311__PTR19), .ZN(_03311__PTR20) );
  AND2_X1 U19275 ( .A1(P3_rEIP_PTR23), .A2(_03311__PTR21), .ZN(_03311__PTR22) );
  AND2_X1 U19276 ( .A1(P3_rEIP_PTR25), .A2(_03311__PTR23), .ZN(_03311__PTR24) );
  AND2_X1 U19277 ( .A1(P3_rEIP_PTR27), .A2(_03311__PTR25), .ZN(_03311__PTR26) );
  AND2_X1 U19278 ( .A1(P3_rEIP_PTR29), .A2(_03311__PTR27), .ZN(_03311__PTR28) );
  AND2_X1 U19279 ( .A1(_03224__PTR1), .A2(_02678__PTR32), .ZN(_03437__PTR1) );
  AND2_X1 U19280 ( .A1(_04850_), .A2(_03437__PTR1), .ZN(_03437__PTR3) );
  AND2_X1 U19281 ( .A1(_04879_), .A2(_03437__PTR3), .ZN(_03437__PTR7) );
  AND2_X1 U19282 ( .A1(_04886_), .A2(_03437__PTR7), .ZN(_03437__PTR15) );
  AND2_X1 U19283 ( .A1(_03224__PTR9), .A2(_03224__PTR8), .ZN(_04867_) );
  AND2_X1 U19284 ( .A1(_03224__PTR17), .A2(_03224__PTR16), .ZN(_04871_) );
  AND2_X1 U19285 ( .A1(_03224__PTR29), .A2(_03224__PTR28), .ZN(_04877_) );
  AND2_X1 U19286 ( .A1(_04887_), .A2(_03437__PTR15), .ZN(_03437__PTR23) );
  AND2_X1 U19287 ( .A1(_04880_), .A2(_03437__PTR7), .ZN(_03437__PTR11) );
  AND2_X1 U19288 ( .A1(_04882_), .A2(_03437__PTR15), .ZN(_03437__PTR19) );
  AND2_X1 U19289 ( .A1(_04884_), .A2(_03437__PTR23), .ZN(_03437__PTR27) );
  AND2_X1 U19290 ( .A1(_04865_), .A2(_03437__PTR3), .ZN(_03437__PTR5) );
  AND2_X1 U19291 ( .A1(_04867_), .A2(_03437__PTR7), .ZN(_03437__PTR9) );
  AND2_X1 U19292 ( .A1(_04869_), .A2(_03437__PTR11), .ZN(_03437__PTR13) );
  AND2_X1 U19293 ( .A1(_04871_), .A2(_03437__PTR15), .ZN(_03437__PTR17) );
  AND2_X1 U19294 ( .A1(_04873_), .A2(_03437__PTR19), .ZN(_03437__PTR21) );
  AND2_X1 U19295 ( .A1(_04875_), .A2(_03437__PTR23), .ZN(_03437__PTR25) );
  AND2_X1 U19296 ( .A1(_04877_), .A2(_03437__PTR27), .ZN(_03437__PTR29) );
  AND2_X1 U19297 ( .A1(_03224__PTR2), .A2(_03437__PTR1), .ZN(_03437__PTR2) );
  AND2_X1 U19298 ( .A1(_03224__PTR4), .A2(_03437__PTR3), .ZN(_03437__PTR4) );
  AND2_X1 U19299 ( .A1(_03224__PTR6), .A2(_03437__PTR5), .ZN(_03437__PTR6) );
  AND2_X1 U19300 ( .A1(_03224__PTR8), .A2(_03437__PTR7), .ZN(_03437__PTR8) );
  AND2_X1 U19301 ( .A1(_03224__PTR10), .A2(_03437__PTR9), .ZN(_03437__PTR10) );
  AND2_X1 U19302 ( .A1(_03224__PTR12), .A2(_03437__PTR11), .ZN(_03437__PTR12) );
  AND2_X1 U19303 ( .A1(_03224__PTR14), .A2(_03437__PTR13), .ZN(_03437__PTR14) );
  AND2_X1 U19304 ( .A1(_03224__PTR16), .A2(_03437__PTR15), .ZN(_03437__PTR16) );
  AND2_X1 U19305 ( .A1(_03224__PTR18), .A2(_03437__PTR17), .ZN(_03437__PTR18) );
  AND2_X1 U19306 ( .A1(_03224__PTR20), .A2(_03437__PTR19), .ZN(_03437__PTR20) );
  AND2_X1 U19307 ( .A1(_03224__PTR22), .A2(_03437__PTR21), .ZN(_03437__PTR22) );
  AND2_X1 U19308 ( .A1(_03224__PTR24), .A2(_03437__PTR23), .ZN(_03437__PTR24) );
  AND2_X1 U19309 ( .A1(_03224__PTR26), .A2(_03437__PTR25), .ZN(_03437__PTR26) );
  AND2_X1 U19310 ( .A1(_03224__PTR28), .A2(_03437__PTR27), .ZN(_03437__PTR28) );
  AND2_X1 U19311 ( .A1(_03224__PTR30), .A2(_03437__PTR29), .ZN(_03437__PTR30) );
  AND2_X1 U19312 ( .A1(_03224__PTR3), .A2(P3_EBX_PTR2), .ZN(_04835_) );
  AND2_X1 U19313 ( .A1(_03224__PTR5), .A2(P3_EBX_PTR4), .ZN(_04836_) );
  AND2_X1 U19314 ( .A1(_03224__PTR7), .A2(P3_EBX_PTR6), .ZN(_04837_) );
  AND2_X1 U19315 ( .A1(_03224__PTR9), .A2(P3_EBX_PTR8), .ZN(_04838_) );
  AND2_X1 U19316 ( .A1(_03224__PTR11), .A2(P3_EBX_PTR10), .ZN(_04839_) );
  AND2_X1 U19317 ( .A1(_03224__PTR13), .A2(P3_EBX_PTR12), .ZN(_04840_) );
  AND2_X1 U19318 ( .A1(_03224__PTR15), .A2(P3_EBX_PTR14), .ZN(_04841_) );
  AND2_X1 U19319 ( .A1(_03224__PTR17), .A2(P3_EBX_PTR16), .ZN(_04842_) );
  AND2_X1 U19320 ( .A1(_03224__PTR19), .A2(P3_EBX_PTR18), .ZN(_04843_) );
  AND2_X1 U19321 ( .A1(_03224__PTR21), .A2(P3_EBX_PTR20), .ZN(_04844_) );
  AND2_X1 U19322 ( .A1(_03224__PTR23), .A2(P3_EBX_PTR22), .ZN(_04845_) );
  AND2_X1 U19323 ( .A1(_03224__PTR25), .A2(P3_EBX_PTR24), .ZN(_04846_) );
  AND2_X1 U19324 ( .A1(_03224__PTR27), .A2(P3_EBX_PTR26), .ZN(_04847_) );
  AND2_X1 U19325 ( .A1(_03224__PTR29), .A2(P3_EBX_PTR28), .ZN(_04848_) );
  AND2_X1 U19326 ( .A1(_03222__PTR31), .A2(P3_EBX_PTR30), .ZN(_04849_) );
  AND2_X1 U19327 ( .A1(_04866_), .A2(_04891_), .ZN(_04851_) );
  AND2_X1 U19328 ( .A1(_04868_), .A2(_04893_), .ZN(_04852_) );
  AND2_X1 U19329 ( .A1(_04870_), .A2(_04895_), .ZN(_04853_) );
  AND2_X1 U19330 ( .A1(_04872_), .A2(_04897_), .ZN(_04854_) );
  AND2_X1 U19331 ( .A1(_04874_), .A2(_04899_), .ZN(_04855_) );
  AND2_X1 U19332 ( .A1(_04876_), .A2(_04901_), .ZN(_04856_) );
  AND2_X1 U19333 ( .A1(_04878_), .A2(_04903_), .ZN(_04857_) );
  AND2_X1 U19334 ( .A1(_04879_), .A2(_03223__PTR3), .ZN(_04858_) );
  AND2_X1 U19335 ( .A1(_04881_), .A2(_04905_), .ZN(_04859_) );
  AND2_X1 U19336 ( .A1(_04883_), .A2(_04907_), .ZN(_04860_) );
  AND2_X1 U19337 ( .A1(_04885_), .A2(_04909_), .ZN(_04861_) );
  AND2_X1 U19338 ( .A1(_04886_), .A2(_03223__PTR7), .ZN(_04862_) );
  AND2_X1 U19339 ( .A1(_04888_), .A2(_04912_), .ZN(_04863_) );
  AND2_X1 U19340 ( .A1(_04889_), .A2(_03223__PTR15), .ZN(_04864_) );
  AND2_X1 U19341 ( .A1(_03224__PTR3), .A2(_03224__PTR2), .ZN(_04850_) );
  AND2_X1 U19342 ( .A1(_03224__PTR5), .A2(_03224__PTR4), .ZN(_04865_) );
  AND2_X1 U19343 ( .A1(_03224__PTR7), .A2(_03224__PTR6), .ZN(_04866_) );
  AND2_X1 U19344 ( .A1(_03224__PTR11), .A2(_03224__PTR10), .ZN(_04868_) );
  AND2_X1 U19345 ( .A1(_03224__PTR13), .A2(_03224__PTR12), .ZN(_04869_) );
  AND2_X1 U19346 ( .A1(_03224__PTR15), .A2(_03224__PTR14), .ZN(_04870_) );
  AND2_X1 U19347 ( .A1(_03224__PTR19), .A2(_03224__PTR18), .ZN(_04872_) );
  AND2_X1 U19348 ( .A1(_03224__PTR21), .A2(_03224__PTR20), .ZN(_04873_) );
  AND2_X1 U19349 ( .A1(_03224__PTR23), .A2(_03224__PTR22), .ZN(_04874_) );
  AND2_X1 U19350 ( .A1(_03224__PTR25), .A2(_03224__PTR24), .ZN(_04875_) );
  AND2_X1 U19351 ( .A1(_03224__PTR27), .A2(_03224__PTR26), .ZN(_04876_) );
  AND2_X1 U19352 ( .A1(_03222__PTR31), .A2(_03224__PTR30), .ZN(_04878_) );
  AND2_X1 U19353 ( .A1(_04866_), .A2(_04865_), .ZN(_04879_) );
  AND2_X1 U19354 ( .A1(_04868_), .A2(_04867_), .ZN(_04880_) );
  AND2_X1 U19355 ( .A1(_04870_), .A2(_04869_), .ZN(_04881_) );
  AND2_X1 U19356 ( .A1(_04872_), .A2(_04871_), .ZN(_04882_) );
  AND2_X1 U19357 ( .A1(_04874_), .A2(_04873_), .ZN(_04883_) );
  AND2_X1 U19358 ( .A1(_04876_), .A2(_04875_), .ZN(_04884_) );
  AND2_X1 U19359 ( .A1(_04878_), .A2(_04877_), .ZN(_04885_) );
  AND2_X1 U19360 ( .A1(_04881_), .A2(_04880_), .ZN(_04886_) );
  AND2_X1 U19361 ( .A1(_04883_), .A2(_04882_), .ZN(_04887_) );
  AND2_X1 U19362 ( .A1(_04885_), .A2(_04884_), .ZN(_04888_) );
  AND2_X1 U19363 ( .A1(_04888_), .A2(_04887_), .ZN(_04889_) );
  OR2_X1 U19364 ( .A1(P3_EBX_PTR3), .A2(_04835_), .ZN(_04890_) );
  OR2_X1 U19365 ( .A1(P3_EBX_PTR5), .A2(_04836_), .ZN(_04891_) );
  OR2_X1 U19366 ( .A1(P3_EBX_PTR7), .A2(_04837_), .ZN(_04892_) );
  OR2_X1 U19367 ( .A1(P3_EBX_PTR9), .A2(_04838_), .ZN(_04893_) );
  OR2_X1 U19368 ( .A1(P3_EBX_PTR11), .A2(_04839_), .ZN(_04894_) );
  OR2_X1 U19369 ( .A1(P3_EBX_PTR13), .A2(_04840_), .ZN(_04895_) );
  OR2_X1 U19370 ( .A1(P3_EBX_PTR15), .A2(_04841_), .ZN(_04896_) );
  OR2_X1 U19371 ( .A1(P3_EBX_PTR17), .A2(_04842_), .ZN(_04897_) );
  OR2_X1 U19372 ( .A1(P3_EBX_PTR19), .A2(_04843_), .ZN(_04898_) );
  OR2_X1 U19373 ( .A1(P3_EBX_PTR21), .A2(_04844_), .ZN(_04899_) );
  OR2_X1 U19374 ( .A1(P3_EBX_PTR23), .A2(_04845_), .ZN(_04900_) );
  OR2_X1 U19375 ( .A1(P3_EBX_PTR25), .A2(_04846_), .ZN(_04901_) );
  OR2_X1 U19376 ( .A1(P3_EBX_PTR27), .A2(_04847_), .ZN(_04902_) );
  OR2_X1 U19377 ( .A1(P3_EBX_PTR29), .A2(_04848_), .ZN(_04903_) );
  OR2_X1 U19378 ( .A1(_04890_), .A2(_04850_), .ZN(_03223__PTR3) );
  OR2_X1 U19379 ( .A1(_04892_), .A2(_04851_), .ZN(_04904_) );
  OR2_X1 U19380 ( .A1(_04894_), .A2(_04852_), .ZN(_04905_) );
  OR2_X1 U19381 ( .A1(_04896_), .A2(_04853_), .ZN(_04906_) );
  OR2_X1 U19382 ( .A1(_04898_), .A2(_04854_), .ZN(_04907_) );
  OR2_X1 U19383 ( .A1(_04900_), .A2(_04855_), .ZN(_04908_) );
  OR2_X1 U19384 ( .A1(_04902_), .A2(_04856_), .ZN(_04909_) );
  OR2_X1 U19385 ( .A1(_04849_), .A2(_04857_), .ZN(_04910_) );
  OR2_X1 U19386 ( .A1(_04904_), .A2(_04858_), .ZN(_03223__PTR7) );
  OR2_X1 U19387 ( .A1(_04906_), .A2(_04859_), .ZN(_04911_) );
  OR2_X1 U19388 ( .A1(_04908_), .A2(_04860_), .ZN(_04912_) );
  OR2_X1 U19389 ( .A1(_04910_), .A2(_04861_), .ZN(_04913_) );
  OR2_X1 U19390 ( .A1(_04911_), .A2(_04862_), .ZN(_03223__PTR15) );
  OR2_X1 U19391 ( .A1(_04913_), .A2(_04863_), .ZN(_04914_) );
  OR2_X1 U19392 ( .A1(_04914_), .A2(_04864_), .ZN(_03223__PTR31) );
  AND2_X1 U19393 ( .A1(_03422__PTR1), .A2(_03421__PTR0), .ZN(_05273_) );
  AND2_X1 U19394 ( .A1(_03422__PTR3), .A2(_03423__PTR2), .ZN(_05274_) );
  AND2_X1 U19395 ( .A1(_05276_), .A2(_03421__PTR1), .ZN(_05275_) );
  AND2_X1 U19396 ( .A1(_03422__PTR3), .A2(_03422__PTR2), .ZN(_05276_) );
  AND2_X1 U19397 ( .A1(_03422__PTR2), .A2(_03421__PTR1), .ZN(_05278_) );
  AND2_X1 U19398 ( .A1(_03422__PTR4), .A2(_03421__PTR3), .ZN(_05277_) );
  OR2_X1 U19399 ( .A1(_03423__PTR0), .A2(_03208__PTR0), .ZN(_03421__PTR0) );
  OR2_X1 U19400 ( .A1(_03423__PTR1), .A2(_05273_), .ZN(_03421__PTR1) );
  OR2_X1 U19401 ( .A1(_03423__PTR3), .A2(_05274_), .ZN(_05279_) );
  OR2_X1 U19402 ( .A1(_05279_), .A2(_05275_), .ZN(_03421__PTR3) );
  OR2_X1 U19403 ( .A1(_03423__PTR4), .A2(_05277_), .ZN(_03210__PTR5) );
  OR2_X1 U19404 ( .A1(_03423__PTR2), .A2(_05278_), .ZN(_03421__PTR2) );
  AND2_X1 U19405 ( .A1(_03207__PTR1), .A2(_03208__PTR0), .ZN(_01266__PTR0) );
  AND2_X1 U19406 ( .A1(_03209__PTR3), .A2(_03219__PTR1), .ZN(_03219__PTR3) );
  AND2_X1 U19407 ( .A1(_01266__PTR2), .A2(_03219__PTR3), .ZN(_04834_) );
  OR2_X1 U19408 ( .A1(_03208__PTR1), .A2(_01266__PTR0), .ZN(_03219__PTR1) );
  OR2_X1 U19409 ( .A1(_03206__PTR5), .A2(_04834_), .ZN(_03219__PTR5) );
  AND2_X1 U19410 ( .A1(P3_P1_InstQueueRd_Addr_PTR1), .A2(P3_P1_InstQueueRd_Addr_PTR0), .ZN(_03240__PTR1) );
  AND2_X1 U19411 ( .A1(_02467__PTR5), .A2(_03240__PTR1), .ZN(_05228_) );
  OR2_X1 U19412 ( .A1(P3_P1_InstQueueRd_Addr_PTR2), .A2(_05228_), .ZN(_03309__PTR2) );
  AND2_X1 U19413 ( .A1(P3_P1_InstQueueRd_Addr_PTR2), .A2(P3_P1_InstQueueRd_Addr_PTR1), .ZN(_03307__PTR1) );
  AND2_X1 U19414 ( .A1(P3_P1_InstQueueRd_Addr_PTR3), .A2(_03307__PTR1), .ZN(_03307__PTR2) );
  AND2_X1 U19415 ( .A1(_02468__PTR1), .A2(_03304__PTR0), .ZN(_03304__PTR1) );
  AND2_X1 U19416 ( .A1(_05224_), .A2(_03304__PTR1), .ZN(_03304__PTR3) );
  AND2_X1 U19417 ( .A1(_05227_), .A2(_03304__PTR3), .ZN(_03304__PTR7) );
  AND2_X1 U19418 ( .A1(_02468__PTR3), .A2(_02468__PTR2), .ZN(_05224_) );
  AND2_X1 U19419 ( .A1(_02468__PTR5), .A2(_02468__PTR4), .ZN(_05225_) );
  AND2_X1 U19420 ( .A1(_02468__PTR7), .A2(_02468__PTR6), .ZN(_05226_) );
  AND2_X1 U19421 ( .A1(_05226_), .A2(_05225_), .ZN(_05227_) );
  AND2_X1 U19422 ( .A1(_05225_), .A2(_03304__PTR3), .ZN(_03304__PTR5) );
  AND2_X1 U19423 ( .A1(_02468__PTR2), .A2(_03304__PTR1), .ZN(_03304__PTR2) );
  AND2_X1 U19424 ( .A1(_02468__PTR4), .A2(_03304__PTR3), .ZN(_03304__PTR4) );
  AND2_X1 U19425 ( .A1(_02468__PTR6), .A2(_03304__PTR5), .ZN(_03304__PTR6) );
  AND2_X1 U19426 ( .A1(_02471__PTR4), .A2(P3_P1_InstQueueRd_Addr_PTR0), .ZN(_05223_) );
  AND2_X1 U19427 ( .A1(P3_P1_InstQueueRd_Addr_PTR3), .A2(P3_P1_InstQueueRd_Addr_PTR2), .ZN(_03302__PTR1) );
  AND2_X1 U19428 ( .A1(P3_P1_InstQueueRd_Addr_PTR2), .A2(_03303__PTR1), .ZN(_03303__PTR2) );
  OR2_X1 U19429 ( .A1(P3_P1_InstQueueRd_Addr_PTR1), .A2(_05223_), .ZN(_03303__PTR1) );
  AND2_X1 U19430 ( .A1(_05184_), .A2(_03288__PTR1), .ZN(_05183_) );
  AND2_X1 U19431 ( .A1(_05116_), .A2(_03296__PTR3), .ZN(_03296__PTR7) );
  AND2_X1 U19432 ( .A1(_05122_), .A2(_03296__PTR7), .ZN(_03296__PTR15) );
  AND2_X1 U19433 ( .A1(P3_P1_InstAddrPointer_PTR3), .A2(_03235__PTR2), .ZN(_05184_) );
  AND2_X1 U19434 ( .A1(P3_P1_InstAddrPointer_PTR11), .A2(P3_P1_InstAddrPointer_PTR10), .ZN(_05106_) );
  AND2_X1 U19435 ( .A1(P3_P1_InstAddrPointer_PTR25), .A2(P3_P1_InstAddrPointer_PTR24), .ZN(_05113_) );
  AND2_X1 U19436 ( .A1(_05106_), .A2(_05105_), .ZN(_05117_) );
  AND2_X1 U19437 ( .A1(_05110_), .A2(_05109_), .ZN(_05119_) );
  AND2_X1 U19438 ( .A1(_05123_), .A2(_03296__PTR15), .ZN(_03296__PTR23) );
  AND2_X1 U19439 ( .A1(_05117_), .A2(_03296__PTR7), .ZN(_03296__PTR11) );
  AND2_X1 U19440 ( .A1(_05119_), .A2(_03296__PTR15), .ZN(_03296__PTR19) );
  AND2_X1 U19441 ( .A1(_05121_), .A2(_03296__PTR23), .ZN(_03296__PTR27) );
  AND2_X1 U19442 ( .A1(_05103_), .A2(_03296__PTR3), .ZN(_03296__PTR5) );
  AND2_X1 U19443 ( .A1(_05105_), .A2(_03296__PTR7), .ZN(_03296__PTR9) );
  AND2_X1 U19444 ( .A1(_05107_), .A2(_03296__PTR11), .ZN(_03296__PTR13) );
  AND2_X1 U19445 ( .A1(_05109_), .A2(_03296__PTR15), .ZN(_03296__PTR17) );
  AND2_X1 U19446 ( .A1(_05111_), .A2(_03296__PTR19), .ZN(_03296__PTR21) );
  AND2_X1 U19447 ( .A1(_05113_), .A2(_03296__PTR23), .ZN(_03296__PTR25) );
  AND2_X1 U19448 ( .A1(_05115_), .A2(_03296__PTR27), .ZN(_03296__PTR29) );
  AND2_X1 U19449 ( .A1(_03235__PTR2), .A2(_03288__PTR1), .ZN(_05185_) );
  AND2_X1 U19450 ( .A1(P3_P1_InstAddrPointer_PTR4), .A2(_03296__PTR3), .ZN(_03296__PTR4) );
  AND2_X1 U19451 ( .A1(P3_P1_InstAddrPointer_PTR6), .A2(_03296__PTR5), .ZN(_03296__PTR6) );
  AND2_X1 U19452 ( .A1(P3_P1_InstAddrPointer_PTR8), .A2(_03296__PTR7), .ZN(_03296__PTR8) );
  AND2_X1 U19453 ( .A1(P3_P1_InstAddrPointer_PTR10), .A2(_03296__PTR9), .ZN(_03296__PTR10) );
  AND2_X1 U19454 ( .A1(P3_P1_InstAddrPointer_PTR12), .A2(_03296__PTR11), .ZN(_03296__PTR12) );
  AND2_X1 U19455 ( .A1(P3_P1_InstAddrPointer_PTR14), .A2(_03296__PTR13), .ZN(_03296__PTR14) );
  AND2_X1 U19456 ( .A1(P3_P1_InstAddrPointer_PTR16), .A2(_03296__PTR15), .ZN(_03296__PTR16) );
  AND2_X1 U19457 ( .A1(P3_P1_InstAddrPointer_PTR18), .A2(_03296__PTR17), .ZN(_03296__PTR18) );
  AND2_X1 U19458 ( .A1(P3_P1_InstAddrPointer_PTR20), .A2(_03296__PTR19), .ZN(_03296__PTR20) );
  AND2_X1 U19459 ( .A1(P3_P1_InstAddrPointer_PTR22), .A2(_03296__PTR21), .ZN(_03296__PTR22) );
  AND2_X1 U19460 ( .A1(P3_P1_InstAddrPointer_PTR24), .A2(_03296__PTR23), .ZN(_03296__PTR24) );
  AND2_X1 U19461 ( .A1(P3_P1_InstAddrPointer_PTR26), .A2(_03296__PTR25), .ZN(_03296__PTR26) );
  AND2_X1 U19462 ( .A1(P3_P1_InstAddrPointer_PTR28), .A2(_03296__PTR27), .ZN(_03296__PTR28) );
  AND2_X1 U19463 ( .A1(P3_P1_InstAddrPointer_PTR30), .A2(_03296__PTR29), .ZN(_03296__PTR30) );
  OR2_X1 U19464 ( .A1(_05102_), .A2(_05183_), .ZN(_03296__PTR3) );
  OR2_X1 U19465 ( .A1(P3_P1_InstAddrPointer_PTR2), .A2(_05185_), .ZN(_03296__PTR2) );
  AND2_X1 U19466 ( .A1(_03299__PTR1), .A2(_03298__PTR0), .ZN(_05186_) );
  AND2_X1 U19467 ( .A1(_03299__PTR3), .A2(_03301__PTR2), .ZN(_05187_) );
  AND2_X1 U19468 ( .A1(_03299__PTR5), .A2(_03301__PTR4), .ZN(_05188_) );
  AND2_X1 U19469 ( .A1(_03299__PTR7), .A2(_03301__PTR6), .ZN(_05189_) );
  AND2_X1 U19470 ( .A1(_05193_), .A2(_03298__PTR1), .ZN(_05190_) );
  AND2_X1 U19471 ( .A1(_05195_), .A2(_05220_), .ZN(_05191_) );
  AND2_X1 U19472 ( .A1(_05207_), .A2(_03298__PTR3), .ZN(_05192_) );
  AND2_X1 U19473 ( .A1(_05213_), .A2(_03298__PTR7), .ZN(_03298__PTR15) );
  AND2_X1 U19474 ( .A1(_03299__PTR3), .A2(_03299__PTR2), .ZN(_05193_) );
  AND2_X1 U19475 ( .A1(_03299__PTR5), .A2(_03299__PTR4), .ZN(_05194_) );
  AND2_X1 U19476 ( .A1(_03299__PTR7), .A2(_03299__PTR6), .ZN(_05195_) );
  AND2_X1 U19477 ( .A1(_03297__PTR9), .A2(_03297__PTR8), .ZN(_05196_) );
  AND2_X1 U19478 ( .A1(_03297__PTR11), .A2(_03297__PTR10), .ZN(_05197_) );
  AND2_X1 U19479 ( .A1(_03297__PTR13), .A2(_03297__PTR12), .ZN(_05198_) );
  AND2_X1 U19480 ( .A1(_03297__PTR15), .A2(_03297__PTR14), .ZN(_05199_) );
  AND2_X1 U19481 ( .A1(_03297__PTR17), .A2(_03297__PTR16), .ZN(_05200_) );
  AND2_X1 U19482 ( .A1(_03297__PTR19), .A2(_03297__PTR18), .ZN(_05201_) );
  AND2_X1 U19483 ( .A1(_03297__PTR21), .A2(_03297__PTR20), .ZN(_05202_) );
  AND2_X1 U19484 ( .A1(_03297__PTR23), .A2(_03297__PTR22), .ZN(_05203_) );
  AND2_X1 U19485 ( .A1(_03297__PTR25), .A2(_03297__PTR24), .ZN(_05204_) );
  AND2_X1 U19486 ( .A1(_03297__PTR27), .A2(_03297__PTR26), .ZN(_05205_) );
  AND2_X1 U19487 ( .A1(_03297__PTR29), .A2(_03297__PTR28), .ZN(_05206_) );
  AND2_X1 U19488 ( .A1(_05195_), .A2(_05194_), .ZN(_05207_) );
  AND2_X1 U19489 ( .A1(_05197_), .A2(_05196_), .ZN(_05208_) );
  AND2_X1 U19490 ( .A1(_05199_), .A2(_05198_), .ZN(_05209_) );
  AND2_X1 U19491 ( .A1(_05201_), .A2(_05200_), .ZN(_05210_) );
  AND2_X1 U19492 ( .A1(_05203_), .A2(_05202_), .ZN(_05211_) );
  AND2_X1 U19493 ( .A1(_05205_), .A2(_05204_), .ZN(_05212_) );
  AND2_X1 U19494 ( .A1(_05209_), .A2(_05208_), .ZN(_05213_) );
  AND2_X1 U19495 ( .A1(_05211_), .A2(_05210_), .ZN(_05214_) );
  AND2_X1 U19496 ( .A1(_05214_), .A2(_03298__PTR15), .ZN(_03298__PTR23) );
  AND2_X1 U19497 ( .A1(_05208_), .A2(_03298__PTR7), .ZN(_03298__PTR11) );
  AND2_X1 U19498 ( .A1(_05210_), .A2(_03298__PTR15), .ZN(_03298__PTR19) );
  AND2_X1 U19499 ( .A1(_05212_), .A2(_03298__PTR23), .ZN(_03298__PTR27) );
  AND2_X1 U19500 ( .A1(_05194_), .A2(_03298__PTR3), .ZN(_05215_) );
  AND2_X1 U19501 ( .A1(_05196_), .A2(_03298__PTR7), .ZN(_03298__PTR9) );
  AND2_X1 U19502 ( .A1(_05198_), .A2(_03298__PTR11), .ZN(_03298__PTR13) );
  AND2_X1 U19503 ( .A1(_05200_), .A2(_03298__PTR15), .ZN(_03298__PTR17) );
  AND2_X1 U19504 ( .A1(_05202_), .A2(_03298__PTR19), .ZN(_03298__PTR21) );
  AND2_X1 U19505 ( .A1(_05204_), .A2(_03298__PTR23), .ZN(_03298__PTR25) );
  AND2_X1 U19506 ( .A1(_05206_), .A2(_03298__PTR27), .ZN(_03298__PTR29) );
  AND2_X1 U19507 ( .A1(_03299__PTR2), .A2(_03298__PTR1), .ZN(_05216_) );
  AND2_X1 U19508 ( .A1(_03299__PTR4), .A2(_03298__PTR3), .ZN(_05217_) );
  AND2_X1 U19509 ( .A1(_03299__PTR6), .A2(_03298__PTR5), .ZN(_05218_) );
  AND2_X1 U19510 ( .A1(_03297__PTR8), .A2(_03298__PTR7), .ZN(_03298__PTR8) );
  AND2_X1 U19511 ( .A1(_03297__PTR10), .A2(_03298__PTR9), .ZN(_03298__PTR10) );
  AND2_X1 U19512 ( .A1(_03297__PTR12), .A2(_03298__PTR11), .ZN(_03298__PTR12) );
  AND2_X1 U19513 ( .A1(_03297__PTR14), .A2(_03298__PTR13), .ZN(_03298__PTR14) );
  AND2_X1 U19514 ( .A1(_03297__PTR16), .A2(_03298__PTR15), .ZN(_03298__PTR16) );
  AND2_X1 U19515 ( .A1(_03297__PTR18), .A2(_03298__PTR17), .ZN(_03298__PTR18) );
  AND2_X1 U19516 ( .A1(_03297__PTR20), .A2(_03298__PTR19), .ZN(_03298__PTR20) );
  AND2_X1 U19517 ( .A1(_03297__PTR22), .A2(_03298__PTR21), .ZN(_03298__PTR22) );
  AND2_X1 U19518 ( .A1(_03297__PTR24), .A2(_03298__PTR23), .ZN(_03298__PTR24) );
  AND2_X1 U19519 ( .A1(_03297__PTR26), .A2(_03298__PTR25), .ZN(_03298__PTR26) );
  AND2_X1 U19520 ( .A1(_03297__PTR28), .A2(_03298__PTR27), .ZN(_03298__PTR28) );
  AND2_X1 U19521 ( .A1(_03297__PTR30), .A2(_03298__PTR29), .ZN(_03298__PTR30) );
  OR2_X1 U19522 ( .A1(_03301__PTR1), .A2(_05186_), .ZN(_03298__PTR1) );
  OR2_X1 U19523 ( .A1(_03301__PTR3), .A2(_05187_), .ZN(_05219_) );
  OR2_X1 U19524 ( .A1(_03301__PTR5), .A2(_05188_), .ZN(_05220_) );
  OR2_X1 U19525 ( .A1(_03301__PTR7), .A2(_05189_), .ZN(_05221_) );
  OR2_X1 U19526 ( .A1(_05219_), .A2(_05190_), .ZN(_03298__PTR3) );
  OR2_X1 U19527 ( .A1(_05221_), .A2(_05191_), .ZN(_05222_) );
  OR2_X1 U19528 ( .A1(_05222_), .A2(_05192_), .ZN(_03298__PTR7) );
  OR2_X1 U19529 ( .A1(_05220_), .A2(_05215_), .ZN(_03298__PTR5) );
  OR2_X1 U19530 ( .A1(_03301__PTR2), .A2(_05216_), .ZN(_03298__PTR2) );
  OR2_X1 U19531 ( .A1(_03301__PTR4), .A2(_05217_), .ZN(_03298__PTR4) );
  OR2_X1 U19532 ( .A1(_03301__PTR6), .A2(_05218_), .ZN(_03298__PTR6) );
  AND2_X1 U19533 ( .A1(_03208__PTR3), .A2(_03208__PTR2), .ZN(_03209__PTR3) );
  AND2_X1 U19534 ( .A1(_01268__PTR1), .A2(_03208__PTR1), .ZN(_04832_) );
  AND2_X1 U19535 ( .A1(_03208__PTR3), .A2(_03207__PTR2), .ZN(_01268__PTR1) );
  AND2_X1 U19536 ( .A1(_03210__PTR5), .A2(_03208__PTR4), .ZN(_01266__PTR2) );
  AND2_X1 U19537 ( .A1(_01266__PTR2), .A2(_03216__PTR3), .ZN(_04833_) );
  OR2_X1 U19538 ( .A1(_03209__PTR3), .A2(_04832_), .ZN(_03216__PTR3) );
  OR2_X1 U19539 ( .A1(_03206__PTR5), .A2(_04833_), .ZN(_03216__PTR5) );
  AND2_X1 U19540 ( .A1(P3_P1_InstAddrPointer_PTR2), .A2(P3_P1_InstAddrPointer_PTR1), .ZN(_03291__PTR1) );
  AND2_X1 U19541 ( .A1(_05124_), .A2(_03291__PTR1), .ZN(_03291__PTR3) );
  AND2_X1 U19542 ( .A1(_05138_), .A2(_03291__PTR3), .ZN(_03291__PTR7) );
  AND2_X1 U19543 ( .A1(_05144_), .A2(_03291__PTR7), .ZN(_03291__PTR15) );
  AND2_X1 U19544 ( .A1(P3_P1_InstAddrPointer_PTR4), .A2(P3_P1_InstAddrPointer_PTR3), .ZN(_05124_) );
  AND2_X1 U19545 ( .A1(P3_P1_InstAddrPointer_PTR6), .A2(P3_P1_InstAddrPointer_PTR5), .ZN(_05125_) );
  AND2_X1 U19546 ( .A1(P3_P1_InstAddrPointer_PTR8), .A2(P3_P1_InstAddrPointer_PTR7), .ZN(_05126_) );
  AND2_X1 U19547 ( .A1(P3_P1_InstAddrPointer_PTR10), .A2(P3_P1_InstAddrPointer_PTR9), .ZN(_05127_) );
  AND2_X1 U19548 ( .A1(P3_P1_InstAddrPointer_PTR12), .A2(P3_P1_InstAddrPointer_PTR11), .ZN(_05128_) );
  AND2_X1 U19549 ( .A1(P3_P1_InstAddrPointer_PTR14), .A2(P3_P1_InstAddrPointer_PTR13), .ZN(_05129_) );
  AND2_X1 U19550 ( .A1(P3_P1_InstAddrPointer_PTR16), .A2(P3_P1_InstAddrPointer_PTR15), .ZN(_05130_) );
  AND2_X1 U19551 ( .A1(P3_P1_InstAddrPointer_PTR18), .A2(P3_P1_InstAddrPointer_PTR17), .ZN(_05131_) );
  AND2_X1 U19552 ( .A1(P3_P1_InstAddrPointer_PTR20), .A2(P3_P1_InstAddrPointer_PTR19), .ZN(_05132_) );
  AND2_X1 U19553 ( .A1(P3_P1_InstAddrPointer_PTR22), .A2(P3_P1_InstAddrPointer_PTR21), .ZN(_05133_) );
  AND2_X1 U19554 ( .A1(P3_P1_InstAddrPointer_PTR24), .A2(P3_P1_InstAddrPointer_PTR23), .ZN(_05134_) );
  AND2_X1 U19555 ( .A1(P3_P1_InstAddrPointer_PTR26), .A2(P3_P1_InstAddrPointer_PTR25), .ZN(_05135_) );
  AND2_X1 U19556 ( .A1(P3_P1_InstAddrPointer_PTR28), .A2(P3_P1_InstAddrPointer_PTR27), .ZN(_05136_) );
  AND2_X1 U19557 ( .A1(P3_P1_InstAddrPointer_PTR30), .A2(P3_P1_InstAddrPointer_PTR29), .ZN(_05137_) );
  AND2_X1 U19558 ( .A1(_05126_), .A2(_05125_), .ZN(_05138_) );
  AND2_X1 U19559 ( .A1(_05128_), .A2(_05127_), .ZN(_05139_) );
  AND2_X1 U19560 ( .A1(_05130_), .A2(_05129_), .ZN(_05140_) );
  AND2_X1 U19561 ( .A1(_05132_), .A2(_05131_), .ZN(_05141_) );
  AND2_X1 U19562 ( .A1(_05134_), .A2(_05133_), .ZN(_05142_) );
  AND2_X1 U19563 ( .A1(_05136_), .A2(_05135_), .ZN(_05143_) );
  AND2_X1 U19564 ( .A1(_05140_), .A2(_05139_), .ZN(_05144_) );
  AND2_X1 U19565 ( .A1(_05142_), .A2(_05141_), .ZN(_05145_) );
  AND2_X1 U19566 ( .A1(_05145_), .A2(_03291__PTR15), .ZN(_03291__PTR23) );
  AND2_X1 U19567 ( .A1(_05139_), .A2(_03291__PTR7), .ZN(_03291__PTR11) );
  AND2_X1 U19568 ( .A1(_05141_), .A2(_03291__PTR15), .ZN(_03291__PTR19) );
  AND2_X1 U19569 ( .A1(_05143_), .A2(_03291__PTR23), .ZN(_03291__PTR27) );
  AND2_X1 U19570 ( .A1(_05125_), .A2(_03291__PTR3), .ZN(_03291__PTR5) );
  AND2_X1 U19571 ( .A1(_05127_), .A2(_03291__PTR7), .ZN(_03291__PTR9) );
  AND2_X1 U19572 ( .A1(_05129_), .A2(_03291__PTR11), .ZN(_03291__PTR13) );
  AND2_X1 U19573 ( .A1(_05131_), .A2(_03291__PTR15), .ZN(_03291__PTR17) );
  AND2_X1 U19574 ( .A1(_05133_), .A2(_03291__PTR19), .ZN(_03291__PTR21) );
  AND2_X1 U19575 ( .A1(_05135_), .A2(_03291__PTR23), .ZN(_03291__PTR25) );
  AND2_X1 U19576 ( .A1(_05137_), .A2(_03291__PTR27), .ZN(_03291__PTR29) );
  AND2_X1 U19577 ( .A1(P3_P1_InstAddrPointer_PTR3), .A2(_03291__PTR1), .ZN(_03291__PTR2) );
  AND2_X1 U19578 ( .A1(P3_P1_InstAddrPointer_PTR5), .A2(_03291__PTR3), .ZN(_03291__PTR4) );
  AND2_X1 U19579 ( .A1(P3_P1_InstAddrPointer_PTR7), .A2(_03291__PTR5), .ZN(_03291__PTR6) );
  AND2_X1 U19580 ( .A1(P3_P1_InstAddrPointer_PTR9), .A2(_03291__PTR7), .ZN(_03291__PTR8) );
  AND2_X1 U19581 ( .A1(P3_P1_InstAddrPointer_PTR11), .A2(_03291__PTR9), .ZN(_03291__PTR10) );
  AND2_X1 U19582 ( .A1(P3_P1_InstAddrPointer_PTR13), .A2(_03291__PTR11), .ZN(_03291__PTR12) );
  AND2_X1 U19583 ( .A1(P3_P1_InstAddrPointer_PTR15), .A2(_03291__PTR13), .ZN(_03291__PTR14) );
  AND2_X1 U19584 ( .A1(P3_P1_InstAddrPointer_PTR17), .A2(_03291__PTR15), .ZN(_03291__PTR16) );
  AND2_X1 U19585 ( .A1(P3_P1_InstAddrPointer_PTR19), .A2(_03291__PTR17), .ZN(_03291__PTR18) );
  AND2_X1 U19586 ( .A1(P3_P1_InstAddrPointer_PTR21), .A2(_03291__PTR19), .ZN(_03291__PTR20) );
  AND2_X1 U19587 ( .A1(P3_P1_InstAddrPointer_PTR23), .A2(_03291__PTR21), .ZN(_03291__PTR22) );
  AND2_X1 U19588 ( .A1(P3_P1_InstAddrPointer_PTR25), .A2(_03291__PTR23), .ZN(_03291__PTR24) );
  AND2_X1 U19589 ( .A1(P3_P1_InstAddrPointer_PTR27), .A2(_03291__PTR25), .ZN(_03291__PTR26) );
  AND2_X1 U19590 ( .A1(P3_P1_InstAddrPointer_PTR29), .A2(_03291__PTR27), .ZN(_03291__PTR28) );
  AND2_X1 U19591 ( .A1(_03293__PTR1), .A2(_03292__PTR0), .ZN(_05146_) );
  AND2_X1 U19592 ( .A1(_03293__PTR3), .A2(_03295__PTR2), .ZN(_05147_) );
  AND2_X1 U19593 ( .A1(_03293__PTR5), .A2(_03295__PTR4), .ZN(_05148_) );
  AND2_X1 U19594 ( .A1(_03293__PTR7), .A2(_03295__PTR6), .ZN(_05149_) );
  AND2_X1 U19595 ( .A1(_05153_), .A2(_03292__PTR1), .ZN(_05150_) );
  AND2_X1 U19596 ( .A1(_05155_), .A2(_05180_), .ZN(_05151_) );
  AND2_X1 U19597 ( .A1(_05167_), .A2(_03292__PTR3), .ZN(_05152_) );
  AND2_X1 U19598 ( .A1(_05173_), .A2(_03292__PTR7), .ZN(_03292__PTR15) );
  AND2_X1 U19599 ( .A1(_03293__PTR3), .A2(_03293__PTR2), .ZN(_05153_) );
  AND2_X1 U19600 ( .A1(_03293__PTR5), .A2(_03293__PTR4), .ZN(_05154_) );
  AND2_X1 U19601 ( .A1(_03293__PTR7), .A2(_03293__PTR6), .ZN(_05155_) );
  AND2_X1 U19602 ( .A1(_02662__PTR41), .A2(_02662__PTR40), .ZN(_05156_) );
  AND2_X1 U19603 ( .A1(_02662__PTR43), .A2(_02662__PTR42), .ZN(_05157_) );
  AND2_X1 U19604 ( .A1(_02662__PTR45), .A2(_02662__PTR44), .ZN(_05158_) );
  AND2_X1 U19605 ( .A1(_02662__PTR47), .A2(_02662__PTR46), .ZN(_05159_) );
  AND2_X1 U19606 ( .A1(_02662__PTR49), .A2(_02662__PTR48), .ZN(_05160_) );
  AND2_X1 U19607 ( .A1(_02662__PTR51), .A2(_02662__PTR50), .ZN(_05161_) );
  AND2_X1 U19608 ( .A1(_02662__PTR53), .A2(_02662__PTR52), .ZN(_05162_) );
  AND2_X1 U19609 ( .A1(_02662__PTR55), .A2(_02662__PTR54), .ZN(_05163_) );
  AND2_X1 U19610 ( .A1(_02662__PTR57), .A2(_02662__PTR56), .ZN(_05164_) );
  AND2_X1 U19611 ( .A1(_02662__PTR59), .A2(_02662__PTR58), .ZN(_05165_) );
  AND2_X1 U19612 ( .A1(_02662__PTR61), .A2(_02662__PTR60), .ZN(_05166_) );
  AND2_X1 U19613 ( .A1(_05155_), .A2(_05154_), .ZN(_05167_) );
  AND2_X1 U19614 ( .A1(_05157_), .A2(_05156_), .ZN(_05168_) );
  AND2_X1 U19615 ( .A1(_05159_), .A2(_05158_), .ZN(_05169_) );
  AND2_X1 U19616 ( .A1(_05161_), .A2(_05160_), .ZN(_05170_) );
  AND2_X1 U19617 ( .A1(_05163_), .A2(_05162_), .ZN(_05171_) );
  AND2_X1 U19618 ( .A1(_05165_), .A2(_05164_), .ZN(_05172_) );
  AND2_X1 U19619 ( .A1(_05169_), .A2(_05168_), .ZN(_05173_) );
  AND2_X1 U19620 ( .A1(_05171_), .A2(_05170_), .ZN(_05174_) );
  AND2_X1 U19621 ( .A1(_05174_), .A2(_03292__PTR15), .ZN(_03292__PTR23) );
  AND2_X1 U19622 ( .A1(_05168_), .A2(_03292__PTR7), .ZN(_03292__PTR11) );
  AND2_X1 U19623 ( .A1(_05170_), .A2(_03292__PTR15), .ZN(_03292__PTR19) );
  AND2_X1 U19624 ( .A1(_05172_), .A2(_03292__PTR23), .ZN(_03292__PTR27) );
  AND2_X1 U19625 ( .A1(_05154_), .A2(_03292__PTR3), .ZN(_05175_) );
  AND2_X1 U19626 ( .A1(_05156_), .A2(_03292__PTR7), .ZN(_03292__PTR9) );
  AND2_X1 U19627 ( .A1(_05158_), .A2(_03292__PTR11), .ZN(_03292__PTR13) );
  AND2_X1 U19628 ( .A1(_05160_), .A2(_03292__PTR15), .ZN(_03292__PTR17) );
  AND2_X1 U19629 ( .A1(_05162_), .A2(_03292__PTR19), .ZN(_03292__PTR21) );
  AND2_X1 U19630 ( .A1(_05164_), .A2(_03292__PTR23), .ZN(_03292__PTR25) );
  AND2_X1 U19631 ( .A1(_05166_), .A2(_03292__PTR27), .ZN(_03292__PTR29) );
  AND2_X1 U19632 ( .A1(_03293__PTR2), .A2(_03292__PTR1), .ZN(_05176_) );
  AND2_X1 U19633 ( .A1(_03293__PTR4), .A2(_03292__PTR3), .ZN(_05177_) );
  AND2_X1 U19634 ( .A1(_03293__PTR6), .A2(_03292__PTR5), .ZN(_05178_) );
  AND2_X1 U19635 ( .A1(_02662__PTR40), .A2(_03292__PTR7), .ZN(_03292__PTR8) );
  AND2_X1 U19636 ( .A1(_02662__PTR42), .A2(_03292__PTR9), .ZN(_03292__PTR10) );
  AND2_X1 U19637 ( .A1(_02662__PTR44), .A2(_03292__PTR11), .ZN(_03292__PTR12) );
  AND2_X1 U19638 ( .A1(_02662__PTR46), .A2(_03292__PTR13), .ZN(_03292__PTR14) );
  AND2_X1 U19639 ( .A1(_02662__PTR48), .A2(_03292__PTR15), .ZN(_03292__PTR16) );
  AND2_X1 U19640 ( .A1(_02662__PTR50), .A2(_03292__PTR17), .ZN(_03292__PTR18) );
  AND2_X1 U19641 ( .A1(_02662__PTR52), .A2(_03292__PTR19), .ZN(_03292__PTR20) );
  AND2_X1 U19642 ( .A1(_02662__PTR54), .A2(_03292__PTR21), .ZN(_03292__PTR22) );
  AND2_X1 U19643 ( .A1(_02662__PTR56), .A2(_03292__PTR23), .ZN(_03292__PTR24) );
  AND2_X1 U19644 ( .A1(_02662__PTR58), .A2(_03292__PTR25), .ZN(_03292__PTR26) );
  AND2_X1 U19645 ( .A1(_02662__PTR60), .A2(_03292__PTR27), .ZN(_03292__PTR28) );
  AND2_X1 U19646 ( .A1(_02662__PTR62), .A2(_03292__PTR29), .ZN(_03292__PTR30) );
  OR2_X1 U19647 ( .A1(_03295__PTR1), .A2(_05146_), .ZN(_03292__PTR1) );
  OR2_X1 U19648 ( .A1(_03295__PTR3), .A2(_05147_), .ZN(_05179_) );
  OR2_X1 U19649 ( .A1(_03295__PTR5), .A2(_05148_), .ZN(_05180_) );
  OR2_X1 U19650 ( .A1(_03295__PTR7), .A2(_05149_), .ZN(_05181_) );
  OR2_X1 U19651 ( .A1(_05179_), .A2(_05150_), .ZN(_03292__PTR3) );
  OR2_X1 U19652 ( .A1(_05181_), .A2(_05151_), .ZN(_05182_) );
  OR2_X1 U19653 ( .A1(_05182_), .A2(_05152_), .ZN(_03292__PTR7) );
  OR2_X1 U19654 ( .A1(_05180_), .A2(_05175_), .ZN(_03292__PTR5) );
  OR2_X1 U19655 ( .A1(_03295__PTR2), .A2(_05176_), .ZN(_03292__PTR2) );
  OR2_X1 U19656 ( .A1(_03295__PTR4), .A2(_05177_), .ZN(_03292__PTR4) );
  OR2_X1 U19657 ( .A1(_03295__PTR6), .A2(_05178_), .ZN(_03292__PTR6) );
  AND2_X1 U19658 ( .A1(_02466__PTR7), .A2(_03213__PTR6), .ZN(_05280_) );
  AND2_X1 U19659 ( .A1(_05283_), .A2(_04830_), .ZN(_05281_) );
  AND2_X1 U19660 ( .A1(_05284_), .A2(_03214__PTR3), .ZN(_05282_) );
  AND2_X1 U19661 ( .A1(_02466__PTR3), .A2(_02466__PTR2), .ZN(_04820_) );
  AND2_X1 U19662 ( .A1(_02466__PTR5), .A2(_02466__PTR4), .ZN(_04823_) );
  AND2_X1 U19663 ( .A1(_02466__PTR7), .A2(_02466__PTR6), .ZN(_05283_) );
  AND2_X1 U19664 ( .A1(_05283_), .A2(_04823_), .ZN(_05284_) );
  AND2_X1 U19665 ( .A1(_02466__PTR4), .A2(_03214__PTR3), .ZN(_04827_) );
  OR2_X1 U19666 ( .A1(_03213__PTR5), .A2(_04818_), .ZN(_04830_) );
  OR2_X1 U19667 ( .A1(_03213__PTR7), .A2(_05280_), .ZN(_05285_) );
  OR2_X1 U19668 ( .A1(_04829_), .A2(_04820_), .ZN(_03214__PTR3) );
  OR2_X1 U19669 ( .A1(_05285_), .A2(_05281_), .ZN(_05286_) );
  OR2_X1 U19670 ( .A1(_05286_), .A2(_05282_), .ZN(_03424__PTR8) );
  OR2_X1 U19671 ( .A1(_04830_), .A2(_04826_), .ZN(_03214__PTR5) );
  AND2_X1 U19672 ( .A1(P3_P1_InstAddrPointer_PTR1), .A2(P3_P1_InstAddrPointer_PTR0), .ZN(_03288__PTR1) );
  AND2_X1 U19673 ( .A1(_05102_), .A2(_03288__PTR1), .ZN(_03288__PTR3) );
  AND2_X1 U19674 ( .A1(_05116_), .A2(_03288__PTR3), .ZN(_03288__PTR7) );
  AND2_X1 U19675 ( .A1(_05122_), .A2(_03288__PTR7), .ZN(_03288__PTR15) );
  AND2_X1 U19676 ( .A1(P3_P1_InstAddrPointer_PTR3), .A2(P3_P1_InstAddrPointer_PTR2), .ZN(_05102_) );
  AND2_X1 U19677 ( .A1(P3_P1_InstAddrPointer_PTR5), .A2(P3_P1_InstAddrPointer_PTR4), .ZN(_05103_) );
  AND2_X1 U19678 ( .A1(P3_P1_InstAddrPointer_PTR7), .A2(P3_P1_InstAddrPointer_PTR6), .ZN(_05104_) );
  AND2_X1 U19679 ( .A1(P3_P1_InstAddrPointer_PTR9), .A2(P3_P1_InstAddrPointer_PTR8), .ZN(_05105_) );
  AND2_X1 U19680 ( .A1(P3_P1_InstAddrPointer_PTR13), .A2(P3_P1_InstAddrPointer_PTR12), .ZN(_05107_) );
  AND2_X1 U19681 ( .A1(P3_P1_InstAddrPointer_PTR15), .A2(P3_P1_InstAddrPointer_PTR14), .ZN(_05108_) );
  AND2_X1 U19682 ( .A1(P3_P1_InstAddrPointer_PTR17), .A2(P3_P1_InstAddrPointer_PTR16), .ZN(_05109_) );
  AND2_X1 U19683 ( .A1(P3_P1_InstAddrPointer_PTR19), .A2(P3_P1_InstAddrPointer_PTR18), .ZN(_05110_) );
  AND2_X1 U19684 ( .A1(P3_P1_InstAddrPointer_PTR21), .A2(P3_P1_InstAddrPointer_PTR20), .ZN(_05111_) );
  AND2_X1 U19685 ( .A1(P3_P1_InstAddrPointer_PTR23), .A2(P3_P1_InstAddrPointer_PTR22), .ZN(_05112_) );
  AND2_X1 U19686 ( .A1(P3_P1_InstAddrPointer_PTR27), .A2(P3_P1_InstAddrPointer_PTR26), .ZN(_05114_) );
  AND2_X1 U19687 ( .A1(P3_P1_InstAddrPointer_PTR29), .A2(P3_P1_InstAddrPointer_PTR28), .ZN(_05115_) );
  AND2_X1 U19688 ( .A1(_05104_), .A2(_05103_), .ZN(_05116_) );
  AND2_X1 U19689 ( .A1(_05108_), .A2(_05107_), .ZN(_05118_) );
  AND2_X1 U19690 ( .A1(_05112_), .A2(_05111_), .ZN(_05120_) );
  AND2_X1 U19691 ( .A1(_05114_), .A2(_05113_), .ZN(_05121_) );
  AND2_X1 U19692 ( .A1(_05118_), .A2(_05117_), .ZN(_05122_) );
  AND2_X1 U19693 ( .A1(_05120_), .A2(_05119_), .ZN(_05123_) );
  AND2_X1 U19694 ( .A1(_05123_), .A2(_03288__PTR15), .ZN(_03288__PTR23) );
  AND2_X1 U19695 ( .A1(_05117_), .A2(_03288__PTR7), .ZN(_03288__PTR11) );
  AND2_X1 U19696 ( .A1(_05119_), .A2(_03288__PTR15), .ZN(_03288__PTR19) );
  AND2_X1 U19697 ( .A1(_05121_), .A2(_03288__PTR23), .ZN(_03288__PTR27) );
  AND2_X1 U19698 ( .A1(_05103_), .A2(_03288__PTR3), .ZN(_03288__PTR5) );
  AND2_X1 U19699 ( .A1(_05105_), .A2(_03288__PTR7), .ZN(_03288__PTR9) );
  AND2_X1 U19700 ( .A1(_05107_), .A2(_03288__PTR11), .ZN(_03288__PTR13) );
  AND2_X1 U19701 ( .A1(_05109_), .A2(_03288__PTR15), .ZN(_03288__PTR17) );
  AND2_X1 U19702 ( .A1(_05111_), .A2(_03288__PTR19), .ZN(_03288__PTR21) );
  AND2_X1 U19703 ( .A1(_05113_), .A2(_03288__PTR23), .ZN(_03288__PTR25) );
  AND2_X1 U19704 ( .A1(_05115_), .A2(_03288__PTR27), .ZN(_03288__PTR29) );
  AND2_X1 U19705 ( .A1(P3_P1_InstAddrPointer_PTR2), .A2(_03288__PTR1), .ZN(_03288__PTR2) );
  AND2_X1 U19706 ( .A1(P3_P1_InstAddrPointer_PTR4), .A2(_03288__PTR3), .ZN(_03288__PTR4) );
  AND2_X1 U19707 ( .A1(P3_P1_InstAddrPointer_PTR6), .A2(_03288__PTR5), .ZN(_03288__PTR6) );
  AND2_X1 U19708 ( .A1(P3_P1_InstAddrPointer_PTR8), .A2(_03288__PTR7), .ZN(_03288__PTR8) );
  AND2_X1 U19709 ( .A1(P3_P1_InstAddrPointer_PTR10), .A2(_03288__PTR9), .ZN(_03288__PTR10) );
  AND2_X1 U19710 ( .A1(P3_P1_InstAddrPointer_PTR12), .A2(_03288__PTR11), .ZN(_03288__PTR12) );
  AND2_X1 U19711 ( .A1(P3_P1_InstAddrPointer_PTR14), .A2(_03288__PTR13), .ZN(_03288__PTR14) );
  AND2_X1 U19712 ( .A1(P3_P1_InstAddrPointer_PTR16), .A2(_03288__PTR15), .ZN(_03288__PTR16) );
  AND2_X1 U19713 ( .A1(P3_P1_InstAddrPointer_PTR18), .A2(_03288__PTR17), .ZN(_03288__PTR18) );
  AND2_X1 U19714 ( .A1(P3_P1_InstAddrPointer_PTR20), .A2(_03288__PTR19), .ZN(_03288__PTR20) );
  AND2_X1 U19715 ( .A1(P3_P1_InstAddrPointer_PTR22), .A2(_03288__PTR21), .ZN(_03288__PTR22) );
  AND2_X1 U19716 ( .A1(P3_P1_InstAddrPointer_PTR24), .A2(_03288__PTR23), .ZN(_03288__PTR24) );
  AND2_X1 U19717 ( .A1(P3_P1_InstAddrPointer_PTR26), .A2(_03288__PTR25), .ZN(_03288__PTR26) );
  AND2_X1 U19718 ( .A1(P3_P1_InstAddrPointer_PTR28), .A2(_03288__PTR27), .ZN(_03288__PTR28) );
  AND2_X1 U19719 ( .A1(P3_P1_InstAddrPointer_PTR30), .A2(_03288__PTR29), .ZN(_03288__PTR30) );
  AND2_X1 U19720 ( .A1(_03299__PTR1), .A2(_03427__PTR0), .ZN(_05287_) );
  AND2_X1 U19721 ( .A1(_03428__PTR3), .A2(_03430__PTR2), .ZN(_05288_) );
  AND2_X1 U19722 ( .A1(_03428__PTR5), .A2(_03430__PTR4), .ZN(_05289_) );
  AND2_X1 U19723 ( .A1(_03428__PTR7), .A2(_03430__PTR6), .ZN(_05290_) );
  AND2_X1 U19724 ( .A1(_03428__PTR9), .A2(_03430__PTR8), .ZN(_05291_) );
  AND2_X1 U19725 ( .A1(_03428__PTR11), .A2(_03430__PTR10), .ZN(_05292_) );
  AND2_X1 U19726 ( .A1(_03428__PTR13), .A2(_03430__PTR12), .ZN(_05293_) );
  AND2_X1 U19727 ( .A1(_03428__PTR15), .A2(_03430__PTR14), .ZN(_05294_) );
  AND2_X1 U19728 ( .A1(_03428__PTR17), .A2(_03430__PTR16), .ZN(_05295_) );
  AND2_X1 U19729 ( .A1(_03428__PTR19), .A2(_03430__PTR18), .ZN(_05296_) );
  AND2_X1 U19730 ( .A1(_03428__PTR21), .A2(_03430__PTR20), .ZN(_05297_) );
  AND2_X1 U19731 ( .A1(_03428__PTR23), .A2(_03430__PTR22), .ZN(_05298_) );
  AND2_X1 U19732 ( .A1(_03428__PTR25), .A2(_03430__PTR24), .ZN(_05299_) );
  AND2_X1 U19733 ( .A1(_03428__PTR27), .A2(_03430__PTR26), .ZN(_05300_) );
  AND2_X1 U19734 ( .A1(_03428__PTR29), .A2(_03430__PTR28), .ZN(_05301_) );
  AND2_X1 U19735 ( .A1(_05313_), .A2(_03427__PTR1), .ZN(_05302_) );
  AND2_X1 U19736 ( .A1(_05315_), .A2(_05362_), .ZN(_05303_) );
  AND2_X1 U19737 ( .A1(_05317_), .A2(_05364_), .ZN(_05304_) );
  AND2_X1 U19738 ( .A1(_05319_), .A2(_05366_), .ZN(_05305_) );
  AND2_X1 U19739 ( .A1(_05321_), .A2(_05368_), .ZN(_05306_) );
  AND2_X1 U19740 ( .A1(_05323_), .A2(_05370_), .ZN(_05307_) );
  AND2_X1 U19741 ( .A1(_05325_), .A2(_05372_), .ZN(_05308_) );
  AND2_X1 U19742 ( .A1(_05327_), .A2(_03427__PTR3), .ZN(_05309_) );
  AND2_X1 U19743 ( .A1(_05329_), .A2(_05376_), .ZN(_05310_) );
  AND2_X1 U19744 ( .A1(_05331_), .A2(_05378_), .ZN(_05311_) );
  AND2_X1 U19745 ( .A1(_05333_), .A2(_03427__PTR7), .ZN(_05312_) );
  AND2_X1 U19746 ( .A1(_03428__PTR3), .A2(_03428__PTR2), .ZN(_05313_) );
  AND2_X1 U19747 ( .A1(_03428__PTR5), .A2(_03428__PTR4), .ZN(_05314_) );
  AND2_X1 U19748 ( .A1(_03428__PTR7), .A2(_03428__PTR6), .ZN(_05315_) );
  AND2_X1 U19749 ( .A1(_03428__PTR9), .A2(_03428__PTR8), .ZN(_05316_) );
  AND2_X1 U19750 ( .A1(_03428__PTR11), .A2(_03428__PTR10), .ZN(_05317_) );
  AND2_X1 U19751 ( .A1(_03428__PTR13), .A2(_03428__PTR12), .ZN(_05318_) );
  AND2_X1 U19752 ( .A1(_03428__PTR15), .A2(_03428__PTR14), .ZN(_05319_) );
  AND2_X1 U19753 ( .A1(_03428__PTR17), .A2(_03428__PTR16), .ZN(_05320_) );
  AND2_X1 U19754 ( .A1(_03428__PTR19), .A2(_03428__PTR18), .ZN(_05321_) );
  AND2_X1 U19755 ( .A1(_03428__PTR21), .A2(_03428__PTR20), .ZN(_05322_) );
  AND2_X1 U19756 ( .A1(_03428__PTR23), .A2(_03428__PTR22), .ZN(_05323_) );
  AND2_X1 U19757 ( .A1(_03428__PTR25), .A2(_03428__PTR24), .ZN(_05324_) );
  AND2_X1 U19758 ( .A1(_03428__PTR27), .A2(_03428__PTR26), .ZN(_05325_) );
  AND2_X1 U19759 ( .A1(_03428__PTR29), .A2(_03428__PTR28), .ZN(_05326_) );
  AND2_X1 U19760 ( .A1(_05315_), .A2(_05314_), .ZN(_05327_) );
  AND2_X1 U19761 ( .A1(_05317_), .A2(_05316_), .ZN(_05328_) );
  AND2_X1 U19762 ( .A1(_05319_), .A2(_05318_), .ZN(_05329_) );
  AND2_X1 U19763 ( .A1(_05321_), .A2(_05320_), .ZN(_05330_) );
  AND2_X1 U19764 ( .A1(_05323_), .A2(_05322_), .ZN(_05331_) );
  AND2_X1 U19765 ( .A1(_05325_), .A2(_05324_), .ZN(_05332_) );
  AND2_X1 U19766 ( .A1(_05329_), .A2(_05328_), .ZN(_05333_) );
  AND2_X1 U19767 ( .A1(_05331_), .A2(_05330_), .ZN(_05334_) );
  AND2_X1 U19768 ( .A1(_05334_), .A2(_03427__PTR15), .ZN(_05335_) );
  AND2_X1 U19769 ( .A1(_05328_), .A2(_03427__PTR7), .ZN(_05336_) );
  AND2_X1 U19770 ( .A1(_05330_), .A2(_03427__PTR15), .ZN(_05337_) );
  AND2_X1 U19771 ( .A1(_05332_), .A2(_03427__PTR23), .ZN(_05338_) );
  AND2_X1 U19772 ( .A1(_05314_), .A2(_03427__PTR3), .ZN(_05339_) );
  AND2_X1 U19773 ( .A1(_05316_), .A2(_03427__PTR7), .ZN(_05340_) );
  AND2_X1 U19774 ( .A1(_05318_), .A2(_03427__PTR11), .ZN(_05341_) );
  AND2_X1 U19775 ( .A1(_05320_), .A2(_03427__PTR15), .ZN(_05342_) );
  AND2_X1 U19776 ( .A1(_05322_), .A2(_03427__PTR19), .ZN(_05343_) );
  AND2_X1 U19777 ( .A1(_05324_), .A2(_03427__PTR23), .ZN(_05344_) );
  AND2_X1 U19778 ( .A1(_05326_), .A2(_03427__PTR27), .ZN(_05345_) );
  AND2_X1 U19779 ( .A1(_03428__PTR2), .A2(_03427__PTR1), .ZN(_05346_) );
  AND2_X1 U19780 ( .A1(_03428__PTR4), .A2(_03427__PTR3), .ZN(_05347_) );
  AND2_X1 U19781 ( .A1(_03428__PTR6), .A2(_03427__PTR5), .ZN(_05348_) );
  AND2_X1 U19782 ( .A1(_03428__PTR8), .A2(_03427__PTR7), .ZN(_05349_) );
  AND2_X1 U19783 ( .A1(_03428__PTR10), .A2(_03427__PTR9), .ZN(_05350_) );
  AND2_X1 U19784 ( .A1(_03428__PTR12), .A2(_03427__PTR11), .ZN(_05351_) );
  AND2_X1 U19785 ( .A1(_03428__PTR14), .A2(_03427__PTR13), .ZN(_05352_) );
  AND2_X1 U19786 ( .A1(_03428__PTR16), .A2(_03427__PTR15), .ZN(_05353_) );
  AND2_X1 U19787 ( .A1(_03428__PTR18), .A2(_03427__PTR17), .ZN(_05354_) );
  AND2_X1 U19788 ( .A1(_03428__PTR20), .A2(_03427__PTR19), .ZN(_05355_) );
  AND2_X1 U19789 ( .A1(_03428__PTR22), .A2(_03427__PTR21), .ZN(_05356_) );
  AND2_X1 U19790 ( .A1(_03428__PTR24), .A2(_03427__PTR23), .ZN(_05357_) );
  AND2_X1 U19791 ( .A1(_03428__PTR26), .A2(_03427__PTR25), .ZN(_05358_) );
  AND2_X1 U19792 ( .A1(_03428__PTR28), .A2(_03427__PTR27), .ZN(_05359_) );
  AND2_X1 U19793 ( .A1(_03428__PTR30), .A2(_03427__PTR29), .ZN(_05360_) );
  OR2_X1 U19794 ( .A1(_03298__PTR0), .A2(_03299__PTR0), .ZN(_03427__PTR0) );
  OR2_X1 U19795 ( .A1(_03301__PTR1), .A2(_05287_), .ZN(_03427__PTR1) );
  OR2_X1 U19796 ( .A1(_03430__PTR3), .A2(_05288_), .ZN(_05361_) );
  OR2_X1 U19797 ( .A1(_03430__PTR5), .A2(_05289_), .ZN(_05362_) );
  OR2_X1 U19798 ( .A1(_03430__PTR7), .A2(_05290_), .ZN(_05363_) );
  OR2_X1 U19799 ( .A1(_03430__PTR9), .A2(_05291_), .ZN(_05364_) );
  OR2_X1 U19800 ( .A1(_03430__PTR11), .A2(_05292_), .ZN(_05365_) );
  OR2_X1 U19801 ( .A1(_03430__PTR13), .A2(_05293_), .ZN(_05366_) );
  OR2_X1 U19802 ( .A1(_03430__PTR15), .A2(_05294_), .ZN(_05367_) );
  OR2_X1 U19803 ( .A1(_03430__PTR17), .A2(_05295_), .ZN(_05368_) );
  OR2_X1 U19804 ( .A1(_03430__PTR19), .A2(_05296_), .ZN(_05369_) );
  OR2_X1 U19805 ( .A1(_03430__PTR21), .A2(_05297_), .ZN(_05370_) );
  OR2_X1 U19806 ( .A1(_03430__PTR23), .A2(_05298_), .ZN(_05371_) );
  OR2_X1 U19807 ( .A1(_03430__PTR25), .A2(_05299_), .ZN(_05372_) );
  OR2_X1 U19808 ( .A1(_03430__PTR27), .A2(_05300_), .ZN(_05373_) );
  OR2_X1 U19809 ( .A1(_03430__PTR29), .A2(_05301_), .ZN(_05374_) );
  OR2_X1 U19810 ( .A1(_05361_), .A2(_05302_), .ZN(_03427__PTR3) );
  OR2_X1 U19811 ( .A1(_05363_), .A2(_05303_), .ZN(_05375_) );
  OR2_X1 U19812 ( .A1(_05365_), .A2(_05304_), .ZN(_05376_) );
  OR2_X1 U19813 ( .A1(_05367_), .A2(_05305_), .ZN(_05377_) );
  OR2_X1 U19814 ( .A1(_05369_), .A2(_05306_), .ZN(_05378_) );
  OR2_X1 U19815 ( .A1(_05371_), .A2(_05307_), .ZN(_05379_) );
  OR2_X1 U19816 ( .A1(_05373_), .A2(_05308_), .ZN(_05380_) );
  OR2_X1 U19817 ( .A1(_05375_), .A2(_05309_), .ZN(_03427__PTR7) );
  OR2_X1 U19818 ( .A1(_05377_), .A2(_05310_), .ZN(_05381_) );
  OR2_X1 U19819 ( .A1(_05379_), .A2(_05311_), .ZN(_05382_) );
  OR2_X1 U19820 ( .A1(_05381_), .A2(_05312_), .ZN(_03427__PTR15) );
  OR2_X1 U19821 ( .A1(_05382_), .A2(_05335_), .ZN(_03427__PTR23) );
  OR2_X1 U19822 ( .A1(_05376_), .A2(_05336_), .ZN(_03427__PTR11) );
  OR2_X1 U19823 ( .A1(_05378_), .A2(_05337_), .ZN(_03427__PTR19) );
  OR2_X1 U19824 ( .A1(_05380_), .A2(_05338_), .ZN(_03427__PTR27) );
  OR2_X1 U19825 ( .A1(_05362_), .A2(_05339_), .ZN(_03427__PTR5) );
  OR2_X1 U19826 ( .A1(_05364_), .A2(_05340_), .ZN(_03427__PTR9) );
  OR2_X1 U19827 ( .A1(_05366_), .A2(_05341_), .ZN(_03427__PTR13) );
  OR2_X1 U19828 ( .A1(_05368_), .A2(_05342_), .ZN(_03427__PTR17) );
  OR2_X1 U19829 ( .A1(_05370_), .A2(_05343_), .ZN(_03427__PTR21) );
  OR2_X1 U19830 ( .A1(_05372_), .A2(_05344_), .ZN(_03427__PTR25) );
  OR2_X1 U19831 ( .A1(_05374_), .A2(_05345_), .ZN(_03427__PTR29) );
  OR2_X1 U19832 ( .A1(_03430__PTR2), .A2(_05346_), .ZN(_03427__PTR2) );
  OR2_X1 U19833 ( .A1(_03430__PTR4), .A2(_05347_), .ZN(_03427__PTR4) );
  OR2_X1 U19834 ( .A1(_03430__PTR6), .A2(_05348_), .ZN(_03427__PTR6) );
  OR2_X1 U19835 ( .A1(_03430__PTR8), .A2(_05349_), .ZN(_03427__PTR8) );
  OR2_X1 U19836 ( .A1(_03430__PTR10), .A2(_05350_), .ZN(_03427__PTR10) );
  OR2_X1 U19837 ( .A1(_03430__PTR12), .A2(_05351_), .ZN(_03427__PTR12) );
  OR2_X1 U19838 ( .A1(_03430__PTR14), .A2(_05352_), .ZN(_03427__PTR14) );
  OR2_X1 U19839 ( .A1(_03430__PTR16), .A2(_05353_), .ZN(_03427__PTR16) );
  OR2_X1 U19840 ( .A1(_03430__PTR18), .A2(_05354_), .ZN(_03427__PTR18) );
  OR2_X1 U19841 ( .A1(_03430__PTR20), .A2(_05355_), .ZN(_03427__PTR20) );
  OR2_X1 U19842 ( .A1(_03430__PTR22), .A2(_05356_), .ZN(_03427__PTR22) );
  OR2_X1 U19843 ( .A1(_03430__PTR24), .A2(_05357_), .ZN(_03427__PTR24) );
  OR2_X1 U19844 ( .A1(_03430__PTR26), .A2(_05358_), .ZN(_03427__PTR26) );
  OR2_X1 U19845 ( .A1(_03430__PTR28), .A2(_05359_), .ZN(_03427__PTR28) );
  OR2_X1 U19846 ( .A1(_03430__PTR30), .A2(_05360_), .ZN(_03427__PTR30) );
  AND2_X1 U19847 ( .A1(_02466__PTR3), .A2(_03213__PTR2), .ZN(_04817_) );
  AND2_X1 U19848 ( .A1(_02466__PTR5), .A2(_03213__PTR4), .ZN(_04818_) );
  AND2_X1 U19849 ( .A1(_03213__PTR7), .A2(_03213__PTR6), .ZN(_04819_) );
  AND2_X1 U19850 ( .A1(_04824_), .A2(_04830_), .ZN(_04821_) );
  AND2_X1 U19851 ( .A1(_04825_), .A2(_03214__PTR3), .ZN(_04822_) );
  AND2_X1 U19852 ( .A1(_03213__PTR7), .A2(_02466__PTR6), .ZN(_04824_) );
  AND2_X1 U19853 ( .A1(_04824_), .A2(_04823_), .ZN(_04825_) );
  AND2_X1 U19854 ( .A1(_04823_), .A2(_03214__PTR3), .ZN(_04826_) );
  AND2_X1 U19855 ( .A1(_02466__PTR6), .A2(_03214__PTR5), .ZN(_04828_) );
  OR2_X1 U19856 ( .A1(_03213__PTR3), .A2(_04817_), .ZN(_04829_) );
  OR2_X1 U19857 ( .A1(_04819_), .A2(_04821_), .ZN(_04831_) );
  OR2_X1 U19858 ( .A1(_04831_), .A2(_04822_), .ZN(_03214__PTR7) );
  OR2_X1 U19859 ( .A1(_03213__PTR4), .A2(_04827_), .ZN(_03214__PTR4) );
  OR2_X1 U19860 ( .A1(_03213__PTR6), .A2(_04828_), .ZN(_03214__PTR6) );
  AND2_X1 U19861 ( .A1(_01266__PTR2), .A2(_03209__PTR3), .ZN(_04816_) );
  OR2_X1 U19862 ( .A1(_03206__PTR5), .A2(_04816_), .ZN(_03209__PTR5) );
  AND2_X1 U19863 ( .A1(P3_P1_InstQueueRd_Addr_PTR2), .A2(_03240__PTR1), .ZN(_03240__PTR2) );
  AND2_X1 U19864 ( .A1(P3_P1_InstQueueRd_Addr_PTR4), .A2(_03240__PTR3), .ZN(_03289__PTR4) );
  AND2_X1 U19865 ( .A1(P3_P1_PhyAddrPointer_PTR2), .A2(P3_P1_PhyAddrPointer_PTR1), .ZN(_03287__PTR1) );
  AND2_X1 U19866 ( .A1(_05080_), .A2(_03287__PTR1), .ZN(_03287__PTR3) );
  AND2_X1 U19867 ( .A1(_05094_), .A2(_03287__PTR3), .ZN(_03287__PTR7) );
  AND2_X1 U19868 ( .A1(_05100_), .A2(_03287__PTR7), .ZN(_03287__PTR15) );
  AND2_X1 U19869 ( .A1(P3_P1_PhyAddrPointer_PTR4), .A2(P3_P1_PhyAddrPointer_PTR3), .ZN(_05080_) );
  AND2_X1 U19870 ( .A1(P3_P1_PhyAddrPointer_PTR6), .A2(P3_P1_PhyAddrPointer_PTR5), .ZN(_05081_) );
  AND2_X1 U19871 ( .A1(P3_P1_PhyAddrPointer_PTR8), .A2(P3_P1_PhyAddrPointer_PTR7), .ZN(_05082_) );
  AND2_X1 U19872 ( .A1(P3_P1_PhyAddrPointer_PTR10), .A2(P3_P1_PhyAddrPointer_PTR9), .ZN(_05083_) );
  AND2_X1 U19873 ( .A1(P3_P1_PhyAddrPointer_PTR12), .A2(P3_P1_PhyAddrPointer_PTR11), .ZN(_05084_) );
  AND2_X1 U19874 ( .A1(P3_P1_PhyAddrPointer_PTR14), .A2(P3_P1_PhyAddrPointer_PTR13), .ZN(_05085_) );
  AND2_X1 U19875 ( .A1(P3_P1_PhyAddrPointer_PTR16), .A2(P3_P1_PhyAddrPointer_PTR15), .ZN(_05086_) );
  AND2_X1 U19876 ( .A1(P3_P1_PhyAddrPointer_PTR18), .A2(P3_P1_PhyAddrPointer_PTR17), .ZN(_05087_) );
  AND2_X1 U19877 ( .A1(P3_P1_PhyAddrPointer_PTR20), .A2(P3_P1_PhyAddrPointer_PTR19), .ZN(_05088_) );
  AND2_X1 U19878 ( .A1(P3_P1_PhyAddrPointer_PTR22), .A2(P3_P1_PhyAddrPointer_PTR21), .ZN(_05089_) );
  AND2_X1 U19879 ( .A1(P3_P1_PhyAddrPointer_PTR24), .A2(P3_P1_PhyAddrPointer_PTR23), .ZN(_05090_) );
  AND2_X1 U19880 ( .A1(P3_P1_PhyAddrPointer_PTR26), .A2(P3_P1_PhyAddrPointer_PTR25), .ZN(_05091_) );
  AND2_X1 U19881 ( .A1(P3_P1_PhyAddrPointer_PTR28), .A2(P3_P1_PhyAddrPointer_PTR27), .ZN(_05092_) );
  AND2_X1 U19882 ( .A1(P3_P1_PhyAddrPointer_PTR30), .A2(P3_P1_PhyAddrPointer_PTR29), .ZN(_05093_) );
  AND2_X1 U19883 ( .A1(_05082_), .A2(_05081_), .ZN(_05094_) );
  AND2_X1 U19884 ( .A1(_05084_), .A2(_05083_), .ZN(_05095_) );
  AND2_X1 U19885 ( .A1(_05086_), .A2(_05085_), .ZN(_05096_) );
  AND2_X1 U19886 ( .A1(_05088_), .A2(_05087_), .ZN(_05097_) );
  AND2_X1 U19887 ( .A1(_05090_), .A2(_05089_), .ZN(_05098_) );
  AND2_X1 U19888 ( .A1(_05092_), .A2(_05091_), .ZN(_05099_) );
  AND2_X1 U19889 ( .A1(_05096_), .A2(_05095_), .ZN(_05100_) );
  AND2_X1 U19890 ( .A1(_05098_), .A2(_05097_), .ZN(_05101_) );
  AND2_X1 U19891 ( .A1(_05101_), .A2(_03287__PTR15), .ZN(_03287__PTR23) );
  AND2_X1 U19892 ( .A1(_05095_), .A2(_03287__PTR7), .ZN(_03287__PTR11) );
  AND2_X1 U19893 ( .A1(_05097_), .A2(_03287__PTR15), .ZN(_03287__PTR19) );
  AND2_X1 U19894 ( .A1(_05099_), .A2(_03287__PTR23), .ZN(_03287__PTR27) );
  AND2_X1 U19895 ( .A1(_05081_), .A2(_03287__PTR3), .ZN(_03287__PTR5) );
  AND2_X1 U19896 ( .A1(_05083_), .A2(_03287__PTR7), .ZN(_03287__PTR9) );
  AND2_X1 U19897 ( .A1(_05085_), .A2(_03287__PTR11), .ZN(_03287__PTR13) );
  AND2_X1 U19898 ( .A1(_05087_), .A2(_03287__PTR15), .ZN(_03287__PTR17) );
  AND2_X1 U19899 ( .A1(_05089_), .A2(_03287__PTR19), .ZN(_03287__PTR21) );
  AND2_X1 U19900 ( .A1(_05091_), .A2(_03287__PTR23), .ZN(_03287__PTR25) );
  AND2_X1 U19901 ( .A1(_05093_), .A2(_03287__PTR27), .ZN(_03287__PTR29) );
  AND2_X1 U19902 ( .A1(P3_P1_PhyAddrPointer_PTR3), .A2(_03287__PTR1), .ZN(_03287__PTR2) );
  AND2_X1 U19903 ( .A1(P3_P1_PhyAddrPointer_PTR5), .A2(_03287__PTR3), .ZN(_03287__PTR4) );
  AND2_X1 U19904 ( .A1(P3_P1_PhyAddrPointer_PTR7), .A2(_03287__PTR5), .ZN(_03287__PTR6) );
  AND2_X1 U19905 ( .A1(P3_P1_PhyAddrPointer_PTR9), .A2(_03287__PTR7), .ZN(_03287__PTR8) );
  AND2_X1 U19906 ( .A1(P3_P1_PhyAddrPointer_PTR11), .A2(_03287__PTR9), .ZN(_03287__PTR10) );
  AND2_X1 U19907 ( .A1(P3_P1_PhyAddrPointer_PTR13), .A2(_03287__PTR11), .ZN(_03287__PTR12) );
  AND2_X1 U19908 ( .A1(P3_P1_PhyAddrPointer_PTR15), .A2(_03287__PTR13), .ZN(_03287__PTR14) );
  AND2_X1 U19909 ( .A1(P3_P1_PhyAddrPointer_PTR17), .A2(_03287__PTR15), .ZN(_03287__PTR16) );
  AND2_X1 U19910 ( .A1(P3_P1_PhyAddrPointer_PTR19), .A2(_03287__PTR17), .ZN(_03287__PTR18) );
  AND2_X1 U19911 ( .A1(P3_P1_PhyAddrPointer_PTR21), .A2(_03287__PTR19), .ZN(_03287__PTR20) );
  AND2_X1 U19912 ( .A1(P3_P1_PhyAddrPointer_PTR23), .A2(_03287__PTR21), .ZN(_03287__PTR22) );
  AND2_X1 U19913 ( .A1(P3_P1_PhyAddrPointer_PTR25), .A2(_03287__PTR23), .ZN(_03287__PTR24) );
  AND2_X1 U19914 ( .A1(P3_P1_PhyAddrPointer_PTR27), .A2(_03287__PTR25), .ZN(_03287__PTR26) );
  AND2_X1 U19915 ( .A1(P3_P1_PhyAddrPointer_PTR29), .A2(_03287__PTR27), .ZN(_03287__PTR28) );
  AND2_X1 U19916 ( .A1(P3_P1_PhyAddrPointer_PTR1), .A2(_03205__PTR0), .ZN(_03435__PTR1) );
  AND2_X1 U19917 ( .A1(_04751_), .A2(_03435__PTR1), .ZN(_03435__PTR3) );
  AND2_X1 U19918 ( .A1(_04780_), .A2(_03435__PTR3), .ZN(_03435__PTR7) );
  AND2_X1 U19919 ( .A1(_04787_), .A2(_03435__PTR7), .ZN(_03435__PTR15) );
  AND2_X1 U19920 ( .A1(_03205__PTR7), .A2(_03205__PTR6), .ZN(_04767_) );
  AND2_X1 U19921 ( .A1(_03205__PTR9), .A2(_03205__PTR8), .ZN(_04768_) );
  AND2_X1 U19922 ( .A1(_03205__PTR11), .A2(_03205__PTR10), .ZN(_04769_) );
  AND2_X1 U19923 ( .A1(_03205__PTR13), .A2(_03205__PTR12), .ZN(_04770_) );
  AND2_X1 U19924 ( .A1(_03205__PTR15), .A2(_03205__PTR14), .ZN(_04771_) );
  AND2_X1 U19925 ( .A1(_03205__PTR17), .A2(_03205__PTR16), .ZN(_04772_) );
  AND2_X1 U19926 ( .A1(_03205__PTR19), .A2(_03205__PTR18), .ZN(_04773_) );
  AND2_X1 U19927 ( .A1(_03205__PTR21), .A2(_03205__PTR20), .ZN(_04774_) );
  AND2_X1 U19928 ( .A1(_03205__PTR23), .A2(_03205__PTR22), .ZN(_04775_) );
  AND2_X1 U19929 ( .A1(_03205__PTR25), .A2(_03205__PTR24), .ZN(_04776_) );
  AND2_X1 U19930 ( .A1(_04788_), .A2(_03435__PTR15), .ZN(_03435__PTR23) );
  AND2_X1 U19931 ( .A1(_04781_), .A2(_03435__PTR7), .ZN(_03435__PTR11) );
  AND2_X1 U19932 ( .A1(_04783_), .A2(_03435__PTR15), .ZN(_03435__PTR19) );
  AND2_X1 U19933 ( .A1(_04785_), .A2(_03435__PTR23), .ZN(_03435__PTR27) );
  AND2_X1 U19934 ( .A1(_04766_), .A2(_03435__PTR3), .ZN(_03435__PTR5) );
  AND2_X1 U19935 ( .A1(_04768_), .A2(_03435__PTR7), .ZN(_03435__PTR9) );
  AND2_X1 U19936 ( .A1(_04770_), .A2(_03435__PTR11), .ZN(_03435__PTR13) );
  AND2_X1 U19937 ( .A1(_04772_), .A2(_03435__PTR15), .ZN(_03435__PTR17) );
  AND2_X1 U19938 ( .A1(_04774_), .A2(_03435__PTR19), .ZN(_03435__PTR21) );
  AND2_X1 U19939 ( .A1(_04776_), .A2(_03435__PTR23), .ZN(_03435__PTR25) );
  AND2_X1 U19940 ( .A1(_04778_), .A2(_03435__PTR27), .ZN(_03435__PTR29) );
  AND2_X1 U19941 ( .A1(_03205__PTR2), .A2(_03435__PTR1), .ZN(_03435__PTR2) );
  AND2_X1 U19942 ( .A1(_03205__PTR4), .A2(_03435__PTR3), .ZN(_03435__PTR4) );
  AND2_X1 U19943 ( .A1(_03205__PTR6), .A2(_03435__PTR5), .ZN(_03435__PTR6) );
  AND2_X1 U19944 ( .A1(_03205__PTR8), .A2(_03435__PTR7), .ZN(_03435__PTR8) );
  AND2_X1 U19945 ( .A1(_03205__PTR10), .A2(_03435__PTR9), .ZN(_03435__PTR10) );
  AND2_X1 U19946 ( .A1(_03205__PTR12), .A2(_03435__PTR11), .ZN(_03435__PTR12) );
  AND2_X1 U19947 ( .A1(_03205__PTR14), .A2(_03435__PTR13), .ZN(_03435__PTR14) );
  AND2_X1 U19948 ( .A1(_03205__PTR16), .A2(_03435__PTR15), .ZN(_03435__PTR16) );
  AND2_X1 U19949 ( .A1(_03205__PTR18), .A2(_03435__PTR17), .ZN(_03435__PTR18) );
  AND2_X1 U19950 ( .A1(_03205__PTR20), .A2(_03435__PTR19), .ZN(_03435__PTR20) );
  AND2_X1 U19951 ( .A1(_03205__PTR22), .A2(_03435__PTR21), .ZN(_03435__PTR22) );
  AND2_X1 U19952 ( .A1(_03205__PTR24), .A2(_03435__PTR23), .ZN(_03435__PTR24) );
  AND2_X1 U19953 ( .A1(_03205__PTR26), .A2(_03435__PTR25), .ZN(_03435__PTR26) );
  AND2_X1 U19954 ( .A1(_03205__PTR28), .A2(_03435__PTR27), .ZN(_03435__PTR28) );
  AND2_X1 U19955 ( .A1(_03205__PTR30), .A2(_03435__PTR29), .ZN(_03435__PTR30) );
  AND2_X1 U19956 ( .A1(_03205__PTR3), .A2(_02473__PTR130), .ZN(_04736_) );
  AND2_X1 U19957 ( .A1(_03205__PTR5), .A2(_02473__PTR132), .ZN(_04737_) );
  AND2_X1 U19958 ( .A1(_03205__PTR7), .A2(_02473__PTR134), .ZN(_04738_) );
  AND2_X1 U19959 ( .A1(_03205__PTR9), .A2(_02473__PTR136), .ZN(_04739_) );
  AND2_X1 U19960 ( .A1(_03205__PTR11), .A2(_02473__PTR138), .ZN(_04740_) );
  AND2_X1 U19961 ( .A1(_03205__PTR13), .A2(_02473__PTR140), .ZN(_04741_) );
  AND2_X1 U19962 ( .A1(_03205__PTR15), .A2(_02473__PTR142), .ZN(_04742_) );
  AND2_X1 U19963 ( .A1(_03205__PTR17), .A2(_02473__PTR144), .ZN(_04743_) );
  AND2_X1 U19964 ( .A1(_03205__PTR19), .A2(_02473__PTR146), .ZN(_04744_) );
  AND2_X1 U19965 ( .A1(_03205__PTR21), .A2(_02473__PTR148), .ZN(_04745_) );
  AND2_X1 U19966 ( .A1(_03205__PTR23), .A2(_02473__PTR150), .ZN(_04746_) );
  AND2_X1 U19967 ( .A1(_03205__PTR25), .A2(_02473__PTR152), .ZN(_04747_) );
  AND2_X1 U19968 ( .A1(_03205__PTR27), .A2(_02473__PTR154), .ZN(_04748_) );
  AND2_X1 U19969 ( .A1(_03205__PTR29), .A2(_02473__PTR156), .ZN(_04749_) );
  AND2_X1 U19970 ( .A1(_03203__PTR31), .A2(_02473__PTR158), .ZN(_04750_) );
  AND2_X1 U19971 ( .A1(_04767_), .A2(_04792_), .ZN(_04752_) );
  AND2_X1 U19972 ( .A1(_04769_), .A2(_04794_), .ZN(_04753_) );
  AND2_X1 U19973 ( .A1(_04771_), .A2(_04796_), .ZN(_04754_) );
  AND2_X1 U19974 ( .A1(_04773_), .A2(_04798_), .ZN(_04755_) );
  AND2_X1 U19975 ( .A1(_04775_), .A2(_04800_), .ZN(_04756_) );
  AND2_X1 U19976 ( .A1(_04777_), .A2(_04802_), .ZN(_04757_) );
  AND2_X1 U19977 ( .A1(_04779_), .A2(_04804_), .ZN(_04758_) );
  AND2_X1 U19978 ( .A1(_04780_), .A2(_03204__PTR3), .ZN(_04759_) );
  AND2_X1 U19979 ( .A1(_04782_), .A2(_04806_), .ZN(_04760_) );
  AND2_X1 U19980 ( .A1(_04784_), .A2(_04808_), .ZN(_04761_) );
  AND2_X1 U19981 ( .A1(_04786_), .A2(_04810_), .ZN(_04762_) );
  AND2_X1 U19982 ( .A1(_04787_), .A2(_03204__PTR7), .ZN(_04763_) );
  AND2_X1 U19983 ( .A1(_04789_), .A2(_04813_), .ZN(_04764_) );
  AND2_X1 U19984 ( .A1(_04790_), .A2(_03204__PTR15), .ZN(_04765_) );
  AND2_X1 U19985 ( .A1(_03205__PTR3), .A2(_03205__PTR2), .ZN(_04751_) );
  AND2_X1 U19986 ( .A1(_03205__PTR5), .A2(_03205__PTR4), .ZN(_04766_) );
  AND2_X1 U19987 ( .A1(_03205__PTR27), .A2(_03205__PTR26), .ZN(_04777_) );
  AND2_X1 U19988 ( .A1(_03205__PTR29), .A2(_03205__PTR28), .ZN(_04778_) );
  AND2_X1 U19989 ( .A1(_03203__PTR31), .A2(_03205__PTR30), .ZN(_04779_) );
  AND2_X1 U19990 ( .A1(_04767_), .A2(_04766_), .ZN(_04780_) );
  AND2_X1 U19991 ( .A1(_04769_), .A2(_04768_), .ZN(_04781_) );
  AND2_X1 U19992 ( .A1(_04771_), .A2(_04770_), .ZN(_04782_) );
  AND2_X1 U19993 ( .A1(_04773_), .A2(_04772_), .ZN(_04783_) );
  AND2_X1 U19994 ( .A1(_04775_), .A2(_04774_), .ZN(_04784_) );
  AND2_X1 U19995 ( .A1(_04777_), .A2(_04776_), .ZN(_04785_) );
  AND2_X1 U19996 ( .A1(_04779_), .A2(_04778_), .ZN(_04786_) );
  AND2_X1 U19997 ( .A1(_04782_), .A2(_04781_), .ZN(_04787_) );
  AND2_X1 U19998 ( .A1(_04784_), .A2(_04783_), .ZN(_04788_) );
  AND2_X1 U19999 ( .A1(_04786_), .A2(_04785_), .ZN(_04789_) );
  AND2_X1 U20000 ( .A1(_04789_), .A2(_04788_), .ZN(_04790_) );
  OR2_X1 U20001 ( .A1(_02473__PTR131), .A2(_04736_), .ZN(_04791_) );
  OR2_X1 U20002 ( .A1(_02473__PTR133), .A2(_04737_), .ZN(_04792_) );
  OR2_X1 U20003 ( .A1(_02473__PTR135), .A2(_04738_), .ZN(_04793_) );
  OR2_X1 U20004 ( .A1(_02473__PTR137), .A2(_04739_), .ZN(_04794_) );
  OR2_X1 U20005 ( .A1(_02473__PTR139), .A2(_04740_), .ZN(_04795_) );
  OR2_X1 U20006 ( .A1(_02473__PTR141), .A2(_04741_), .ZN(_04796_) );
  OR2_X1 U20007 ( .A1(_02473__PTR143), .A2(_04742_), .ZN(_04797_) );
  OR2_X1 U20008 ( .A1(_02473__PTR145), .A2(_04743_), .ZN(_04798_) );
  OR2_X1 U20009 ( .A1(_02473__PTR147), .A2(_04744_), .ZN(_04799_) );
  OR2_X1 U20010 ( .A1(_02473__PTR149), .A2(_04745_), .ZN(_04800_) );
  OR2_X1 U20011 ( .A1(_02473__PTR151), .A2(_04746_), .ZN(_04801_) );
  OR2_X1 U20012 ( .A1(_02473__PTR153), .A2(_04747_), .ZN(_04802_) );
  OR2_X1 U20013 ( .A1(_02473__PTR155), .A2(_04748_), .ZN(_04803_) );
  OR2_X1 U20014 ( .A1(_02473__PTR157), .A2(_04749_), .ZN(_04804_) );
  OR2_X1 U20015 ( .A1(_04791_), .A2(_04751_), .ZN(_03204__PTR3) );
  OR2_X1 U20016 ( .A1(_04793_), .A2(_04752_), .ZN(_04805_) );
  OR2_X1 U20017 ( .A1(_04795_), .A2(_04753_), .ZN(_04806_) );
  OR2_X1 U20018 ( .A1(_04797_), .A2(_04754_), .ZN(_04807_) );
  OR2_X1 U20019 ( .A1(_04799_), .A2(_04755_), .ZN(_04808_) );
  OR2_X1 U20020 ( .A1(_04801_), .A2(_04756_), .ZN(_04809_) );
  OR2_X1 U20021 ( .A1(_04803_), .A2(_04757_), .ZN(_04810_) );
  OR2_X1 U20022 ( .A1(_04750_), .A2(_04758_), .ZN(_04811_) );
  OR2_X1 U20023 ( .A1(_04805_), .A2(_04759_), .ZN(_03204__PTR7) );
  OR2_X1 U20024 ( .A1(_04807_), .A2(_04760_), .ZN(_04812_) );
  OR2_X1 U20025 ( .A1(_04809_), .A2(_04761_), .ZN(_04813_) );
  OR2_X1 U20026 ( .A1(_04811_), .A2(_04762_), .ZN(_04814_) );
  OR2_X1 U20027 ( .A1(_04812_), .A2(_04763_), .ZN(_03204__PTR15) );
  OR2_X1 U20028 ( .A1(_04814_), .A2(_04764_), .ZN(_04815_) );
  OR2_X1 U20029 ( .A1(_04815_), .A2(_04765_), .ZN(_03204__PTR31) );
  AND2_X1 U20030 ( .A1(P3_P1_PhyAddrPointer_PTR3), .A2(P3_P1_PhyAddrPointer_PTR2), .ZN(_03284__PTR1) );
  AND2_X1 U20031 ( .A1(_05059_), .A2(_03284__PTR1), .ZN(_03284__PTR3) );
  AND2_X1 U20032 ( .A1(_05072_), .A2(_03284__PTR3), .ZN(_03284__PTR7) );
  AND2_X1 U20033 ( .A1(_05078_), .A2(_03284__PTR7), .ZN(_03284__PTR15) );
  AND2_X1 U20034 ( .A1(P3_P1_PhyAddrPointer_PTR5), .A2(P3_P1_PhyAddrPointer_PTR4), .ZN(_05059_) );
  AND2_X1 U20035 ( .A1(P3_P1_PhyAddrPointer_PTR7), .A2(P3_P1_PhyAddrPointer_PTR6), .ZN(_05060_) );
  AND2_X1 U20036 ( .A1(P3_P1_PhyAddrPointer_PTR9), .A2(P3_P1_PhyAddrPointer_PTR8), .ZN(_05061_) );
  AND2_X1 U20037 ( .A1(P3_P1_PhyAddrPointer_PTR11), .A2(P3_P1_PhyAddrPointer_PTR10), .ZN(_05062_) );
  AND2_X1 U20038 ( .A1(P3_P1_PhyAddrPointer_PTR13), .A2(P3_P1_PhyAddrPointer_PTR12), .ZN(_05063_) );
  AND2_X1 U20039 ( .A1(P3_P1_PhyAddrPointer_PTR15), .A2(P3_P1_PhyAddrPointer_PTR14), .ZN(_05064_) );
  AND2_X1 U20040 ( .A1(P3_P1_PhyAddrPointer_PTR17), .A2(P3_P1_PhyAddrPointer_PTR16), .ZN(_05065_) );
  AND2_X1 U20041 ( .A1(P3_P1_PhyAddrPointer_PTR19), .A2(P3_P1_PhyAddrPointer_PTR18), .ZN(_05066_) );
  AND2_X1 U20042 ( .A1(P3_P1_PhyAddrPointer_PTR21), .A2(P3_P1_PhyAddrPointer_PTR20), .ZN(_05067_) );
  AND2_X1 U20043 ( .A1(P3_P1_PhyAddrPointer_PTR23), .A2(P3_P1_PhyAddrPointer_PTR22), .ZN(_05068_) );
  AND2_X1 U20044 ( .A1(P3_P1_PhyAddrPointer_PTR25), .A2(P3_P1_PhyAddrPointer_PTR24), .ZN(_05069_) );
  AND2_X1 U20045 ( .A1(P3_P1_PhyAddrPointer_PTR27), .A2(P3_P1_PhyAddrPointer_PTR26), .ZN(_05070_) );
  AND2_X1 U20046 ( .A1(P3_P1_PhyAddrPointer_PTR29), .A2(P3_P1_PhyAddrPointer_PTR28), .ZN(_05071_) );
  AND2_X1 U20047 ( .A1(_05061_), .A2(_05060_), .ZN(_05072_) );
  AND2_X1 U20048 ( .A1(_05063_), .A2(_05062_), .ZN(_05073_) );
  AND2_X1 U20049 ( .A1(_05065_), .A2(_05064_), .ZN(_05074_) );
  AND2_X1 U20050 ( .A1(_05067_), .A2(_05066_), .ZN(_05075_) );
  AND2_X1 U20051 ( .A1(_05069_), .A2(_05068_), .ZN(_05076_) );
  AND2_X1 U20052 ( .A1(_05071_), .A2(_05070_), .ZN(_05077_) );
  AND2_X1 U20053 ( .A1(_05074_), .A2(_05073_), .ZN(_05078_) );
  AND2_X1 U20054 ( .A1(_05076_), .A2(_05075_), .ZN(_05079_) );
  AND2_X1 U20055 ( .A1(_05079_), .A2(_03284__PTR15), .ZN(_03284__PTR23) );
  AND2_X1 U20056 ( .A1(_05073_), .A2(_03284__PTR7), .ZN(_03284__PTR11) );
  AND2_X1 U20057 ( .A1(_05075_), .A2(_03284__PTR15), .ZN(_03284__PTR19) );
  AND2_X1 U20058 ( .A1(_05077_), .A2(_03284__PTR23), .ZN(_03284__PTR27) );
  AND2_X1 U20059 ( .A1(_05060_), .A2(_03284__PTR3), .ZN(_03284__PTR5) );
  AND2_X1 U20060 ( .A1(_05062_), .A2(_03284__PTR7), .ZN(_03284__PTR9) );
  AND2_X1 U20061 ( .A1(_05064_), .A2(_03284__PTR11), .ZN(_03284__PTR13) );
  AND2_X1 U20062 ( .A1(_05066_), .A2(_03284__PTR15), .ZN(_03284__PTR17) );
  AND2_X1 U20063 ( .A1(_05068_), .A2(_03284__PTR19), .ZN(_03284__PTR21) );
  AND2_X1 U20064 ( .A1(_05070_), .A2(_03284__PTR23), .ZN(_03284__PTR25) );
  AND2_X1 U20065 ( .A1(P3_P1_PhyAddrPointer_PTR4), .A2(_03284__PTR1), .ZN(_03284__PTR2) );
  AND2_X1 U20066 ( .A1(P3_P1_PhyAddrPointer_PTR6), .A2(_03284__PTR3), .ZN(_03284__PTR4) );
  AND2_X1 U20067 ( .A1(P3_P1_PhyAddrPointer_PTR8), .A2(_03284__PTR5), .ZN(_03284__PTR6) );
  AND2_X1 U20068 ( .A1(P3_P1_PhyAddrPointer_PTR10), .A2(_03284__PTR7), .ZN(_03284__PTR8) );
  AND2_X1 U20069 ( .A1(P3_P1_PhyAddrPointer_PTR12), .A2(_03284__PTR9), .ZN(_03284__PTR10) );
  AND2_X1 U20070 ( .A1(P3_P1_PhyAddrPointer_PTR14), .A2(_03284__PTR11), .ZN(_03284__PTR12) );
  AND2_X1 U20071 ( .A1(P3_P1_PhyAddrPointer_PTR16), .A2(_03284__PTR13), .ZN(_03284__PTR14) );
  AND2_X1 U20072 ( .A1(P3_P1_PhyAddrPointer_PTR18), .A2(_03284__PTR15), .ZN(_03284__PTR16) );
  AND2_X1 U20073 ( .A1(P3_P1_PhyAddrPointer_PTR20), .A2(_03284__PTR17), .ZN(_03284__PTR18) );
  AND2_X1 U20074 ( .A1(P3_P1_PhyAddrPointer_PTR22), .A2(_03284__PTR19), .ZN(_03284__PTR20) );
  AND2_X1 U20075 ( .A1(P3_P1_PhyAddrPointer_PTR24), .A2(_03284__PTR21), .ZN(_03284__PTR22) );
  AND2_X1 U20076 ( .A1(P3_P1_PhyAddrPointer_PTR26), .A2(_03284__PTR23), .ZN(_03284__PTR24) );
  AND2_X1 U20077 ( .A1(P3_P1_PhyAddrPointer_PTR28), .A2(_03284__PTR25), .ZN(_03284__PTR26) );
  AND2_X1 U20078 ( .A1(P3_P1_PhyAddrPointer_PTR30), .A2(_03284__PTR27), .ZN(_03284__PTR28) );
  AND2_X1 U20079 ( .A1(P3_P1_InstQueueWr_Addr_PTR1), .A2(P3_P1_InstQueueWr_Addr_PTR0), .ZN(_03269__PTR1) );
  AND2_X1 U20080 ( .A1(P3_P1_InstQueueWr_Addr_PTR2), .A2(_03269__PTR1), .ZN(_03269__PTR2) );
  AND2_X1 U20081 ( .A1(_02418__PTR1), .A2(_02418__PTR0), .ZN(_03270__PTR1) );
  AND2_X1 U20082 ( .A1(_02418__PTR2), .A2(_03270__PTR1), .ZN(_03270__PTR2) );
  AND2_X1 U20083 ( .A1(_02420__PTR1), .A2(P3_P1_InstQueueWr_Addr_PTR0), .ZN(_03275__PTR1) );
  AND2_X1 U20084 ( .A1(_02420__PTR2), .A2(_03275__PTR1), .ZN(_03275__PTR2) );
  AND2_X1 U20085 ( .A1(_02422__PTR1), .A2(_02418__PTR0), .ZN(_03280__PTR1) );
  AND2_X1 U20086 ( .A1(_02422__PTR2), .A2(_03280__PTR1), .ZN(_03280__PTR2) );
  AND2_X1 U20087 ( .A1(buf2_PTR25), .A2(_03277__PTR0), .ZN(_03277__PTR1) );
  AND2_X1 U20088 ( .A1(_05036_), .A2(_03277__PTR1), .ZN(_03277__PTR3) );
  AND2_X1 U20089 ( .A1(_05037_), .A2(_03277__PTR3), .ZN(_03277__PTR5) );
  AND2_X1 U20090 ( .A1(buf2_PTR26), .A2(_03277__PTR1), .ZN(_03277__PTR2) );
  AND2_X1 U20091 ( .A1(buf2_PTR28), .A2(_03277__PTR3), .ZN(_03277__PTR4) );
  AND2_X1 U20092 ( .A1(buf2_PTR30), .A2(_03277__PTR5), .ZN(_03277__PTR6) );
  AND2_X1 U20093 ( .A1(buf2_PTR17), .A2(_03272__PTR0), .ZN(_03272__PTR1) );
  AND2_X1 U20094 ( .A1(_05034_), .A2(_03272__PTR1), .ZN(_03272__PTR3) );
  AND2_X1 U20095 ( .A1(buf2_PTR19), .A2(buf2_PTR18), .ZN(_05034_) );
  AND2_X1 U20096 ( .A1(buf2_PTR21), .A2(buf2_PTR20), .ZN(_05035_) );
  AND2_X1 U20097 ( .A1(buf2_PTR27), .A2(buf2_PTR26), .ZN(_05036_) );
  AND2_X1 U20098 ( .A1(buf2_PTR29), .A2(buf2_PTR28), .ZN(_05037_) );
  AND2_X1 U20099 ( .A1(_05035_), .A2(_03272__PTR3), .ZN(_03272__PTR5) );
  AND2_X1 U20100 ( .A1(buf2_PTR18), .A2(_03272__PTR1), .ZN(_03272__PTR2) );
  AND2_X1 U20101 ( .A1(buf2_PTR20), .A2(_03272__PTR3), .ZN(_03272__PTR4) );
  AND2_X1 U20102 ( .A1(buf2_PTR22), .A2(_03272__PTR5), .ZN(_03272__PTR6) );
  AND2_X1 U20103 ( .A1(P3_rEIP_PTR2), .A2(_03268__PTR0), .ZN(_03268__PTR1) );
  AND2_X1 U20104 ( .A1(_05012_), .A2(_03268__PTR1), .ZN(_03268__PTR3) );
  AND2_X1 U20105 ( .A1(_05026_), .A2(_03268__PTR3), .ZN(_03268__PTR7) );
  AND2_X1 U20106 ( .A1(_05032_), .A2(_03268__PTR7), .ZN(_03268__PTR15) );
  AND2_X1 U20107 ( .A1(_05033_), .A2(_03268__PTR15), .ZN(_03268__PTR23) );
  AND2_X1 U20108 ( .A1(_05027_), .A2(_03268__PTR7), .ZN(_03268__PTR11) );
  AND2_X1 U20109 ( .A1(_05029_), .A2(_03268__PTR15), .ZN(_03268__PTR19) );
  AND2_X1 U20110 ( .A1(_05031_), .A2(_03268__PTR23), .ZN(_03268__PTR27) );
  AND2_X1 U20111 ( .A1(_05013_), .A2(_03268__PTR3), .ZN(_03268__PTR5) );
  AND2_X1 U20112 ( .A1(_05015_), .A2(_03268__PTR7), .ZN(_03268__PTR9) );
  AND2_X1 U20113 ( .A1(_05017_), .A2(_03268__PTR11), .ZN(_03268__PTR13) );
  AND2_X1 U20114 ( .A1(_05019_), .A2(_03268__PTR15), .ZN(_03268__PTR17) );
  AND2_X1 U20115 ( .A1(_05021_), .A2(_03268__PTR19), .ZN(_03268__PTR21) );
  AND2_X1 U20116 ( .A1(_05023_), .A2(_03268__PTR23), .ZN(_03268__PTR25) );
  AND2_X1 U20117 ( .A1(P3_rEIP_PTR3), .A2(_03268__PTR1), .ZN(_03268__PTR2) );
  AND2_X1 U20118 ( .A1(P3_rEIP_PTR5), .A2(_03268__PTR3), .ZN(_03268__PTR4) );
  AND2_X1 U20119 ( .A1(P3_rEIP_PTR7), .A2(_03268__PTR5), .ZN(_03268__PTR6) );
  AND2_X1 U20120 ( .A1(P3_rEIP_PTR9), .A2(_03268__PTR7), .ZN(_03268__PTR8) );
  AND2_X1 U20121 ( .A1(P3_rEIP_PTR11), .A2(_03268__PTR9), .ZN(_03268__PTR10) );
  AND2_X1 U20122 ( .A1(P3_rEIP_PTR13), .A2(_03268__PTR11), .ZN(_03268__PTR12) );
  AND2_X1 U20123 ( .A1(P3_rEIP_PTR15), .A2(_03268__PTR13), .ZN(_03268__PTR14) );
  AND2_X1 U20124 ( .A1(P3_rEIP_PTR17), .A2(_03268__PTR15), .ZN(_03268__PTR16) );
  AND2_X1 U20125 ( .A1(P3_rEIP_PTR19), .A2(_03268__PTR17), .ZN(_03268__PTR18) );
  AND2_X1 U20126 ( .A1(P3_rEIP_PTR21), .A2(_03268__PTR19), .ZN(_03268__PTR20) );
  AND2_X1 U20127 ( .A1(P3_rEIP_PTR23), .A2(_03268__PTR21), .ZN(_03268__PTR22) );
  AND2_X1 U20128 ( .A1(P3_rEIP_PTR25), .A2(_03268__PTR23), .ZN(_03268__PTR24) );
  AND2_X1 U20129 ( .A1(P3_rEIP_PTR27), .A2(_03268__PTR25), .ZN(_03268__PTR26) );
  AND2_X1 U20130 ( .A1(P3_rEIP_PTR29), .A2(_03268__PTR27), .ZN(_03268__PTR28) );
  AND2_X1 U20131 ( .A1(P3_rEIP_PTR3), .A2(_03283__PTR0), .ZN(_03283__PTR1) );
  AND2_X1 U20132 ( .A1(_05038_), .A2(_03283__PTR1), .ZN(_03283__PTR3) );
  AND2_X1 U20133 ( .A1(_05051_), .A2(_03283__PTR3), .ZN(_03283__PTR7) );
  AND2_X1 U20134 ( .A1(_05057_), .A2(_03283__PTR7), .ZN(_03283__PTR15) );
  AND2_X1 U20135 ( .A1(P3_rEIP_PTR5), .A2(P3_rEIP_PTR4), .ZN(_05038_) );
  AND2_X1 U20136 ( .A1(P3_rEIP_PTR7), .A2(P3_rEIP_PTR6), .ZN(_05039_) );
  AND2_X1 U20137 ( .A1(P3_rEIP_PTR9), .A2(P3_rEIP_PTR8), .ZN(_05040_) );
  AND2_X1 U20138 ( .A1(P3_rEIP_PTR11), .A2(P3_rEIP_PTR10), .ZN(_05041_) );
  AND2_X1 U20139 ( .A1(P3_rEIP_PTR13), .A2(P3_rEIP_PTR12), .ZN(_05042_) );
  AND2_X1 U20140 ( .A1(P3_rEIP_PTR15), .A2(P3_rEIP_PTR14), .ZN(_05043_) );
  AND2_X1 U20141 ( .A1(P3_rEIP_PTR17), .A2(P3_rEIP_PTR16), .ZN(_05044_) );
  AND2_X1 U20142 ( .A1(P3_rEIP_PTR19), .A2(P3_rEIP_PTR18), .ZN(_05045_) );
  AND2_X1 U20143 ( .A1(P3_rEIP_PTR21), .A2(P3_rEIP_PTR20), .ZN(_05046_) );
  AND2_X1 U20144 ( .A1(P3_rEIP_PTR23), .A2(P3_rEIP_PTR22), .ZN(_05047_) );
  AND2_X1 U20145 ( .A1(P3_rEIP_PTR25), .A2(P3_rEIP_PTR24), .ZN(_05048_) );
  AND2_X1 U20146 ( .A1(P3_rEIP_PTR27), .A2(P3_rEIP_PTR26), .ZN(_05049_) );
  AND2_X1 U20147 ( .A1(P3_rEIP_PTR29), .A2(P3_rEIP_PTR28), .ZN(_05050_) );
  AND2_X1 U20148 ( .A1(_05040_), .A2(_05039_), .ZN(_05051_) );
  AND2_X1 U20149 ( .A1(_05042_), .A2(_05041_), .ZN(_05052_) );
  AND2_X1 U20150 ( .A1(_05044_), .A2(_05043_), .ZN(_05053_) );
  AND2_X1 U20151 ( .A1(_05046_), .A2(_05045_), .ZN(_05054_) );
  AND2_X1 U20152 ( .A1(_05048_), .A2(_05047_), .ZN(_05055_) );
  AND2_X1 U20153 ( .A1(_05050_), .A2(_05049_), .ZN(_05056_) );
  AND2_X1 U20154 ( .A1(_05053_), .A2(_05052_), .ZN(_05057_) );
  AND2_X1 U20155 ( .A1(_05055_), .A2(_05054_), .ZN(_05058_) );
  AND2_X1 U20156 ( .A1(_05058_), .A2(_03283__PTR15), .ZN(_03283__PTR23) );
  AND2_X1 U20157 ( .A1(_05052_), .A2(_03283__PTR7), .ZN(_03283__PTR11) );
  AND2_X1 U20158 ( .A1(_05054_), .A2(_03283__PTR15), .ZN(_03283__PTR19) );
  AND2_X1 U20159 ( .A1(_05056_), .A2(_03283__PTR23), .ZN(_03283__PTR27) );
  AND2_X1 U20160 ( .A1(_05039_), .A2(_03283__PTR3), .ZN(_03283__PTR5) );
  AND2_X1 U20161 ( .A1(_05041_), .A2(_03283__PTR7), .ZN(_03283__PTR9) );
  AND2_X1 U20162 ( .A1(_05043_), .A2(_03283__PTR11), .ZN(_03283__PTR13) );
  AND2_X1 U20163 ( .A1(_05045_), .A2(_03283__PTR15), .ZN(_03283__PTR17) );
  AND2_X1 U20164 ( .A1(_05047_), .A2(_03283__PTR19), .ZN(_03283__PTR21) );
  AND2_X1 U20165 ( .A1(_05049_), .A2(_03283__PTR23), .ZN(_03283__PTR25) );
  AND2_X1 U20166 ( .A1(P3_rEIP_PTR4), .A2(_03283__PTR1), .ZN(_03283__PTR2) );
  AND2_X1 U20167 ( .A1(P3_rEIP_PTR6), .A2(_03283__PTR3), .ZN(_03283__PTR4) );
  AND2_X1 U20168 ( .A1(P3_rEIP_PTR8), .A2(_03283__PTR5), .ZN(_03283__PTR6) );
  AND2_X1 U20169 ( .A1(P3_rEIP_PTR10), .A2(_03283__PTR7), .ZN(_03283__PTR8) );
  AND2_X1 U20170 ( .A1(P3_rEIP_PTR12), .A2(_03283__PTR9), .ZN(_03283__PTR10) );
  AND2_X1 U20171 ( .A1(P3_rEIP_PTR14), .A2(_03283__PTR11), .ZN(_03283__PTR12) );
  AND2_X1 U20172 ( .A1(P3_rEIP_PTR16), .A2(_03283__PTR13), .ZN(_03283__PTR14) );
  AND2_X1 U20173 ( .A1(P3_rEIP_PTR18), .A2(_03283__PTR15), .ZN(_03283__PTR16) );
  AND2_X1 U20174 ( .A1(P3_rEIP_PTR20), .A2(_03283__PTR17), .ZN(_03283__PTR18) );
  AND2_X1 U20175 ( .A1(P3_rEIP_PTR22), .A2(_03283__PTR19), .ZN(_03283__PTR20) );
  AND2_X1 U20176 ( .A1(P3_rEIP_PTR24), .A2(_03283__PTR21), .ZN(_03283__PTR22) );
  AND2_X1 U20177 ( .A1(P3_rEIP_PTR26), .A2(_03283__PTR23), .ZN(_03283__PTR24) );
  AND2_X1 U20178 ( .A1(P3_rEIP_PTR28), .A2(_03283__PTR25), .ZN(_03283__PTR26) );
  AND2_X1 U20179 ( .A1(P3_rEIP_PTR30), .A2(_03283__PTR27), .ZN(_03283__PTR28) );
  AND2_X1 U20180 ( .A1(_05719_), .A2(_05753_), .ZN(_05756_) );
  AND2_X1 U20181 ( .A1(_05756_), .A2(P1_M_IO_n), .ZN(_05757_) );
  AND2_X1 U20182 ( .A1(_05757_), .A2(_05754_), .ZN(_05758_) );
  AND2_X1 U20183 ( .A1(_05758_), .A2(P1_W_R_n), .ZN(_05759_) );
  AND2_X1 U20184 ( .A1(_05759_), .A2(_05755_), .ZN(_05760_) );
  AND2_X1 U20185 ( .A1(_05714_), .A2(_05763_), .ZN(_05766_) );
  AND2_X1 U20186 ( .A1(_05766_), .A2(P2_M_IO_n), .ZN(_05767_) );
  AND2_X1 U20187 ( .A1(_05767_), .A2(_05764_), .ZN(_05768_) );
  AND2_X1 U20188 ( .A1(_05768_), .A2(P2_W_R_n), .ZN(_05769_) );
  AND2_X1 U20189 ( .A1(_05769_), .A2(_05765_), .ZN(_05770_) );
  AND2_X1 U20190 ( .A1(_05716_), .A2(_05763_), .ZN(_05737_) );
  AND2_X1 U20191 ( .A1(_05737_), .A2(P2_M_IO_n), .ZN(_05738_) );
  AND2_X1 U20192 ( .A1(_05738_), .A2(_05764_), .ZN(_05739_) );
  AND2_X1 U20193 ( .A1(_05739_), .A2(P2_W_R_n), .ZN(_05740_) );
  AND2_X1 U20194 ( .A1(_05740_), .A2(_05765_), .ZN(_05741_) );
  AND2_X1 U20195 ( .A1(_05742_), .A2(P3_M_IO_n), .ZN(_05746_) );
  AND2_X1 U20196 ( .A1(_05746_), .A2(_05743_), .ZN(_05747_) );
  AND2_X1 U20197 ( .A1(_05747_), .A2(_05744_), .ZN(_05748_) );
  AND2_X1 U20198 ( .A1(_05748_), .A2(_05745_), .ZN(_05749_) );
  AND2_X1 U20199 ( .A1(_05723_), .A2(_05727_), .ZN(_05761_) );
  AND2_X1 U20200 ( .A1(_05761_), .A2(_05731_), .ZN(_05762_) );
  AND2_X1 U20201 ( .A1(ready11), .A2(ready1), .ZN(P1_READY_n) );
  AND2_X1 U20202 ( .A1(ready12), .A2(ready21), .ZN(P2_READY_n) );
  AND2_X1 U20203 ( .A1(ready22), .A2(ready2), .ZN(P3_READY_n) );
  OR2_X1 U20204 ( .A1(_02063_), .A2(_01852__PTR5), .ZN(_02064_) );
  OR2_X1 U20205 ( .A1(_02062_), .A2(_01851__PTR5), .ZN(_02063_) );
  OR2_X1 U20206 ( .A1(_02736__PTR4), .A2(_02061_), .ZN(_02062_) );
  OR2_X1 U20207 ( .A1(_02023_), .A2(_02024_), .ZN(_02025_) );
  AND2_X1 U20208 ( .A1(_02022_), .A2(P1_EAX_PTR31), .ZN(_02823_) );
  AND2_X1 U20209 ( .A1(_01979_), .A2(P1_Datai_PTR31), .ZN(_02786_) );
  AND2_X1 U20210 ( .A1(_01615_), .A2(P1_Datai_PTR31), .ZN(_02781_) );
  AND2_X1 U20211 ( .A1(_02000_), .A2(_01876__PTR4), .ZN(_01943_) );
  AND2_X1 U20212 ( .A1(_01894__PTR14), .A2(hold), .ZN(_01942_) );
  AND2_X1 U20213 ( .A1(_01940_), .A2(_01999_), .ZN(_01941_) );
  AND2_X1 U20214 ( .A1(P1_READY_n), .A2(P1_RequestPending), .ZN(_01940_) );
  AND2_X1 U20215 ( .A1(P1_rEIP_PTR0), .A2(P1_rEIP_PTR31), .ZN(_02777_) );
  AND2_X1 U20216 ( .A1(_02003_), .A2(_02059_), .ZN(_02060_) );
  OR2_X1 U20217 ( .A1(hold), .A2(_01876__PTR4), .ZN(_02059_) );
  AND2_X1 U20218 ( .A1(_02048_), .A2(P1_RequestPending), .ZN(_02049_) );
  AND2_X1 U20219 ( .A1(hold), .A2(P1_READY_n), .ZN(_02021_) );
  AND2_X1 U20220 ( .A1(_02011_), .A2(_01894__PTR14), .ZN(_02012_) );
  AND2_X1 U20221 ( .A1(_01876__PTR4), .A2(_01999_), .ZN(_02011_) );
  AND2_X1 U20222 ( .A1(_02007_), .A2(_02003_), .ZN(_02008_) );
  AND2_X1 U20223 ( .A1(_01876__PTR21), .A2(P1_READY_n), .ZN(_02007_) );
  AND2_X1 U20224 ( .A1(P1_RequestPending), .A2(_01999_), .ZN(_01876__PTR21) );
  AND2_X1 U20225 ( .A1(_02004_), .A2(_02003_), .ZN(_02005_) );
  AND2_X1 U20226 ( .A1(_02002_), .A2(P1_READY_n), .ZN(_02004_) );
  OR2_X1 U20227 ( .A1(P1_RequestPending), .A2(hold), .ZN(_02002_) );
  AND2_X1 U20228 ( .A1(P1_READY_n), .A2(na), .ZN(_02001_) );
  AND2_X1 U20229 ( .A1(_02000_), .A2(P1_RequestPending), .ZN(_01769__PTR4) );
  AND2_X1 U20230 ( .A1(_01894__PTR14), .A2(_01999_), .ZN(_02000_) );
  AND2_X1 U20231 ( .A1(_01997_), .A2(P1_rEIP_PTR31), .ZN(_02792_) );
  OR2_X1 U20232 ( .A1(_02352_), .A2(_02145__PTR5), .ZN(_02353_) );
  OR2_X1 U20233 ( .A1(_02351_), .A2(_02144__PTR5), .ZN(_02352_) );
  OR2_X1 U20234 ( .A1(_02981__PTR4), .A2(_02350_), .ZN(_02351_) );
  OR2_X1 U20235 ( .A1(_02313_), .A2(_02314_), .ZN(_02315_) );
  AND2_X1 U20236 ( .A1(_02312_), .A2(P2_EAX_PTR31), .ZN(_03068_) );
  AND2_X1 U20237 ( .A1(_02271_), .A2(P2_Datai_PTR31), .ZN(_03031_) );
  AND2_X1 U20238 ( .A1(_01670_), .A2(P2_Datai_PTR31), .ZN(_03026_) );
  AND2_X1 U20239 ( .A1(_02291_), .A2(_02169__PTR4), .ZN(_02235_) );
  AND2_X1 U20240 ( .A1(_02186__PTR14), .A2(hold), .ZN(_02234_) );
  AND2_X1 U20241 ( .A1(_02232_), .A2(_01999_), .ZN(_02233_) );
  AND2_X1 U20242 ( .A1(P2_READY_n), .A2(P2_RequestPending), .ZN(_02232_) );
  AND2_X1 U20243 ( .A1(P2_rEIP_PTR0), .A2(P2_rEIP_PTR31), .ZN(_03022_) );
  AND2_X1 U20244 ( .A1(_02003_), .A2(_02348_), .ZN(_02349_) );
  OR2_X1 U20245 ( .A1(hold), .A2(_02169__PTR4), .ZN(_02348_) );
  AND2_X1 U20246 ( .A1(_02048_), .A2(P2_RequestPending), .ZN(_02338_) );
  AND2_X1 U20247 ( .A1(_02003_), .A2(_01999_), .ZN(_02048_) );
  AND2_X1 U20248 ( .A1(hold), .A2(P2_READY_n), .ZN(_02311_) );
  AND2_X1 U20249 ( .A1(_02301_), .A2(_02186__PTR14), .ZN(_02302_) );
  AND2_X1 U20250 ( .A1(_02169__PTR4), .A2(_01999_), .ZN(_02301_) );
  AND2_X1 U20251 ( .A1(_02297_), .A2(_02003_), .ZN(_02298_) );
  AND2_X1 U20252 ( .A1(_02169__PTR21), .A2(P2_READY_n), .ZN(_02297_) );
  AND2_X1 U20253 ( .A1(P2_RequestPending), .A2(_01999_), .ZN(_02169__PTR21) );
  AND2_X1 U20254 ( .A1(_02294_), .A2(_02003_), .ZN(_02295_) );
  AND2_X1 U20255 ( .A1(_02293_), .A2(P2_READY_n), .ZN(_02294_) );
  OR2_X1 U20256 ( .A1(P2_RequestPending), .A2(hold), .ZN(_02293_) );
  AND2_X1 U20257 ( .A1(P2_READY_n), .A2(na), .ZN(_02292_) );
  AND2_X1 U20258 ( .A1(_02291_), .A2(P2_RequestPending), .ZN(_01767__PTR4) );
  AND2_X1 U20259 ( .A1(_02186__PTR14), .A2(_01999_), .ZN(_02291_) );
  AND2_X1 U20260 ( .A1(_02289_), .A2(P2_rEIP_PTR31), .ZN(_03037_) );
  OR2_X1 U20261 ( .A1(_02641_), .A2(_02434__PTR5), .ZN(_02642_) );
  OR2_X1 U20262 ( .A1(_02640_), .A2(_02433__PTR5), .ZN(_02641_) );
  OR2_X1 U20263 ( .A1(_03226__PTR4), .A2(_02639_), .ZN(_02640_) );
  OR2_X1 U20264 ( .A1(_02602_), .A2(_02603_), .ZN(_02604_) );
  AND2_X1 U20265 ( .A1(_02601_), .A2(P3_EAX_PTR31), .ZN(_03313_) );
  AND2_X1 U20266 ( .A1(_02560_), .A2(buf2_PTR31), .ZN(_03276_) );
  AND2_X1 U20267 ( .A1(_01723_), .A2(buf2_PTR31), .ZN(_03271_) );
  AND2_X1 U20268 ( .A1(_02580_), .A2(_02458__PTR4), .ZN(_02524_) );
  AND2_X1 U20269 ( .A1(_02475__PTR14), .A2(hold), .ZN(_02523_) );
  AND2_X1 U20270 ( .A1(_02521_), .A2(_01999_), .ZN(_02522_) );
  AND2_X1 U20271 ( .A1(P3_READY_n), .A2(P3_RequestPending), .ZN(_02521_) );
  AND2_X1 U20272 ( .A1(P3_rEIP_PTR0), .A2(P3_rEIP_PTR31), .ZN(_03267_) );
  AND2_X1 U20273 ( .A1(_02003_), .A2(_02637_), .ZN(_02638_) );
  OR2_X1 U20274 ( .A1(hold), .A2(_02458__PTR4), .ZN(_02637_) );
  AND2_X1 U20275 ( .A1(_02048_), .A2(P3_RequestPending), .ZN(_02627_) );
  AND2_X1 U20276 ( .A1(hold), .A2(P3_READY_n), .ZN(_02600_) );
  AND2_X1 U20277 ( .A1(_02590_), .A2(_02475__PTR14), .ZN(_02591_) );
  AND2_X1 U20278 ( .A1(_02458__PTR4), .A2(_01999_), .ZN(_02590_) );
  AND2_X1 U20279 ( .A1(_02586_), .A2(_02003_), .ZN(_02587_) );
  AND2_X1 U20280 ( .A1(_02458__PTR21), .A2(P3_READY_n), .ZN(_02586_) );
  AND2_X1 U20281 ( .A1(P3_RequestPending), .A2(_01999_), .ZN(_02458__PTR21) );
  AND2_X1 U20282 ( .A1(_02583_), .A2(_02003_), .ZN(_02584_) );
  AND2_X1 U20283 ( .A1(_02582_), .A2(P3_READY_n), .ZN(_02583_) );
  OR2_X1 U20284 ( .A1(P3_RequestPending), .A2(hold), .ZN(_02582_) );
  AND2_X1 U20285 ( .A1(P3_READY_n), .A2(na), .ZN(_02581_) );
  AND2_X1 U20286 ( .A1(_02580_), .A2(P3_RequestPending), .ZN(_01765__PTR4) );
  AND2_X1 U20287 ( .A1(_02475__PTR14), .A2(_01999_), .ZN(_02580_) );
  AND2_X1 U20288 ( .A1(_02578_), .A2(P3_rEIP_PTR31), .ZN(_03282_) );
  AND2_X1 U20289 ( .A1(_01882__PTR8), .A2(_02124__PTR3), .ZN(_02123__PTR12) );
  AND2_X1 U20290 ( .A1(_01882__PTR9), .A2(_02124__PTR3), .ZN(_02123__PTR13) );
  AND2_X1 U20291 ( .A1(_01882__PTR10), .A2(_02124__PTR3), .ZN(_02123__PTR14) );
  AND2_X1 U20292 ( .A1(_01882__PTR11), .A2(_02124__PTR3), .ZN(_02123__PTR15) );
  AND2_X1 U20293 ( .A1(_01882__PTR8), .A2(_02124__PTR2), .ZN(_02123__PTR8) );
  AND2_X1 U20294 ( .A1(P1_rEIP_PTR1), .A2(_02124__PTR2), .ZN(_02123__PTR9) );
  AND2_X1 U20295 ( .A1(_01882__PTR6), .A2(_02124__PTR2), .ZN(_02123__PTR10) );
  AND2_X1 U20296 ( .A1(_01882__PTR7), .A2(_02124__PTR2), .ZN(_02123__PTR11) );
  AND2_X1 U20297 ( .A1(_01882__PTR8), .A2(_02124__PTR1), .ZN(_02123__PTR4) );
  AND2_X1 U20298 ( .A1(P1_rEIP_PTR1), .A2(_02124__PTR1), .ZN(_02123__PTR5) );
  AND2_X1 U20299 ( .A1(_01882__PTR2), .A2(_02124__PTR1), .ZN(_02123__PTR6) );
  MUX2_X1 U20300 ( .A(_02706__PTR0), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR0) );
  MUX2_X1 U20301 ( .A(_02706__PTR1), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR1) );
  MUX2_X1 U20302 ( .A(_02706__PTR2), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR2) );
  MUX2_X1 U20303 ( .A(_02706__PTR3), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR3) );
  MUX2_X1 U20304 ( .A(_02706__PTR4), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR4) );
  MUX2_X1 U20305 ( .A(_02706__PTR5), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR5) );
  MUX2_X1 U20306 ( .A(_02706__PTR6), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR6) );
  MUX2_X1 U20307 ( .A(_02706__PTR7), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR7) );
  MUX2_X1 U20308 ( .A(1'b0), .B(_02706__PTR0), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR8) );
  MUX2_X1 U20309 ( .A(1'b0), .B(_02706__PTR1), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR9) );
  MUX2_X1 U20310 ( .A(1'b0), .B(_02706__PTR2), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR10) );
  MUX2_X1 U20311 ( .A(1'b0), .B(_02706__PTR3), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR11) );
  MUX2_X1 U20312 ( .A(1'b0), .B(_02706__PTR4), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR12) );
  MUX2_X1 U20313 ( .A(1'b0), .B(_02706__PTR5), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR13) );
  MUX2_X1 U20314 ( .A(1'b0), .B(_02706__PTR6), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR14) );
  MUX2_X1 U20315 ( .A(1'b0), .B(_02706__PTR7), .S(P1_P1_InstQueueWr_Addr_PTR3), .Z(_01835__PTR15) );
  MUX2_X1 U20316 ( .A(_02705__PTR0), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR2), .Z(_02706__PTR0) );
  MUX2_X1 U20317 ( .A(_02705__PTR1), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR2), .Z(_02706__PTR1) );
  MUX2_X1 U20318 ( .A(_02705__PTR2), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR2), .Z(_02706__PTR2) );
  MUX2_X1 U20319 ( .A(_02705__PTR3), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR2), .Z(_02706__PTR3) );
  MUX2_X1 U20320 ( .A(1'b0), .B(_02705__PTR0), .S(P1_P1_InstQueueWr_Addr_PTR2), .Z(_02706__PTR4) );
  MUX2_X1 U20321 ( .A(1'b0), .B(_02705__PTR1), .S(P1_P1_InstQueueWr_Addr_PTR2), .Z(_02706__PTR5) );
  MUX2_X1 U20322 ( .A(1'b0), .B(_02705__PTR2), .S(P1_P1_InstQueueWr_Addr_PTR2), .Z(_02706__PTR6) );
  MUX2_X1 U20323 ( .A(1'b0), .B(_02705__PTR3), .S(P1_P1_InstQueueWr_Addr_PTR2), .Z(_02706__PTR7) );
  MUX2_X1 U20324 ( .A(_01836__PTR0), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR1), .Z(_02705__PTR0) );
  MUX2_X1 U20325 ( .A(P1_P1_InstQueueWr_Addr_PTR0), .B(1'b0), .S(P1_P1_InstQueueWr_Addr_PTR1), .Z(_02705__PTR1) );
  MUX2_X1 U20326 ( .A(1'b0), .B(_01836__PTR0), .S(P1_P1_InstQueueWr_Addr_PTR1), .Z(_02705__PTR2) );
  MUX2_X1 U20327 ( .A(1'b0), .B(P1_P1_InstQueueWr_Addr_PTR0), .S(P1_P1_InstQueueWr_Addr_PTR1), .Z(_02705__PTR3) );
  MUX2_X1 U20328 ( .A(_02708__PTR0), .B(1'b0), .S(_01836__PTR3), .Z(_01837__PTR0) );
  MUX2_X1 U20329 ( .A(_02708__PTR1), .B(1'b0), .S(_01836__PTR3), .Z(_01837__PTR1) );
  MUX2_X1 U20330 ( .A(_02708__PTR2), .B(1'b0), .S(_01836__PTR3), .Z(_01837__PTR2) );
  MUX2_X1 U20331 ( .A(_02708__PTR3), .B(1'b0), .S(_01836__PTR3), .Z(_01837__PTR3) );
  MUX2_X1 U20332 ( .A(_02708__PTR4), .B(1'b0), .S(_01836__PTR3), .Z(_01837__PTR4) );
  MUX2_X1 U20333 ( .A(_02708__PTR5), .B(1'b0), .S(_01836__PTR3), .Z(_01837__PTR5) );
  MUX2_X1 U20334 ( .A(_02708__PTR6), .B(1'b0), .S(_01836__PTR3), .Z(_01837__PTR6) );
  MUX2_X1 U20335 ( .A(_02708__PTR7), .B(1'b0), .S(_01836__PTR3), .Z(_01837__PTR7) );
  MUX2_X1 U20336 ( .A(1'b0), .B(_02708__PTR0), .S(_01836__PTR3), .Z(_01837__PTR8) );
  MUX2_X1 U20337 ( .A(1'b0), .B(_02708__PTR1), .S(_01836__PTR3), .Z(_01837__PTR9) );
  MUX2_X1 U20338 ( .A(1'b0), .B(_02708__PTR2), .S(_01836__PTR3), .Z(_01837__PTR10) );
  MUX2_X1 U20339 ( .A(1'b0), .B(_02708__PTR3), .S(_01836__PTR3), .Z(_01837__PTR11) );
  MUX2_X1 U20340 ( .A(1'b0), .B(_02708__PTR4), .S(_01836__PTR3), .Z(_01837__PTR12) );
  MUX2_X1 U20341 ( .A(1'b0), .B(_02708__PTR5), .S(_01836__PTR3), .Z(_01837__PTR13) );
  MUX2_X1 U20342 ( .A(1'b0), .B(_02708__PTR6), .S(_01836__PTR3), .Z(_01837__PTR14) );
  MUX2_X1 U20343 ( .A(1'b0), .B(_02708__PTR7), .S(_01836__PTR3), .Z(_01837__PTR15) );
  MUX2_X1 U20344 ( .A(_02707__PTR0), .B(1'b0), .S(_01836__PTR2), .Z(_02708__PTR0) );
  MUX2_X1 U20345 ( .A(_02707__PTR1), .B(1'b0), .S(_01836__PTR2), .Z(_02708__PTR1) );
  MUX2_X1 U20346 ( .A(_02707__PTR2), .B(1'b0), .S(_01836__PTR2), .Z(_02708__PTR2) );
  MUX2_X1 U20347 ( .A(_02707__PTR3), .B(1'b0), .S(_01836__PTR2), .Z(_02708__PTR3) );
  MUX2_X1 U20348 ( .A(1'b0), .B(_02707__PTR0), .S(_01836__PTR2), .Z(_02708__PTR4) );
  MUX2_X1 U20349 ( .A(1'b0), .B(_02707__PTR1), .S(_01836__PTR2), .Z(_02708__PTR5) );
  MUX2_X1 U20350 ( .A(1'b0), .B(_02707__PTR2), .S(_01836__PTR2), .Z(_02708__PTR6) );
  MUX2_X1 U20351 ( .A(1'b0), .B(_02707__PTR3), .S(_01836__PTR2), .Z(_02708__PTR7) );
  MUX2_X1 U20352 ( .A(P1_P1_InstQueueWr_Addr_PTR0), .B(1'b0), .S(_01836__PTR1), .Z(_02707__PTR0) );
  MUX2_X1 U20353 ( .A(_01836__PTR0), .B(1'b0), .S(_01836__PTR1), .Z(_02707__PTR1) );
  MUX2_X1 U20354 ( .A(1'b0), .B(P1_P1_InstQueueWr_Addr_PTR0), .S(_01836__PTR1), .Z(_02707__PTR2) );
  MUX2_X1 U20355 ( .A(1'b0), .B(_01836__PTR0), .S(_01836__PTR1), .Z(_02707__PTR3) );
  MUX2_X1 U20356 ( .A(_02710__PTR0), .B(1'b0), .S(_01838__PTR3), .Z(_01839__PTR0) );
  MUX2_X1 U20357 ( .A(_02710__PTR1), .B(1'b0), .S(_01838__PTR3), .Z(_01839__PTR1) );
  MUX2_X1 U20358 ( .A(_02710__PTR2), .B(1'b0), .S(_01838__PTR3), .Z(_01839__PTR2) );
  MUX2_X1 U20359 ( .A(_02710__PTR3), .B(1'b0), .S(_01838__PTR3), .Z(_01839__PTR3) );
  MUX2_X1 U20360 ( .A(_02710__PTR4), .B(1'b0), .S(_01838__PTR3), .Z(_01839__PTR4) );
  MUX2_X1 U20361 ( .A(_02710__PTR5), .B(1'b0), .S(_01838__PTR3), .Z(_01839__PTR5) );
  MUX2_X1 U20362 ( .A(_02710__PTR6), .B(1'b0), .S(_01838__PTR3), .Z(_01839__PTR6) );
  MUX2_X1 U20363 ( .A(_02710__PTR7), .B(1'b0), .S(_01838__PTR3), .Z(_01839__PTR7) );
  MUX2_X1 U20364 ( .A(1'b0), .B(_02710__PTR0), .S(_01838__PTR3), .Z(_01839__PTR8) );
  MUX2_X1 U20365 ( .A(1'b0), .B(_02710__PTR1), .S(_01838__PTR3), .Z(_01839__PTR9) );
  MUX2_X1 U20366 ( .A(1'b0), .B(_02710__PTR2), .S(_01838__PTR3), .Z(_01839__PTR10) );
  MUX2_X1 U20367 ( .A(1'b0), .B(_02710__PTR3), .S(_01838__PTR3), .Z(_01839__PTR11) );
  MUX2_X1 U20368 ( .A(1'b0), .B(_02710__PTR4), .S(_01838__PTR3), .Z(_01839__PTR12) );
  MUX2_X1 U20369 ( .A(1'b0), .B(_02710__PTR5), .S(_01838__PTR3), .Z(_01839__PTR13) );
  MUX2_X1 U20370 ( .A(1'b0), .B(_02710__PTR6), .S(_01838__PTR3), .Z(_01839__PTR14) );
  MUX2_X1 U20371 ( .A(1'b0), .B(_02710__PTR7), .S(_01838__PTR3), .Z(_01839__PTR15) );
  MUX2_X1 U20372 ( .A(_02709__PTR0), .B(1'b0), .S(_01838__PTR2), .Z(_02710__PTR0) );
  MUX2_X1 U20373 ( .A(_02709__PTR1), .B(1'b0), .S(_01838__PTR2), .Z(_02710__PTR1) );
  MUX2_X1 U20374 ( .A(_02709__PTR2), .B(1'b0), .S(_01838__PTR2), .Z(_02710__PTR2) );
  MUX2_X1 U20375 ( .A(_02709__PTR3), .B(1'b0), .S(_01838__PTR2), .Z(_02710__PTR3) );
  MUX2_X1 U20376 ( .A(1'b0), .B(_02709__PTR0), .S(_01838__PTR2), .Z(_02710__PTR4) );
  MUX2_X1 U20377 ( .A(1'b0), .B(_02709__PTR1), .S(_01838__PTR2), .Z(_02710__PTR5) );
  MUX2_X1 U20378 ( .A(1'b0), .B(_02709__PTR2), .S(_01838__PTR2), .Z(_02710__PTR6) );
  MUX2_X1 U20379 ( .A(1'b0), .B(_02709__PTR3), .S(_01838__PTR2), .Z(_02710__PTR7) );
  MUX2_X1 U20380 ( .A(_01836__PTR0), .B(1'b0), .S(_01838__PTR1), .Z(_02709__PTR0) );
  MUX2_X1 U20381 ( .A(P1_P1_InstQueueWr_Addr_PTR0), .B(1'b0), .S(_01838__PTR1), .Z(_02709__PTR1) );
  MUX2_X1 U20382 ( .A(1'b0), .B(_01836__PTR0), .S(_01838__PTR1), .Z(_02709__PTR2) );
  MUX2_X1 U20383 ( .A(1'b0), .B(P1_P1_InstQueueWr_Addr_PTR0), .S(_01838__PTR1), .Z(_02709__PTR3) );
  MUX2_X1 U20384 ( .A(_02712__PTR0), .B(1'b0), .S(_01840__PTR3), .Z(_01841__PTR0) );
  MUX2_X1 U20385 ( .A(_02712__PTR1), .B(1'b0), .S(_01840__PTR3), .Z(_01841__PTR1) );
  MUX2_X1 U20386 ( .A(_02712__PTR2), .B(1'b0), .S(_01840__PTR3), .Z(_01841__PTR2) );
  MUX2_X1 U20387 ( .A(_02712__PTR3), .B(1'b0), .S(_01840__PTR3), .Z(_01841__PTR3) );
  MUX2_X1 U20388 ( .A(_02712__PTR4), .B(1'b0), .S(_01840__PTR3), .Z(_01841__PTR4) );
  MUX2_X1 U20389 ( .A(_02712__PTR5), .B(1'b0), .S(_01840__PTR3), .Z(_01841__PTR5) );
  MUX2_X1 U20390 ( .A(_02712__PTR6), .B(1'b0), .S(_01840__PTR3), .Z(_01841__PTR6) );
  MUX2_X1 U20391 ( .A(_02712__PTR7), .B(1'b0), .S(_01840__PTR3), .Z(_01841__PTR7) );
  MUX2_X1 U20392 ( .A(1'b0), .B(_02712__PTR0), .S(_01840__PTR3), .Z(_01841__PTR8) );
  MUX2_X1 U20393 ( .A(1'b0), .B(_02712__PTR1), .S(_01840__PTR3), .Z(_01841__PTR9) );
  MUX2_X1 U20394 ( .A(1'b0), .B(_02712__PTR2), .S(_01840__PTR3), .Z(_01841__PTR10) );
  MUX2_X1 U20395 ( .A(1'b0), .B(_02712__PTR3), .S(_01840__PTR3), .Z(_01841__PTR11) );
  MUX2_X1 U20396 ( .A(1'b0), .B(_02712__PTR4), .S(_01840__PTR3), .Z(_01841__PTR12) );
  MUX2_X1 U20397 ( .A(1'b0), .B(_02712__PTR5), .S(_01840__PTR3), .Z(_01841__PTR13) );
  MUX2_X1 U20398 ( .A(1'b0), .B(_02712__PTR6), .S(_01840__PTR3), .Z(_01841__PTR14) );
  MUX2_X1 U20399 ( .A(1'b0), .B(_02712__PTR7), .S(_01840__PTR3), .Z(_01841__PTR15) );
  MUX2_X1 U20400 ( .A(_02711__PTR0), .B(1'b0), .S(_01840__PTR2), .Z(_02712__PTR0) );
  MUX2_X1 U20401 ( .A(_02711__PTR1), .B(1'b0), .S(_01840__PTR2), .Z(_02712__PTR1) );
  MUX2_X1 U20402 ( .A(_02711__PTR2), .B(1'b0), .S(_01840__PTR2), .Z(_02712__PTR2) );
  MUX2_X1 U20403 ( .A(_02711__PTR3), .B(1'b0), .S(_01840__PTR2), .Z(_02712__PTR3) );
  MUX2_X1 U20404 ( .A(1'b0), .B(_02711__PTR0), .S(_01840__PTR2), .Z(_02712__PTR4) );
  MUX2_X1 U20405 ( .A(1'b0), .B(_02711__PTR1), .S(_01840__PTR2), .Z(_02712__PTR5) );
  MUX2_X1 U20406 ( .A(1'b0), .B(_02711__PTR2), .S(_01840__PTR2), .Z(_02712__PTR6) );
  MUX2_X1 U20407 ( .A(1'b0), .B(_02711__PTR3), .S(_01840__PTR2), .Z(_02712__PTR7) );
  MUX2_X1 U20408 ( .A(P1_P1_InstQueueWr_Addr_PTR0), .B(1'b0), .S(_01840__PTR1), .Z(_02711__PTR0) );
  MUX2_X1 U20409 ( .A(_01836__PTR0), .B(1'b0), .S(_01840__PTR1), .Z(_02711__PTR1) );
  MUX2_X1 U20410 ( .A(1'b0), .B(P1_P1_InstQueueWr_Addr_PTR0), .S(_01840__PTR1), .Z(_02711__PTR2) );
  MUX2_X1 U20411 ( .A(1'b0), .B(_01836__PTR0), .S(_01840__PTR1), .Z(_02711__PTR3) );
  MUX2_X1 U20412 ( .A(_02755__PTR0), .B(_02755__PTR4), .S(P1_State_PTR2), .Z(_01843_) );
  MUX2_X1 U20413 ( .A(_02754__PTR0), .B(_02754__PTR6), .S(P1_State_PTR1), .Z(_02755__PTR0) );
  MUX2_X1 U20414 ( .A(1'b0), .B(_02754__PTR6), .S(P1_State_PTR1), .Z(_02755__PTR4) );
  MUX2_X1 U20415 ( .A(1'b1), .B(1'b0), .S(P1_State_PTR0), .Z(_02754__PTR0) );
  MUX2_X1 U20416 ( .A(_01842__PTR6), .B(P1_D_C_n), .S(P1_State_PTR0), .Z(_02754__PTR6) );
  MUX2_X1 U20417 ( .A(_02757__PTR0), .B(_02757__PTR4), .S(P1_State_PTR2), .Z(_01844_) );
  MUX2_X1 U20418 ( .A(_02756__PTR4), .B(P1_State_PTR0), .S(P1_State_PTR1), .Z(_02757__PTR0) );
  MUX2_X1 U20419 ( .A(_02756__PTR4), .B(_02756__PTR6), .S(P1_State_PTR1), .Z(_02757__PTR4) );
  MUX2_X1 U20420 ( .A(1'b1), .B(P1_ADS_n), .S(P1_State_PTR0), .Z(_02756__PTR4) );
  MUX2_X1 U20421 ( .A(1'b0), .B(1'b0), .S(P1_State_PTR0), .Z(_02756__PTR6) );
  MUX2_X1 U20422 ( .A(_02759__PTR0), .B(_02759__PTR4), .S(P1_State_PTR2), .Z(_01845_) );
  MUX2_X1 U20423 ( .A(_02754__PTR0), .B(_02758__PTR2), .S(P1_State_PTR1), .Z(_02759__PTR0) );
  MUX2_X1 U20424 ( .A(_02758__PTR4), .B(1'b0), .S(P1_State_PTR1), .Z(_02759__PTR4) );
  MUX2_X1 U20425 ( .A(1'b0), .B(bs16), .S(P1_State_PTR0), .Z(_02758__PTR2) );
  MUX2_X1 U20426 ( .A(bs16), .B(1'b0), .S(P1_State_PTR0), .Z(_02758__PTR4) );
  MUX2_X1 U20427 ( .A(_02761__PTR0), .B(_02761__PTR4), .S(P1_P1_State2_PTR2), .Z(_02762__PTR0) );
  MUX2_X1 U20428 ( .A(1'b1), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02761__PTR0) );
  MUX2_X1 U20429 ( .A(_02760__PTR4), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02761__PTR4) );
  MUX2_X1 U20430 ( .A(1'b0), .B(_01847__PTR5), .S(P1_P1_State2_PTR0), .Z(_02760__PTR4) );
  MUX2_X1 U20431 ( .A(_02761__PTR0), .B(_02764__PTR4), .S(P1_P1_State2_PTR2), .Z(_02765__PTR0) );
  MUX2_X1 U20432 ( .A(_02763__PTR4), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02764__PTR4) );
  MUX2_X1 U20433 ( .A(1'b0), .B(_01848__PTR5), .S(P1_P1_State2_PTR0), .Z(_02763__PTR4) );
  MUX2_X1 U20434 ( .A(_02767__PTR0), .B(_02767__PTR4), .S(P1_P1_State2_PTR2), .Z(_02768__PTR0) );
  MUX2_X1 U20435 ( .A(1'b1), .B(P1_P1_State2_PTR0), .S(P1_P1_State2_PTR1), .Z(_02767__PTR0) );
  MUX2_X1 U20436 ( .A(_02766__PTR4), .B(_02766__PTR6), .S(P1_P1_State2_PTR1), .Z(_02767__PTR4) );
  MUX2_X1 U20437 ( .A(1'b0), .B(_01849__PTR5), .S(P1_P1_State2_PTR0), .Z(_02766__PTR4) );
  MUX2_X1 U20438 ( .A(_01849__PTR6), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02766__PTR6) );
  MUX2_X1 U20439 ( .A(_02770__PTR0), .B(_02770__PTR4), .S(P1_P1_State2_PTR2), .Z(_02771__PTR0) );
  MUX2_X1 U20440 ( .A(_02769__PTR0), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02770__PTR0) );
  MUX2_X1 U20441 ( .A(_02769__PTR4), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02770__PTR4) );
  MUX2_X1 U20442 ( .A(1'b0), .B(1'b1), .S(P1_P1_State2_PTR0), .Z(_02769__PTR0) );
  MUX2_X1 U20443 ( .A(1'b0), .B(_01850__PTR5), .S(P1_P1_State2_PTR0), .Z(_02769__PTR4) );
  MUX2_X1 U20444 ( .A(_02832__PTR0), .B(_02832__PTR16), .S(P1_State_PTR2), .Z(_01877__PTR0) );
  MUX2_X1 U20445 ( .A(_02832__PTR1), .B(_02832__PTR17), .S(P1_State_PTR2), .Z(_01877__PTR1) );
  MUX2_X1 U20446 ( .A(_02832__PTR2), .B(_02832__PTR18), .S(P1_State_PTR2), .Z(_01877__PTR2) );
  MUX2_X1 U20447 ( .A(_02834__PTR0), .B(_02833__PTR0), .S(P1_State_PTR1), .Z(_02832__PTR0) );
  MUX2_X1 U20448 ( .A(_02834__PTR1), .B(_02833__PTR1), .S(P1_State_PTR1), .Z(_02832__PTR1) );
  MUX2_X1 U20449 ( .A(_02834__PTR2), .B(_02833__PTR2), .S(P1_State_PTR1), .Z(_02832__PTR2) );
  MUX2_X1 U20450 ( .A(_02833__PTR8), .B(_02833__PTR16), .S(P1_State_PTR1), .Z(_02832__PTR16) );
  MUX2_X1 U20451 ( .A(_02833__PTR9), .B(_02833__PTR17), .S(P1_State_PTR1), .Z(_02832__PTR17) );
  MUX2_X1 U20452 ( .A(_02833__PTR10), .B(_02833__PTR18), .S(P1_State_PTR1), .Z(_02832__PTR18) );
  MUX2_X1 U20453 ( .A(1'b1), .B(_01876__PTR4), .S(P1_State_PTR0), .Z(_02834__PTR0) );
  MUX2_X1 U20454 ( .A(1'b0), .B(P1_RequestPending), .S(P1_State_PTR0), .Z(_02834__PTR1) );
  MUX2_X1 U20455 ( .A(1'b0), .B(_01876__PTR6), .S(P1_State_PTR0), .Z(_02834__PTR2) );
  MUX2_X1 U20456 ( .A(1'b1), .B(_01876__PTR12), .S(P1_State_PTR0), .Z(_02833__PTR0) );
  MUX2_X1 U20457 ( .A(1'b1), .B(_01876__PTR13), .S(P1_State_PTR0), .Z(_02833__PTR1) );
  MUX2_X1 U20458 ( .A(1'b0), .B(_01876__PTR14), .S(P1_State_PTR0), .Z(_02833__PTR2) );
  MUX2_X1 U20459 ( .A(_01876__PTR16), .B(_01876__PTR20), .S(P1_State_PTR0), .Z(_02833__PTR8) );
  MUX2_X1 U20460 ( .A(_01876__PTR17), .B(_01876__PTR21), .S(P1_State_PTR0), .Z(_02833__PTR9) );
  MUX2_X1 U20461 ( .A(_01876__PTR18), .B(_01876__PTR22), .S(P1_State_PTR0), .Z(_02833__PTR10) );
  MUX2_X1 U20462 ( .A(1'b0), .B(_01876__PTR28), .S(P1_State_PTR0), .Z(_02833__PTR16) );
  MUX2_X1 U20463 ( .A(P1_READY_n), .B(_01876__PTR29), .S(P1_State_PTR0), .Z(_02833__PTR17) );
  MUX2_X1 U20464 ( .A(1'b1), .B(_01876__PTR30), .S(P1_State_PTR0), .Z(_02833__PTR18) );
  MUX2_X1 U20465 ( .A(_02836__PTR0), .B(_02836__PTR256), .S(P1_State_PTR2), .Z(_01879__PTR0) );
  MUX2_X1 U20466 ( .A(_02836__PTR2), .B(_02836__PTR258), .S(P1_State_PTR2), .Z(_01879__PTR2) );
  MUX2_X1 U20467 ( .A(_02836__PTR3), .B(_02836__PTR259), .S(P1_State_PTR2), .Z(_01879__PTR3) );
  MUX2_X1 U20468 ( .A(_02836__PTR4), .B(_02836__PTR260), .S(P1_State_PTR2), .Z(_01879__PTR4) );
  MUX2_X1 U20469 ( .A(_02836__PTR5), .B(_02836__PTR261), .S(P1_State_PTR2), .Z(_01879__PTR5) );
  MUX2_X1 U20470 ( .A(_02836__PTR6), .B(_02836__PTR262), .S(P1_State_PTR2), .Z(_01879__PTR6) );
  MUX2_X1 U20471 ( .A(_02836__PTR7), .B(_02836__PTR263), .S(P1_State_PTR2), .Z(_01879__PTR7) );
  MUX2_X1 U20472 ( .A(_02836__PTR8), .B(_02836__PTR264), .S(P1_State_PTR2), .Z(_01879__PTR8) );
  MUX2_X1 U20473 ( .A(_02836__PTR9), .B(_02836__PTR265), .S(P1_State_PTR2), .Z(_01879__PTR9) );
  MUX2_X1 U20474 ( .A(_02836__PTR10), .B(_02836__PTR266), .S(P1_State_PTR2), .Z(_01879__PTR10) );
  MUX2_X1 U20475 ( .A(_02836__PTR11), .B(_02836__PTR267), .S(P1_State_PTR2), .Z(_01879__PTR11) );
  MUX2_X1 U20476 ( .A(_02836__PTR12), .B(_02836__PTR268), .S(P1_State_PTR2), .Z(_01879__PTR12) );
  MUX2_X1 U20477 ( .A(_02836__PTR13), .B(_02836__PTR269), .S(P1_State_PTR2), .Z(_01879__PTR13) );
  MUX2_X1 U20478 ( .A(_02836__PTR14), .B(_02836__PTR270), .S(P1_State_PTR2), .Z(_01879__PTR14) );
  MUX2_X1 U20479 ( .A(_02836__PTR15), .B(_02836__PTR271), .S(P1_State_PTR2), .Z(_01879__PTR15) );
  MUX2_X1 U20480 ( .A(_02836__PTR16), .B(_02836__PTR272), .S(P1_State_PTR2), .Z(_01879__PTR16) );
  MUX2_X1 U20481 ( .A(_02836__PTR17), .B(_02836__PTR273), .S(P1_State_PTR2), .Z(_01879__PTR17) );
  MUX2_X1 U20482 ( .A(_02836__PTR18), .B(_02836__PTR274), .S(P1_State_PTR2), .Z(_01879__PTR18) );
  MUX2_X1 U20483 ( .A(_02836__PTR19), .B(_02836__PTR275), .S(P1_State_PTR2), .Z(_01879__PTR19) );
  MUX2_X1 U20484 ( .A(_02836__PTR20), .B(_02836__PTR276), .S(P1_State_PTR2), .Z(_01879__PTR20) );
  MUX2_X1 U20485 ( .A(_02836__PTR21), .B(_02836__PTR277), .S(P1_State_PTR2), .Z(_01879__PTR21) );
  MUX2_X1 U20486 ( .A(_02836__PTR22), .B(_02836__PTR278), .S(P1_State_PTR2), .Z(_01879__PTR22) );
  MUX2_X1 U20487 ( .A(_02836__PTR23), .B(_02836__PTR279), .S(P1_State_PTR2), .Z(_01879__PTR23) );
  MUX2_X1 U20488 ( .A(_02836__PTR24), .B(_02836__PTR280), .S(P1_State_PTR2), .Z(_01879__PTR24) );
  MUX2_X1 U20489 ( .A(_02836__PTR25), .B(_02836__PTR281), .S(P1_State_PTR2), .Z(_01879__PTR25) );
  MUX2_X1 U20490 ( .A(_02836__PTR26), .B(_02836__PTR282), .S(P1_State_PTR2), .Z(_01879__PTR26) );
  MUX2_X1 U20491 ( .A(_02836__PTR27), .B(_02836__PTR283), .S(P1_State_PTR2), .Z(_01879__PTR27) );
  MUX2_X1 U20492 ( .A(_02836__PTR28), .B(_02836__PTR284), .S(P1_State_PTR2), .Z(_01879__PTR28) );
  MUX2_X1 U20493 ( .A(_02836__PTR29), .B(_02836__PTR285), .S(P1_State_PTR2), .Z(_01879__PTR29) );
  MUX2_X1 U20494 ( .A(_02836__PTR30), .B(_02836__PTR286), .S(P1_State_PTR2), .Z(_01879__PTR30) );
  MUX2_X1 U20495 ( .A(_02836__PTR32), .B(_02836__PTR288), .S(P1_State_PTR2), .Z(_01879__PTR32) );
  MUX2_X1 U20496 ( .A(_02756__PTR6), .B(_02835__PTR128), .S(P1_State_PTR1), .Z(_02836__PTR0) );
  MUX2_X1 U20497 ( .A(_02835__PTR258), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR2) );
  MUX2_X1 U20498 ( .A(_02835__PTR259), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR3) );
  MUX2_X1 U20499 ( .A(_02835__PTR260), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR4) );
  MUX2_X1 U20500 ( .A(_02835__PTR261), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR5) );
  MUX2_X1 U20501 ( .A(_02835__PTR262), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR6) );
  MUX2_X1 U20502 ( .A(_02835__PTR263), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR7) );
  MUX2_X1 U20503 ( .A(_02835__PTR264), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR8) );
  MUX2_X1 U20504 ( .A(_02835__PTR265), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR9) );
  MUX2_X1 U20505 ( .A(_02835__PTR266), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR10) );
  MUX2_X1 U20506 ( .A(_02835__PTR267), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR11) );
  MUX2_X1 U20507 ( .A(_02835__PTR268), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR12) );
  MUX2_X1 U20508 ( .A(_02835__PTR269), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR13) );
  MUX2_X1 U20509 ( .A(_02835__PTR270), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR14) );
  MUX2_X1 U20510 ( .A(_02835__PTR271), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR15) );
  MUX2_X1 U20511 ( .A(_02835__PTR272), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR16) );
  MUX2_X1 U20512 ( .A(_02835__PTR273), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR17) );
  MUX2_X1 U20513 ( .A(_02835__PTR274), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR18) );
  MUX2_X1 U20514 ( .A(_02835__PTR275), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR19) );
  MUX2_X1 U20515 ( .A(_02835__PTR276), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR20) );
  MUX2_X1 U20516 ( .A(_02835__PTR277), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR21) );
  MUX2_X1 U20517 ( .A(_02835__PTR278), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR22) );
  MUX2_X1 U20518 ( .A(_02835__PTR279), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR23) );
  MUX2_X1 U20519 ( .A(_02835__PTR280), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR24) );
  MUX2_X1 U20520 ( .A(_02835__PTR281), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR25) );
  MUX2_X1 U20521 ( .A(_02835__PTR282), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR26) );
  MUX2_X1 U20522 ( .A(_02835__PTR283), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR27) );
  MUX2_X1 U20523 ( .A(_02835__PTR284), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR28) );
  MUX2_X1 U20524 ( .A(_02835__PTR285), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR29) );
  MUX2_X1 U20525 ( .A(_02835__PTR286), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR30) );
  MUX2_X1 U20526 ( .A(_02835__PTR288), .B(_02835__PTR160), .S(P1_State_PTR1), .Z(_02836__PTR32) );
  MUX2_X1 U20527 ( .A(_02835__PTR256), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR256) );
  MUX2_X1 U20528 ( .A(_02835__PTR258), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR258) );
  MUX2_X1 U20529 ( .A(_02835__PTR259), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR259) );
  MUX2_X1 U20530 ( .A(_02835__PTR260), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR260) );
  MUX2_X1 U20531 ( .A(_02835__PTR261), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR261) );
  MUX2_X1 U20532 ( .A(_02835__PTR262), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR262) );
  MUX2_X1 U20533 ( .A(_02835__PTR263), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR263) );
  MUX2_X1 U20534 ( .A(_02835__PTR264), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR264) );
  MUX2_X1 U20535 ( .A(_02835__PTR265), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR265) );
  MUX2_X1 U20536 ( .A(_02835__PTR266), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR266) );
  MUX2_X1 U20537 ( .A(_02835__PTR267), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR267) );
  MUX2_X1 U20538 ( .A(_02835__PTR268), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR268) );
  MUX2_X1 U20539 ( .A(_02835__PTR269), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR269) );
  MUX2_X1 U20540 ( .A(_02835__PTR270), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR270) );
  MUX2_X1 U20541 ( .A(_02835__PTR271), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR271) );
  MUX2_X1 U20542 ( .A(_02835__PTR272), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR272) );
  MUX2_X1 U20543 ( .A(_02835__PTR273), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR273) );
  MUX2_X1 U20544 ( .A(_02835__PTR274), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR274) );
  MUX2_X1 U20545 ( .A(_02835__PTR275), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR275) );
  MUX2_X1 U20546 ( .A(_02835__PTR276), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR276) );
  MUX2_X1 U20547 ( .A(_02835__PTR277), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR277) );
  MUX2_X1 U20548 ( .A(_02835__PTR278), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR278) );
  MUX2_X1 U20549 ( .A(_02835__PTR279), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR279) );
  MUX2_X1 U20550 ( .A(_02835__PTR280), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR280) );
  MUX2_X1 U20551 ( .A(_02835__PTR281), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR281) );
  MUX2_X1 U20552 ( .A(_02835__PTR282), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR282) );
  MUX2_X1 U20553 ( .A(_02835__PTR283), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR283) );
  MUX2_X1 U20554 ( .A(_02835__PTR284), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR284) );
  MUX2_X1 U20555 ( .A(_02835__PTR285), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR285) );
  MUX2_X1 U20556 ( .A(_02835__PTR286), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR286) );
  MUX2_X1 U20557 ( .A(_02835__PTR288), .B(1'b0), .S(P1_State_PTR1), .Z(_02836__PTR288) );
  MUX2_X1 U20558 ( .A(1'b0), .B(_01878__PTR256), .S(P1_State_PTR0), .Z(_02835__PTR128) );
  MUX2_X1 U20559 ( .A(1'b0), .B(1'b0), .S(P1_State_PTR0), .Z(_02835__PTR160) );
  MUX2_X1 U20560 ( .A(_01878__PTR256), .B(1'b0), .S(P1_State_PTR0), .Z(_02835__PTR256) );
  MUX2_X1 U20561 ( .A(1'b0), .B(P1_DataWidth_PTR2), .S(P1_State_PTR0), .Z(_02835__PTR258) );
  MUX2_X1 U20562 ( .A(1'b0), .B(P1_DataWidth_PTR3), .S(P1_State_PTR0), .Z(_02835__PTR259) );
  MUX2_X1 U20563 ( .A(1'b0), .B(P1_DataWidth_PTR4), .S(P1_State_PTR0), .Z(_02835__PTR260) );
  MUX2_X1 U20564 ( .A(1'b0), .B(P1_DataWidth_PTR5), .S(P1_State_PTR0), .Z(_02835__PTR261) );
  MUX2_X1 U20565 ( .A(1'b0), .B(P1_DataWidth_PTR6), .S(P1_State_PTR0), .Z(_02835__PTR262) );
  MUX2_X1 U20566 ( .A(1'b0), .B(P1_DataWidth_PTR7), .S(P1_State_PTR0), .Z(_02835__PTR263) );
  MUX2_X1 U20567 ( .A(1'b0), .B(P1_DataWidth_PTR8), .S(P1_State_PTR0), .Z(_02835__PTR264) );
  MUX2_X1 U20568 ( .A(1'b0), .B(P1_DataWidth_PTR9), .S(P1_State_PTR0), .Z(_02835__PTR265) );
  MUX2_X1 U20569 ( .A(1'b0), .B(P1_DataWidth_PTR10), .S(P1_State_PTR0), .Z(_02835__PTR266) );
  MUX2_X1 U20570 ( .A(1'b0), .B(P1_DataWidth_PTR11), .S(P1_State_PTR0), .Z(_02835__PTR267) );
  MUX2_X1 U20571 ( .A(1'b0), .B(P1_DataWidth_PTR12), .S(P1_State_PTR0), .Z(_02835__PTR268) );
  MUX2_X1 U20572 ( .A(1'b0), .B(P1_DataWidth_PTR13), .S(P1_State_PTR0), .Z(_02835__PTR269) );
  MUX2_X1 U20573 ( .A(1'b0), .B(P1_DataWidth_PTR14), .S(P1_State_PTR0), .Z(_02835__PTR270) );
  MUX2_X1 U20574 ( .A(1'b0), .B(P1_DataWidth_PTR15), .S(P1_State_PTR0), .Z(_02835__PTR271) );
  MUX2_X1 U20575 ( .A(1'b0), .B(P1_DataWidth_PTR16), .S(P1_State_PTR0), .Z(_02835__PTR272) );
  MUX2_X1 U20576 ( .A(1'b0), .B(P1_DataWidth_PTR17), .S(P1_State_PTR0), .Z(_02835__PTR273) );
  MUX2_X1 U20577 ( .A(1'b0), .B(P1_DataWidth_PTR18), .S(P1_State_PTR0), .Z(_02835__PTR274) );
  MUX2_X1 U20578 ( .A(1'b0), .B(P1_DataWidth_PTR19), .S(P1_State_PTR0), .Z(_02835__PTR275) );
  MUX2_X1 U20579 ( .A(1'b0), .B(P1_DataWidth_PTR20), .S(P1_State_PTR0), .Z(_02835__PTR276) );
  MUX2_X1 U20580 ( .A(1'b0), .B(P1_DataWidth_PTR21), .S(P1_State_PTR0), .Z(_02835__PTR277) );
  MUX2_X1 U20581 ( .A(1'b0), .B(P1_DataWidth_PTR22), .S(P1_State_PTR0), .Z(_02835__PTR278) );
  MUX2_X1 U20582 ( .A(1'b0), .B(P1_DataWidth_PTR23), .S(P1_State_PTR0), .Z(_02835__PTR279) );
  MUX2_X1 U20583 ( .A(1'b0), .B(P1_DataWidth_PTR24), .S(P1_State_PTR0), .Z(_02835__PTR280) );
  MUX2_X1 U20584 ( .A(1'b0), .B(P1_DataWidth_PTR25), .S(P1_State_PTR0), .Z(_02835__PTR281) );
  MUX2_X1 U20585 ( .A(1'b0), .B(P1_DataWidth_PTR26), .S(P1_State_PTR0), .Z(_02835__PTR282) );
  MUX2_X1 U20586 ( .A(1'b0), .B(P1_DataWidth_PTR27), .S(P1_State_PTR0), .Z(_02835__PTR283) );
  MUX2_X1 U20587 ( .A(1'b0), .B(P1_DataWidth_PTR28), .S(P1_State_PTR0), .Z(_02835__PTR284) );
  MUX2_X1 U20588 ( .A(1'b0), .B(P1_DataWidth_PTR29), .S(P1_State_PTR0), .Z(_02835__PTR285) );
  MUX2_X1 U20589 ( .A(1'b0), .B(P1_DataWidth_PTR30), .S(P1_State_PTR0), .Z(_02835__PTR286) );
  MUX2_X1 U20590 ( .A(1'b0), .B(P1_DataWidth_PTR31), .S(P1_State_PTR0), .Z(_02835__PTR288) );
  MUX2_X1 U20591 ( .A(_02838__PTR0), .B(_02838__PTR128), .S(P1_State_PTR2), .Z(_01881__PTR0) );
  MUX2_X1 U20592 ( .A(_02838__PTR1), .B(_02838__PTR129), .S(P1_State_PTR2), .Z(_01881__PTR1) );
  MUX2_X1 U20593 ( .A(_02838__PTR2), .B(_02838__PTR130), .S(P1_State_PTR2), .Z(_01881__PTR2) );
  MUX2_X1 U20594 ( .A(_02838__PTR3), .B(_02838__PTR131), .S(P1_State_PTR2), .Z(_01881__PTR3) );
  MUX2_X1 U20595 ( .A(_02838__PTR4), .B(_02838__PTR132), .S(P1_State_PTR2), .Z(_01881__PTR4) );
  MUX2_X1 U20596 ( .A(_02838__PTR5), .B(_02838__PTR133), .S(P1_State_PTR2), .Z(_01881__PTR5) );
  MUX2_X1 U20597 ( .A(_02838__PTR6), .B(_02838__PTR134), .S(P1_State_PTR2), .Z(_01881__PTR6) );
  MUX2_X1 U20598 ( .A(_02838__PTR7), .B(_02838__PTR135), .S(P1_State_PTR2), .Z(_01881__PTR7) );
  MUX2_X1 U20599 ( .A(_02838__PTR8), .B(_02838__PTR136), .S(P1_State_PTR2), .Z(_01881__PTR8) );
  MUX2_X1 U20600 ( .A(_02838__PTR9), .B(_02838__PTR137), .S(P1_State_PTR2), .Z(_01881__PTR9) );
  MUX2_X1 U20601 ( .A(_02838__PTR10), .B(_02838__PTR138), .S(P1_State_PTR2), .Z(_01881__PTR10) );
  MUX2_X1 U20602 ( .A(_02838__PTR11), .B(_02838__PTR139), .S(P1_State_PTR2), .Z(_01881__PTR11) );
  MUX2_X1 U20603 ( .A(_02838__PTR12), .B(_02838__PTR140), .S(P1_State_PTR2), .Z(_01881__PTR12) );
  MUX2_X1 U20604 ( .A(_02838__PTR13), .B(_02838__PTR141), .S(P1_State_PTR2), .Z(_01881__PTR13) );
  MUX2_X1 U20605 ( .A(_02838__PTR14), .B(_02838__PTR142), .S(P1_State_PTR2), .Z(_01881__PTR14) );
  MUX2_X1 U20606 ( .A(_02838__PTR15), .B(_02838__PTR143), .S(P1_State_PTR2), .Z(_01881__PTR15) );
  MUX2_X1 U20607 ( .A(_02838__PTR16), .B(_02838__PTR144), .S(P1_State_PTR2), .Z(_01881__PTR16) );
  MUX2_X1 U20608 ( .A(_02838__PTR17), .B(_02838__PTR145), .S(P1_State_PTR2), .Z(_01881__PTR17) );
  MUX2_X1 U20609 ( .A(_02838__PTR18), .B(_02838__PTR146), .S(P1_State_PTR2), .Z(_01881__PTR18) );
  MUX2_X1 U20610 ( .A(_02838__PTR19), .B(_02838__PTR147), .S(P1_State_PTR2), .Z(_01881__PTR19) );
  MUX2_X1 U20611 ( .A(_02838__PTR20), .B(_02838__PTR148), .S(P1_State_PTR2), .Z(_01881__PTR20) );
  MUX2_X1 U20612 ( .A(_02838__PTR21), .B(_02838__PTR149), .S(P1_State_PTR2), .Z(_01881__PTR21) );
  MUX2_X1 U20613 ( .A(_02838__PTR22), .B(_02838__PTR150), .S(P1_State_PTR2), .Z(_01881__PTR22) );
  MUX2_X1 U20614 ( .A(_02838__PTR23), .B(_02838__PTR151), .S(P1_State_PTR2), .Z(_01881__PTR23) );
  MUX2_X1 U20615 ( .A(_02838__PTR24), .B(_02838__PTR152), .S(P1_State_PTR2), .Z(_01881__PTR24) );
  MUX2_X1 U20616 ( .A(_02838__PTR25), .B(_02838__PTR153), .S(P1_State_PTR2), .Z(_01881__PTR25) );
  MUX2_X1 U20617 ( .A(_02838__PTR26), .B(_02838__PTR154), .S(P1_State_PTR2), .Z(_01881__PTR26) );
  MUX2_X1 U20618 ( .A(_02838__PTR27), .B(_02838__PTR155), .S(P1_State_PTR2), .Z(_01881__PTR27) );
  MUX2_X1 U20619 ( .A(_02838__PTR28), .B(_02838__PTR156), .S(P1_State_PTR2), .Z(_01881__PTR28) );
  MUX2_X1 U20620 ( .A(_02838__PTR29), .B(_02838__PTR157), .S(P1_State_PTR2), .Z(_01881__PTR29) );
  MUX2_X1 U20621 ( .A(1'b0), .B(_02837__PTR64), .S(P1_State_PTR1), .Z(_02838__PTR0) );
  MUX2_X1 U20622 ( .A(1'b0), .B(_02837__PTR65), .S(P1_State_PTR1), .Z(_02838__PTR1) );
  MUX2_X1 U20623 ( .A(1'b0), .B(_02837__PTR66), .S(P1_State_PTR1), .Z(_02838__PTR2) );
  MUX2_X1 U20624 ( .A(1'b0), .B(_02837__PTR67), .S(P1_State_PTR1), .Z(_02838__PTR3) );
  MUX2_X1 U20625 ( .A(1'b0), .B(_02837__PTR68), .S(P1_State_PTR1), .Z(_02838__PTR4) );
  MUX2_X1 U20626 ( .A(1'b0), .B(_02837__PTR69), .S(P1_State_PTR1), .Z(_02838__PTR5) );
  MUX2_X1 U20627 ( .A(1'b0), .B(_02837__PTR70), .S(P1_State_PTR1), .Z(_02838__PTR6) );
  MUX2_X1 U20628 ( .A(1'b0), .B(_02837__PTR71), .S(P1_State_PTR1), .Z(_02838__PTR7) );
  MUX2_X1 U20629 ( .A(1'b0), .B(_02837__PTR72), .S(P1_State_PTR1), .Z(_02838__PTR8) );
  MUX2_X1 U20630 ( .A(1'b0), .B(_02837__PTR73), .S(P1_State_PTR1), .Z(_02838__PTR9) );
  MUX2_X1 U20631 ( .A(1'b0), .B(_02837__PTR74), .S(P1_State_PTR1), .Z(_02838__PTR10) );
  MUX2_X1 U20632 ( .A(1'b0), .B(_02837__PTR75), .S(P1_State_PTR1), .Z(_02838__PTR11) );
  MUX2_X1 U20633 ( .A(1'b0), .B(_02837__PTR76), .S(P1_State_PTR1), .Z(_02838__PTR12) );
  MUX2_X1 U20634 ( .A(1'b0), .B(_02837__PTR77), .S(P1_State_PTR1), .Z(_02838__PTR13) );
  MUX2_X1 U20635 ( .A(1'b0), .B(_02837__PTR78), .S(P1_State_PTR1), .Z(_02838__PTR14) );
  MUX2_X1 U20636 ( .A(1'b0), .B(_02837__PTR79), .S(P1_State_PTR1), .Z(_02838__PTR15) );
  MUX2_X1 U20637 ( .A(1'b0), .B(_02837__PTR80), .S(P1_State_PTR1), .Z(_02838__PTR16) );
  MUX2_X1 U20638 ( .A(1'b0), .B(_02837__PTR81), .S(P1_State_PTR1), .Z(_02838__PTR17) );
  MUX2_X1 U20639 ( .A(1'b0), .B(_02837__PTR82), .S(P1_State_PTR1), .Z(_02838__PTR18) );
  MUX2_X1 U20640 ( .A(1'b0), .B(_02837__PTR83), .S(P1_State_PTR1), .Z(_02838__PTR19) );
  MUX2_X1 U20641 ( .A(1'b0), .B(_02837__PTR84), .S(P1_State_PTR1), .Z(_02838__PTR20) );
  MUX2_X1 U20642 ( .A(1'b0), .B(_02837__PTR85), .S(P1_State_PTR1), .Z(_02838__PTR21) );
  MUX2_X1 U20643 ( .A(1'b0), .B(_02837__PTR86), .S(P1_State_PTR1), .Z(_02838__PTR22) );
  MUX2_X1 U20644 ( .A(1'b0), .B(_02837__PTR87), .S(P1_State_PTR1), .Z(_02838__PTR23) );
  MUX2_X1 U20645 ( .A(1'b0), .B(_02837__PTR88), .S(P1_State_PTR1), .Z(_02838__PTR24) );
  MUX2_X1 U20646 ( .A(1'b0), .B(_02837__PTR89), .S(P1_State_PTR1), .Z(_02838__PTR25) );
  MUX2_X1 U20647 ( .A(1'b0), .B(_02837__PTR90), .S(P1_State_PTR1), .Z(_02838__PTR26) );
  MUX2_X1 U20648 ( .A(1'b0), .B(_02837__PTR91), .S(P1_State_PTR1), .Z(_02838__PTR27) );
  MUX2_X1 U20649 ( .A(1'b0), .B(_02837__PTR92), .S(P1_State_PTR1), .Z(_02838__PTR28) );
  MUX2_X1 U20650 ( .A(1'b0), .B(_02837__PTR93), .S(P1_State_PTR1), .Z(_02838__PTR29) );
  MUX2_X1 U20651 ( .A(1'b0), .B(_02837__PTR192), .S(P1_State_PTR1), .Z(_02838__PTR128) );
  MUX2_X1 U20652 ( .A(1'b0), .B(_02837__PTR193), .S(P1_State_PTR1), .Z(_02838__PTR129) );
  MUX2_X1 U20653 ( .A(1'b0), .B(_02837__PTR194), .S(P1_State_PTR1), .Z(_02838__PTR130) );
  MUX2_X1 U20654 ( .A(1'b0), .B(_02837__PTR195), .S(P1_State_PTR1), .Z(_02838__PTR131) );
  MUX2_X1 U20655 ( .A(1'b0), .B(_02837__PTR196), .S(P1_State_PTR1), .Z(_02838__PTR132) );
  MUX2_X1 U20656 ( .A(1'b0), .B(_02837__PTR197), .S(P1_State_PTR1), .Z(_02838__PTR133) );
  MUX2_X1 U20657 ( .A(1'b0), .B(_02837__PTR198), .S(P1_State_PTR1), .Z(_02838__PTR134) );
  MUX2_X1 U20658 ( .A(1'b0), .B(_02837__PTR199), .S(P1_State_PTR1), .Z(_02838__PTR135) );
  MUX2_X1 U20659 ( .A(1'b0), .B(_02837__PTR200), .S(P1_State_PTR1), .Z(_02838__PTR136) );
  MUX2_X1 U20660 ( .A(1'b0), .B(_02837__PTR201), .S(P1_State_PTR1), .Z(_02838__PTR137) );
  MUX2_X1 U20661 ( .A(1'b0), .B(_02837__PTR202), .S(P1_State_PTR1), .Z(_02838__PTR138) );
  MUX2_X1 U20662 ( .A(1'b0), .B(_02837__PTR203), .S(P1_State_PTR1), .Z(_02838__PTR139) );
  MUX2_X1 U20663 ( .A(1'b0), .B(_02837__PTR204), .S(P1_State_PTR1), .Z(_02838__PTR140) );
  MUX2_X1 U20664 ( .A(1'b0), .B(_02837__PTR205), .S(P1_State_PTR1), .Z(_02838__PTR141) );
  MUX2_X1 U20665 ( .A(1'b0), .B(_02837__PTR206), .S(P1_State_PTR1), .Z(_02838__PTR142) );
  MUX2_X1 U20666 ( .A(1'b0), .B(_02837__PTR207), .S(P1_State_PTR1), .Z(_02838__PTR143) );
  MUX2_X1 U20667 ( .A(1'b0), .B(_02837__PTR208), .S(P1_State_PTR1), .Z(_02838__PTR144) );
  MUX2_X1 U20668 ( .A(1'b0), .B(_02837__PTR209), .S(P1_State_PTR1), .Z(_02838__PTR145) );
  MUX2_X1 U20669 ( .A(1'b0), .B(_02837__PTR210), .S(P1_State_PTR1), .Z(_02838__PTR146) );
  MUX2_X1 U20670 ( .A(1'b0), .B(_02837__PTR211), .S(P1_State_PTR1), .Z(_02838__PTR147) );
  MUX2_X1 U20671 ( .A(1'b0), .B(_02837__PTR212), .S(P1_State_PTR1), .Z(_02838__PTR148) );
  MUX2_X1 U20672 ( .A(1'b0), .B(_02837__PTR213), .S(P1_State_PTR1), .Z(_02838__PTR149) );
  MUX2_X1 U20673 ( .A(1'b0), .B(_02837__PTR214), .S(P1_State_PTR1), .Z(_02838__PTR150) );
  MUX2_X1 U20674 ( .A(1'b0), .B(_02837__PTR215), .S(P1_State_PTR1), .Z(_02838__PTR151) );
  MUX2_X1 U20675 ( .A(1'b0), .B(_02837__PTR216), .S(P1_State_PTR1), .Z(_02838__PTR152) );
  MUX2_X1 U20676 ( .A(1'b0), .B(_02837__PTR217), .S(P1_State_PTR1), .Z(_02838__PTR153) );
  MUX2_X1 U20677 ( .A(1'b0), .B(_02837__PTR218), .S(P1_State_PTR1), .Z(_02838__PTR154) );
  MUX2_X1 U20678 ( .A(1'b0), .B(_02837__PTR219), .S(P1_State_PTR1), .Z(_02838__PTR155) );
  MUX2_X1 U20679 ( .A(1'b0), .B(_02837__PTR220), .S(P1_State_PTR1), .Z(_02838__PTR156) );
  MUX2_X1 U20680 ( .A(1'b0), .B(_02837__PTR221), .S(P1_State_PTR1), .Z(_02838__PTR157) );
  MUX2_X1 U20681 ( .A(_01880__PTR64), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR64) );
  MUX2_X1 U20682 ( .A(_01880__PTR65), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR65) );
  MUX2_X1 U20683 ( .A(_01880__PTR66), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR66) );
  MUX2_X1 U20684 ( .A(_01880__PTR67), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR67) );
  MUX2_X1 U20685 ( .A(_01880__PTR68), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR68) );
  MUX2_X1 U20686 ( .A(_01880__PTR69), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR69) );
  MUX2_X1 U20687 ( .A(_01880__PTR70), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR70) );
  MUX2_X1 U20688 ( .A(_01880__PTR71), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR71) );
  MUX2_X1 U20689 ( .A(_01880__PTR72), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR72) );
  MUX2_X1 U20690 ( .A(_01880__PTR73), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR73) );
  MUX2_X1 U20691 ( .A(_01880__PTR74), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR74) );
  MUX2_X1 U20692 ( .A(_01880__PTR75), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR75) );
  MUX2_X1 U20693 ( .A(_01880__PTR76), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR76) );
  MUX2_X1 U20694 ( .A(_01880__PTR77), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR77) );
  MUX2_X1 U20695 ( .A(_01880__PTR78), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR78) );
  MUX2_X1 U20696 ( .A(_01880__PTR79), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR79) );
  MUX2_X1 U20697 ( .A(_01880__PTR80), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR80) );
  MUX2_X1 U20698 ( .A(_01880__PTR81), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR81) );
  MUX2_X1 U20699 ( .A(_01880__PTR82), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR82) );
  MUX2_X1 U20700 ( .A(_01880__PTR83), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR83) );
  MUX2_X1 U20701 ( .A(_01880__PTR84), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR84) );
  MUX2_X1 U20702 ( .A(_01880__PTR85), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR85) );
  MUX2_X1 U20703 ( .A(_01880__PTR86), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR86) );
  MUX2_X1 U20704 ( .A(_01880__PTR87), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR87) );
  MUX2_X1 U20705 ( .A(_01880__PTR88), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR88) );
  MUX2_X1 U20706 ( .A(_01880__PTR89), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR89) );
  MUX2_X1 U20707 ( .A(_01880__PTR90), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR90) );
  MUX2_X1 U20708 ( .A(_01880__PTR91), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR91) );
  MUX2_X1 U20709 ( .A(_01880__PTR92), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR92) );
  MUX2_X1 U20710 ( .A(_01880__PTR93), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR93) );
  MUX2_X1 U20711 ( .A(_01880__PTR192), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR192) );
  MUX2_X1 U20712 ( .A(_01880__PTR193), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR193) );
  MUX2_X1 U20713 ( .A(_01880__PTR194), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR194) );
  MUX2_X1 U20714 ( .A(_01880__PTR195), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR195) );
  MUX2_X1 U20715 ( .A(_01880__PTR196), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR196) );
  MUX2_X1 U20716 ( .A(_01880__PTR197), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR197) );
  MUX2_X1 U20717 ( .A(_01880__PTR198), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR198) );
  MUX2_X1 U20718 ( .A(_01880__PTR199), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR199) );
  MUX2_X1 U20719 ( .A(_01880__PTR200), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR200) );
  MUX2_X1 U20720 ( .A(_01880__PTR201), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR201) );
  MUX2_X1 U20721 ( .A(_01880__PTR202), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR202) );
  MUX2_X1 U20722 ( .A(_01880__PTR203), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR203) );
  MUX2_X1 U20723 ( .A(_01880__PTR204), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR204) );
  MUX2_X1 U20724 ( .A(_01880__PTR205), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR205) );
  MUX2_X1 U20725 ( .A(_01880__PTR206), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR206) );
  MUX2_X1 U20726 ( .A(_01880__PTR207), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR207) );
  MUX2_X1 U20727 ( .A(_01880__PTR208), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR208) );
  MUX2_X1 U20728 ( .A(_01880__PTR209), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR209) );
  MUX2_X1 U20729 ( .A(_01880__PTR210), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR210) );
  MUX2_X1 U20730 ( .A(_01880__PTR211), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR211) );
  MUX2_X1 U20731 ( .A(_01880__PTR212), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR212) );
  MUX2_X1 U20732 ( .A(_01880__PTR213), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR213) );
  MUX2_X1 U20733 ( .A(_01880__PTR214), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR214) );
  MUX2_X1 U20734 ( .A(_01880__PTR215), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR215) );
  MUX2_X1 U20735 ( .A(_01880__PTR216), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR216) );
  MUX2_X1 U20736 ( .A(_01880__PTR217), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR217) );
  MUX2_X1 U20737 ( .A(_01880__PTR218), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR218) );
  MUX2_X1 U20738 ( .A(_01880__PTR219), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR219) );
  MUX2_X1 U20739 ( .A(_01880__PTR220), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR220) );
  MUX2_X1 U20740 ( .A(_01880__PTR221), .B(1'b0), .S(P1_State_PTR0), .Z(_02837__PTR221) );
  INV_X1 U20741 ( .A(P1_rEIP_PTR0), .ZN(_02839__PTR43) );
  MUX2_X1 U20742 ( .A(1'b0), .B(P1_rEIP_PTR0), .S(P1_rEIP_PTR1), .Z(_01882__PTR2) );
  MUX2_X1 U20743 ( .A(_02839__PTR43), .B(P1_rEIP_PTR0), .S(P1_rEIP_PTR1), .Z(_01882__PTR6) );
  MUX2_X1 U20744 ( .A(P1_rEIP_PTR0), .B(1'b1), .S(P1_rEIP_PTR1), .Z(_01882__PTR8) );
  MUX2_X1 U20745 ( .A(_02839__PTR43), .B(1'b1), .S(P1_rEIP_PTR1), .Z(_01882__PTR9) );
  MUX2_X1 U20746 ( .A(1'b1), .B(P1_rEIP_PTR0), .S(P1_rEIP_PTR1), .Z(_01882__PTR10) );
  MUX2_X1 U20747 ( .A(1'b1), .B(_02839__PTR43), .S(P1_rEIP_PTR1), .Z(_01882__PTR11) );
  MUX2_X1 U20748 ( .A(_02842__PTR0), .B(_02842__PTR64), .S(P1_P1_InstQueueRd_Addr_PTR3), .Z(_01883__PTR0) );
  MUX2_X1 U20749 ( .A(_02842__PTR1), .B(_02842__PTR65), .S(P1_P1_InstQueueRd_Addr_PTR3), .Z(_01883__PTR1) );
  MUX2_X1 U20750 ( .A(_02842__PTR2), .B(_02842__PTR66), .S(P1_P1_InstQueueRd_Addr_PTR3), .Z(_01883__PTR2) );
  MUX2_X1 U20751 ( .A(_02842__PTR3), .B(_02842__PTR67), .S(P1_P1_InstQueueRd_Addr_PTR3), .Z(_01883__PTR3) );
  MUX2_X1 U20752 ( .A(_02842__PTR4), .B(_02842__PTR68), .S(P1_P1_InstQueueRd_Addr_PTR3), .Z(_01883__PTR4) );
  MUX2_X1 U20753 ( .A(_02842__PTR5), .B(_02842__PTR69), .S(P1_P1_InstQueueRd_Addr_PTR3), .Z(_01883__PTR5) );
  MUX2_X1 U20754 ( .A(_02842__PTR6), .B(_02842__PTR70), .S(P1_P1_InstQueueRd_Addr_PTR3), .Z(_01883__PTR6) );
  MUX2_X1 U20755 ( .A(_02842__PTR7), .B(_02842__PTR71), .S(P1_P1_InstQueueRd_Addr_PTR3), .Z(_01883__PTR7) );
  MUX2_X1 U20756 ( .A(_02841__PTR0), .B(_02841__PTR32), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR0) );
  MUX2_X1 U20757 ( .A(_02841__PTR1), .B(_02841__PTR33), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR1) );
  MUX2_X1 U20758 ( .A(_02841__PTR2), .B(_02841__PTR34), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR2) );
  MUX2_X1 U20759 ( .A(_02841__PTR3), .B(_02841__PTR35), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR3) );
  MUX2_X1 U20760 ( .A(_02841__PTR4), .B(_02841__PTR36), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR4) );
  MUX2_X1 U20761 ( .A(_02841__PTR5), .B(_02841__PTR37), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR5) );
  MUX2_X1 U20762 ( .A(_02841__PTR6), .B(_02841__PTR38), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR6) );
  MUX2_X1 U20763 ( .A(_02841__PTR7), .B(_02841__PTR39), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR7) );
  MUX2_X1 U20764 ( .A(_02841__PTR64), .B(_02841__PTR96), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR64) );
  MUX2_X1 U20765 ( .A(_02841__PTR65), .B(_02841__PTR97), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR65) );
  MUX2_X1 U20766 ( .A(_02841__PTR66), .B(_02841__PTR98), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR66) );
  MUX2_X1 U20767 ( .A(_02841__PTR67), .B(_02841__PTR99), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR67) );
  MUX2_X1 U20768 ( .A(_02841__PTR68), .B(_02841__PTR100), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR68) );
  MUX2_X1 U20769 ( .A(_02841__PTR69), .B(_02841__PTR101), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR69) );
  MUX2_X1 U20770 ( .A(_02841__PTR70), .B(_02841__PTR102), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR70) );
  MUX2_X1 U20771 ( .A(_02841__PTR71), .B(_02841__PTR103), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02842__PTR71) );
  MUX2_X1 U20772 ( .A(_02840__PTR0), .B(_02840__PTR16), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR0) );
  MUX2_X1 U20773 ( .A(_02840__PTR1), .B(_02840__PTR17), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR1) );
  MUX2_X1 U20774 ( .A(_02840__PTR2), .B(_02840__PTR18), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR2) );
  MUX2_X1 U20775 ( .A(_02840__PTR3), .B(_02840__PTR19), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR3) );
  MUX2_X1 U20776 ( .A(_02840__PTR4), .B(_02840__PTR20), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR4) );
  MUX2_X1 U20777 ( .A(_02840__PTR5), .B(_02840__PTR21), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR5) );
  MUX2_X1 U20778 ( .A(_02840__PTR6), .B(_02840__PTR22), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR6) );
  MUX2_X1 U20779 ( .A(_02840__PTR7), .B(_02840__PTR23), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR7) );
  MUX2_X1 U20780 ( .A(_02840__PTR32), .B(_02840__PTR48), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR32) );
  MUX2_X1 U20781 ( .A(_02840__PTR33), .B(_02840__PTR49), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR33) );
  MUX2_X1 U20782 ( .A(_02840__PTR34), .B(_02840__PTR50), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR34) );
  MUX2_X1 U20783 ( .A(_02840__PTR35), .B(_02840__PTR51), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR35) );
  MUX2_X1 U20784 ( .A(_02840__PTR36), .B(_02840__PTR52), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR36) );
  MUX2_X1 U20785 ( .A(_02840__PTR37), .B(_02840__PTR53), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR37) );
  MUX2_X1 U20786 ( .A(_02840__PTR38), .B(_02840__PTR54), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR38) );
  MUX2_X1 U20787 ( .A(_02840__PTR39), .B(_02840__PTR55), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR39) );
  MUX2_X1 U20788 ( .A(_02840__PTR64), .B(_02840__PTR80), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR64) );
  MUX2_X1 U20789 ( .A(_02840__PTR65), .B(_02840__PTR81), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR65) );
  MUX2_X1 U20790 ( .A(_02840__PTR66), .B(_02840__PTR82), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR66) );
  MUX2_X1 U20791 ( .A(_02840__PTR67), .B(_02840__PTR83), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR67) );
  MUX2_X1 U20792 ( .A(_02840__PTR68), .B(_02840__PTR84), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR68) );
  MUX2_X1 U20793 ( .A(_02840__PTR69), .B(_02840__PTR85), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR69) );
  MUX2_X1 U20794 ( .A(_02840__PTR70), .B(_02840__PTR86), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR70) );
  MUX2_X1 U20795 ( .A(_02840__PTR71), .B(_02840__PTR87), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR71) );
  MUX2_X1 U20796 ( .A(_02840__PTR96), .B(_02840__PTR112), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR96) );
  MUX2_X1 U20797 ( .A(_02840__PTR97), .B(_02840__PTR113), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR97) );
  MUX2_X1 U20798 ( .A(_02840__PTR98), .B(_02840__PTR114), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR98) );
  MUX2_X1 U20799 ( .A(_02840__PTR99), .B(_02840__PTR115), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR99) );
  MUX2_X1 U20800 ( .A(_02840__PTR100), .B(_02840__PTR116), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR100) );
  MUX2_X1 U20801 ( .A(_02840__PTR101), .B(_02840__PTR117), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR101) );
  MUX2_X1 U20802 ( .A(_02840__PTR102), .B(_02840__PTR118), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR102) );
  MUX2_X1 U20803 ( .A(_02840__PTR103), .B(_02840__PTR119), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02841__PTR103) );
  MUX2_X1 U20804 ( .A(P1_P1_InstQueue_PTR0_PTR0), .B(P1_P1_InstQueue_PTR1_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR0) );
  MUX2_X1 U20805 ( .A(P1_P1_InstQueue_PTR0_PTR1), .B(P1_P1_InstQueue_PTR1_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR1) );
  MUX2_X1 U20806 ( .A(P1_P1_InstQueue_PTR0_PTR2), .B(P1_P1_InstQueue_PTR1_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR2) );
  MUX2_X1 U20807 ( .A(P1_P1_InstQueue_PTR0_PTR3), .B(P1_P1_InstQueue_PTR1_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR3) );
  MUX2_X1 U20808 ( .A(P1_P1_InstQueue_PTR0_PTR4), .B(P1_P1_InstQueue_PTR1_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR4) );
  MUX2_X1 U20809 ( .A(P1_P1_InstQueue_PTR0_PTR5), .B(P1_P1_InstQueue_PTR1_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR5) );
  MUX2_X1 U20810 ( .A(P1_P1_InstQueue_PTR0_PTR6), .B(P1_P1_InstQueue_PTR1_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR6) );
  MUX2_X1 U20811 ( .A(P1_P1_InstQueue_PTR0_PTR7), .B(P1_P1_InstQueue_PTR1_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR7) );
  MUX2_X1 U20812 ( .A(P1_P1_InstQueue_PTR2_PTR0), .B(P1_P1_InstQueue_PTR3_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR16) );
  MUX2_X1 U20813 ( .A(P1_P1_InstQueue_PTR2_PTR1), .B(P1_P1_InstQueue_PTR3_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR17) );
  MUX2_X1 U20814 ( .A(P1_P1_InstQueue_PTR2_PTR2), .B(P1_P1_InstQueue_PTR3_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR18) );
  MUX2_X1 U20815 ( .A(P1_P1_InstQueue_PTR2_PTR3), .B(P1_P1_InstQueue_PTR3_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR19) );
  MUX2_X1 U20816 ( .A(P1_P1_InstQueue_PTR2_PTR4), .B(P1_P1_InstQueue_PTR3_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR20) );
  MUX2_X1 U20817 ( .A(P1_P1_InstQueue_PTR2_PTR5), .B(P1_P1_InstQueue_PTR3_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR21) );
  MUX2_X1 U20818 ( .A(P1_P1_InstQueue_PTR2_PTR6), .B(P1_P1_InstQueue_PTR3_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR22) );
  MUX2_X1 U20819 ( .A(P1_P1_InstQueue_PTR2_PTR7), .B(P1_P1_InstQueue_PTR3_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR23) );
  MUX2_X1 U20820 ( .A(P1_P1_InstQueue_PTR4_PTR0), .B(P1_P1_InstQueue_PTR5_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR32) );
  MUX2_X1 U20821 ( .A(P1_P1_InstQueue_PTR4_PTR1), .B(P1_P1_InstQueue_PTR5_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR33) );
  MUX2_X1 U20822 ( .A(P1_P1_InstQueue_PTR4_PTR2), .B(P1_P1_InstQueue_PTR5_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR34) );
  MUX2_X1 U20823 ( .A(P1_P1_InstQueue_PTR4_PTR3), .B(P1_P1_InstQueue_PTR5_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR35) );
  MUX2_X1 U20824 ( .A(P1_P1_InstQueue_PTR4_PTR4), .B(P1_P1_InstQueue_PTR5_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR36) );
  MUX2_X1 U20825 ( .A(P1_P1_InstQueue_PTR4_PTR5), .B(P1_P1_InstQueue_PTR5_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR37) );
  MUX2_X1 U20826 ( .A(P1_P1_InstQueue_PTR4_PTR6), .B(P1_P1_InstQueue_PTR5_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR38) );
  MUX2_X1 U20827 ( .A(P1_P1_InstQueue_PTR4_PTR7), .B(P1_P1_InstQueue_PTR5_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR39) );
  MUX2_X1 U20828 ( .A(P1_P1_InstQueue_PTR6_PTR0), .B(P1_P1_InstQueue_PTR7_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR48) );
  MUX2_X1 U20829 ( .A(P1_P1_InstQueue_PTR6_PTR1), .B(P1_P1_InstQueue_PTR7_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR49) );
  MUX2_X1 U20830 ( .A(P1_P1_InstQueue_PTR6_PTR2), .B(P1_P1_InstQueue_PTR7_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR50) );
  MUX2_X1 U20831 ( .A(P1_P1_InstQueue_PTR6_PTR3), .B(P1_P1_InstQueue_PTR7_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR51) );
  MUX2_X1 U20832 ( .A(P1_P1_InstQueue_PTR6_PTR4), .B(P1_P1_InstQueue_PTR7_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR52) );
  MUX2_X1 U20833 ( .A(P1_P1_InstQueue_PTR6_PTR5), .B(P1_P1_InstQueue_PTR7_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR53) );
  MUX2_X1 U20834 ( .A(P1_P1_InstQueue_PTR6_PTR6), .B(P1_P1_InstQueue_PTR7_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR54) );
  MUX2_X1 U20835 ( .A(P1_P1_InstQueue_PTR6_PTR7), .B(P1_P1_InstQueue_PTR7_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR55) );
  MUX2_X1 U20836 ( .A(P1_P1_InstQueue_PTR8_PTR0), .B(P1_P1_InstQueue_PTR9_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR64) );
  MUX2_X1 U20837 ( .A(P1_P1_InstQueue_PTR8_PTR1), .B(P1_P1_InstQueue_PTR9_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR65) );
  MUX2_X1 U20838 ( .A(P1_P1_InstQueue_PTR8_PTR2), .B(P1_P1_InstQueue_PTR9_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR66) );
  MUX2_X1 U20839 ( .A(P1_P1_InstQueue_PTR8_PTR3), .B(P1_P1_InstQueue_PTR9_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR67) );
  MUX2_X1 U20840 ( .A(P1_P1_InstQueue_PTR8_PTR4), .B(P1_P1_InstQueue_PTR9_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR68) );
  MUX2_X1 U20841 ( .A(P1_P1_InstQueue_PTR8_PTR5), .B(P1_P1_InstQueue_PTR9_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR69) );
  MUX2_X1 U20842 ( .A(P1_P1_InstQueue_PTR8_PTR6), .B(P1_P1_InstQueue_PTR9_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR70) );
  MUX2_X1 U20843 ( .A(P1_P1_InstQueue_PTR8_PTR7), .B(P1_P1_InstQueue_PTR9_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR71) );
  MUX2_X1 U20844 ( .A(P1_P1_InstQueue_PTR10_PTR0), .B(P1_P1_InstQueue_PTR11_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR80) );
  MUX2_X1 U20845 ( .A(P1_P1_InstQueue_PTR10_PTR1), .B(P1_P1_InstQueue_PTR11_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR81) );
  MUX2_X1 U20846 ( .A(P1_P1_InstQueue_PTR10_PTR2), .B(P1_P1_InstQueue_PTR11_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR82) );
  MUX2_X1 U20847 ( .A(P1_P1_InstQueue_PTR10_PTR3), .B(P1_P1_InstQueue_PTR11_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR83) );
  MUX2_X1 U20848 ( .A(P1_P1_InstQueue_PTR10_PTR4), .B(P1_P1_InstQueue_PTR11_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR84) );
  MUX2_X1 U20849 ( .A(P1_P1_InstQueue_PTR10_PTR5), .B(P1_P1_InstQueue_PTR11_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR85) );
  MUX2_X1 U20850 ( .A(P1_P1_InstQueue_PTR10_PTR6), .B(P1_P1_InstQueue_PTR11_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR86) );
  MUX2_X1 U20851 ( .A(P1_P1_InstQueue_PTR10_PTR7), .B(P1_P1_InstQueue_PTR11_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR87) );
  MUX2_X1 U20852 ( .A(P1_P1_InstQueue_PTR12_PTR0), .B(P1_P1_InstQueue_PTR13_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR96) );
  MUX2_X1 U20853 ( .A(P1_P1_InstQueue_PTR12_PTR1), .B(P1_P1_InstQueue_PTR13_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR97) );
  MUX2_X1 U20854 ( .A(P1_P1_InstQueue_PTR12_PTR2), .B(P1_P1_InstQueue_PTR13_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR98) );
  MUX2_X1 U20855 ( .A(P1_P1_InstQueue_PTR12_PTR3), .B(P1_P1_InstQueue_PTR13_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR99) );
  MUX2_X1 U20856 ( .A(P1_P1_InstQueue_PTR12_PTR4), .B(P1_P1_InstQueue_PTR13_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR100) );
  MUX2_X1 U20857 ( .A(P1_P1_InstQueue_PTR12_PTR5), .B(P1_P1_InstQueue_PTR13_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR101) );
  MUX2_X1 U20858 ( .A(P1_P1_InstQueue_PTR12_PTR6), .B(P1_P1_InstQueue_PTR13_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR102) );
  MUX2_X1 U20859 ( .A(P1_P1_InstQueue_PTR12_PTR7), .B(P1_P1_InstQueue_PTR13_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR103) );
  MUX2_X1 U20860 ( .A(P1_P1_InstQueue_PTR14_PTR0), .B(P1_P1_InstQueue_PTR15_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR112) );
  MUX2_X1 U20861 ( .A(P1_P1_InstQueue_PTR14_PTR1), .B(P1_P1_InstQueue_PTR15_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR113) );
  MUX2_X1 U20862 ( .A(P1_P1_InstQueue_PTR14_PTR2), .B(P1_P1_InstQueue_PTR15_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR114) );
  MUX2_X1 U20863 ( .A(P1_P1_InstQueue_PTR14_PTR3), .B(P1_P1_InstQueue_PTR15_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR115) );
  MUX2_X1 U20864 ( .A(P1_P1_InstQueue_PTR14_PTR4), .B(P1_P1_InstQueue_PTR15_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR116) );
  MUX2_X1 U20865 ( .A(P1_P1_InstQueue_PTR14_PTR5), .B(P1_P1_InstQueue_PTR15_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR117) );
  MUX2_X1 U20866 ( .A(P1_P1_InstQueue_PTR14_PTR6), .B(P1_P1_InstQueue_PTR15_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR118) );
  MUX2_X1 U20867 ( .A(P1_P1_InstQueue_PTR14_PTR7), .B(P1_P1_InstQueue_PTR15_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02840__PTR119) );
  MUX2_X1 U20868 ( .A(_02845__PTR0), .B(_02845__PTR64), .S(_01884__PTR6), .Z(_01885__PTR0) );
  MUX2_X1 U20869 ( .A(_02845__PTR1), .B(_02845__PTR65), .S(_01884__PTR6), .Z(_01885__PTR1) );
  MUX2_X1 U20870 ( .A(_02845__PTR2), .B(_02845__PTR66), .S(_01884__PTR6), .Z(_01885__PTR2) );
  MUX2_X1 U20871 ( .A(_02845__PTR3), .B(_02845__PTR67), .S(_01884__PTR6), .Z(_01885__PTR3) );
  MUX2_X1 U20872 ( .A(_02845__PTR4), .B(_02845__PTR68), .S(_01884__PTR6), .Z(_01885__PTR4) );
  MUX2_X1 U20873 ( .A(_02845__PTR5), .B(_02845__PTR69), .S(_01884__PTR6), .Z(_01885__PTR5) );
  MUX2_X1 U20874 ( .A(_02845__PTR6), .B(_02845__PTR70), .S(_01884__PTR6), .Z(_01885__PTR6) );
  MUX2_X1 U20875 ( .A(_02845__PTR7), .B(_02845__PTR71), .S(_01884__PTR6), .Z(_01885__PTR7) );
  MUX2_X1 U20876 ( .A(_02844__PTR0), .B(_02844__PTR32), .S(_01884__PTR5), .Z(_02845__PTR0) );
  MUX2_X1 U20877 ( .A(_02844__PTR1), .B(_02844__PTR33), .S(_01884__PTR5), .Z(_02845__PTR1) );
  MUX2_X1 U20878 ( .A(_02844__PTR2), .B(_02844__PTR34), .S(_01884__PTR5), .Z(_02845__PTR2) );
  MUX2_X1 U20879 ( .A(_02844__PTR3), .B(_02844__PTR35), .S(_01884__PTR5), .Z(_02845__PTR3) );
  MUX2_X1 U20880 ( .A(_02844__PTR4), .B(_02844__PTR36), .S(_01884__PTR5), .Z(_02845__PTR4) );
  MUX2_X1 U20881 ( .A(_02844__PTR5), .B(_02844__PTR37), .S(_01884__PTR5), .Z(_02845__PTR5) );
  MUX2_X1 U20882 ( .A(_02844__PTR6), .B(_02844__PTR38), .S(_01884__PTR5), .Z(_02845__PTR6) );
  MUX2_X1 U20883 ( .A(_02844__PTR7), .B(_02844__PTR39), .S(_01884__PTR5), .Z(_02845__PTR7) );
  MUX2_X1 U20884 ( .A(_02844__PTR64), .B(_02844__PTR96), .S(_01884__PTR5), .Z(_02845__PTR64) );
  MUX2_X1 U20885 ( .A(_02844__PTR65), .B(_02844__PTR97), .S(_01884__PTR5), .Z(_02845__PTR65) );
  MUX2_X1 U20886 ( .A(_02844__PTR66), .B(_02844__PTR98), .S(_01884__PTR5), .Z(_02845__PTR66) );
  MUX2_X1 U20887 ( .A(_02844__PTR67), .B(_02844__PTR99), .S(_01884__PTR5), .Z(_02845__PTR67) );
  MUX2_X1 U20888 ( .A(_02844__PTR68), .B(_02844__PTR100), .S(_01884__PTR5), .Z(_02845__PTR68) );
  MUX2_X1 U20889 ( .A(_02844__PTR69), .B(_02844__PTR101), .S(_01884__PTR5), .Z(_02845__PTR69) );
  MUX2_X1 U20890 ( .A(_02844__PTR70), .B(_02844__PTR102), .S(_01884__PTR5), .Z(_02845__PTR70) );
  MUX2_X1 U20891 ( .A(_02844__PTR71), .B(_02844__PTR103), .S(_01884__PTR5), .Z(_02845__PTR71) );
  MUX2_X1 U20892 ( .A(_02843__PTR0), .B(_02843__PTR16), .S(_01884__PTR4), .Z(_02844__PTR0) );
  MUX2_X1 U20893 ( .A(_02843__PTR1), .B(_02843__PTR17), .S(_01884__PTR4), .Z(_02844__PTR1) );
  MUX2_X1 U20894 ( .A(_02843__PTR2), .B(_02843__PTR18), .S(_01884__PTR4), .Z(_02844__PTR2) );
  MUX2_X1 U20895 ( .A(_02843__PTR3), .B(_02843__PTR19), .S(_01884__PTR4), .Z(_02844__PTR3) );
  MUX2_X1 U20896 ( .A(_02843__PTR4), .B(_02843__PTR20), .S(_01884__PTR4), .Z(_02844__PTR4) );
  MUX2_X1 U20897 ( .A(_02843__PTR5), .B(_02843__PTR21), .S(_01884__PTR4), .Z(_02844__PTR5) );
  MUX2_X1 U20898 ( .A(_02843__PTR6), .B(_02843__PTR22), .S(_01884__PTR4), .Z(_02844__PTR6) );
  MUX2_X1 U20899 ( .A(_02843__PTR7), .B(_02843__PTR23), .S(_01884__PTR4), .Z(_02844__PTR7) );
  MUX2_X1 U20900 ( .A(_02843__PTR32), .B(_02843__PTR48), .S(_01884__PTR4), .Z(_02844__PTR32) );
  MUX2_X1 U20901 ( .A(_02843__PTR33), .B(_02843__PTR49), .S(_01884__PTR4), .Z(_02844__PTR33) );
  MUX2_X1 U20902 ( .A(_02843__PTR34), .B(_02843__PTR50), .S(_01884__PTR4), .Z(_02844__PTR34) );
  MUX2_X1 U20903 ( .A(_02843__PTR35), .B(_02843__PTR51), .S(_01884__PTR4), .Z(_02844__PTR35) );
  MUX2_X1 U20904 ( .A(_02843__PTR36), .B(_02843__PTR52), .S(_01884__PTR4), .Z(_02844__PTR36) );
  MUX2_X1 U20905 ( .A(_02843__PTR37), .B(_02843__PTR53), .S(_01884__PTR4), .Z(_02844__PTR37) );
  MUX2_X1 U20906 ( .A(_02843__PTR38), .B(_02843__PTR54), .S(_01884__PTR4), .Z(_02844__PTR38) );
  MUX2_X1 U20907 ( .A(_02843__PTR39), .B(_02843__PTR55), .S(_01884__PTR4), .Z(_02844__PTR39) );
  MUX2_X1 U20908 ( .A(_02843__PTR64), .B(_02843__PTR80), .S(_01884__PTR4), .Z(_02844__PTR64) );
  MUX2_X1 U20909 ( .A(_02843__PTR65), .B(_02843__PTR81), .S(_01884__PTR4), .Z(_02844__PTR65) );
  MUX2_X1 U20910 ( .A(_02843__PTR66), .B(_02843__PTR82), .S(_01884__PTR4), .Z(_02844__PTR66) );
  MUX2_X1 U20911 ( .A(_02843__PTR67), .B(_02843__PTR83), .S(_01884__PTR4), .Z(_02844__PTR67) );
  MUX2_X1 U20912 ( .A(_02843__PTR68), .B(_02843__PTR84), .S(_01884__PTR4), .Z(_02844__PTR68) );
  MUX2_X1 U20913 ( .A(_02843__PTR69), .B(_02843__PTR85), .S(_01884__PTR4), .Z(_02844__PTR69) );
  MUX2_X1 U20914 ( .A(_02843__PTR70), .B(_02843__PTR86), .S(_01884__PTR4), .Z(_02844__PTR70) );
  MUX2_X1 U20915 ( .A(_02843__PTR71), .B(_02843__PTR87), .S(_01884__PTR4), .Z(_02844__PTR71) );
  MUX2_X1 U20916 ( .A(_02843__PTR96), .B(_02843__PTR112), .S(_01884__PTR4), .Z(_02844__PTR96) );
  MUX2_X1 U20917 ( .A(_02843__PTR97), .B(_02843__PTR113), .S(_01884__PTR4), .Z(_02844__PTR97) );
  MUX2_X1 U20918 ( .A(_02843__PTR98), .B(_02843__PTR114), .S(_01884__PTR4), .Z(_02844__PTR98) );
  MUX2_X1 U20919 ( .A(_02843__PTR99), .B(_02843__PTR115), .S(_01884__PTR4), .Z(_02844__PTR99) );
  MUX2_X1 U20920 ( .A(_02843__PTR100), .B(_02843__PTR116), .S(_01884__PTR4), .Z(_02844__PTR100) );
  MUX2_X1 U20921 ( .A(_02843__PTR101), .B(_02843__PTR117), .S(_01884__PTR4), .Z(_02844__PTR101) );
  MUX2_X1 U20922 ( .A(_02843__PTR102), .B(_02843__PTR118), .S(_01884__PTR4), .Z(_02844__PTR102) );
  MUX2_X1 U20923 ( .A(_02843__PTR103), .B(_02843__PTR119), .S(_01884__PTR4), .Z(_02844__PTR103) );
  MUX2_X1 U20924 ( .A(P1_P1_InstQueue_PTR1_PTR0), .B(P1_P1_InstQueue_PTR0_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR0) );
  MUX2_X1 U20925 ( .A(P1_P1_InstQueue_PTR1_PTR1), .B(P1_P1_InstQueue_PTR0_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR1) );
  MUX2_X1 U20926 ( .A(P1_P1_InstQueue_PTR1_PTR2), .B(P1_P1_InstQueue_PTR0_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR2) );
  MUX2_X1 U20927 ( .A(P1_P1_InstQueue_PTR1_PTR3), .B(P1_P1_InstQueue_PTR0_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR3) );
  MUX2_X1 U20928 ( .A(P1_P1_InstQueue_PTR1_PTR4), .B(P1_P1_InstQueue_PTR0_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR4) );
  MUX2_X1 U20929 ( .A(P1_P1_InstQueue_PTR1_PTR5), .B(P1_P1_InstQueue_PTR0_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR5) );
  MUX2_X1 U20930 ( .A(P1_P1_InstQueue_PTR1_PTR6), .B(P1_P1_InstQueue_PTR0_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR6) );
  MUX2_X1 U20931 ( .A(P1_P1_InstQueue_PTR1_PTR7), .B(P1_P1_InstQueue_PTR0_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR7) );
  MUX2_X1 U20932 ( .A(P1_P1_InstQueue_PTR3_PTR0), .B(P1_P1_InstQueue_PTR2_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR16) );
  MUX2_X1 U20933 ( .A(P1_P1_InstQueue_PTR3_PTR1), .B(P1_P1_InstQueue_PTR2_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR17) );
  MUX2_X1 U20934 ( .A(P1_P1_InstQueue_PTR3_PTR2), .B(P1_P1_InstQueue_PTR2_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR18) );
  MUX2_X1 U20935 ( .A(P1_P1_InstQueue_PTR3_PTR3), .B(P1_P1_InstQueue_PTR2_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR19) );
  MUX2_X1 U20936 ( .A(P1_P1_InstQueue_PTR3_PTR4), .B(P1_P1_InstQueue_PTR2_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR20) );
  MUX2_X1 U20937 ( .A(P1_P1_InstQueue_PTR3_PTR5), .B(P1_P1_InstQueue_PTR2_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR21) );
  MUX2_X1 U20938 ( .A(P1_P1_InstQueue_PTR3_PTR6), .B(P1_P1_InstQueue_PTR2_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR22) );
  MUX2_X1 U20939 ( .A(P1_P1_InstQueue_PTR3_PTR7), .B(P1_P1_InstQueue_PTR2_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR23) );
  MUX2_X1 U20940 ( .A(P1_P1_InstQueue_PTR5_PTR0), .B(P1_P1_InstQueue_PTR4_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR32) );
  MUX2_X1 U20941 ( .A(P1_P1_InstQueue_PTR5_PTR1), .B(P1_P1_InstQueue_PTR4_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR33) );
  MUX2_X1 U20942 ( .A(P1_P1_InstQueue_PTR5_PTR2), .B(P1_P1_InstQueue_PTR4_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR34) );
  MUX2_X1 U20943 ( .A(P1_P1_InstQueue_PTR5_PTR3), .B(P1_P1_InstQueue_PTR4_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR35) );
  MUX2_X1 U20944 ( .A(P1_P1_InstQueue_PTR5_PTR4), .B(P1_P1_InstQueue_PTR4_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR36) );
  MUX2_X1 U20945 ( .A(P1_P1_InstQueue_PTR5_PTR5), .B(P1_P1_InstQueue_PTR4_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR37) );
  MUX2_X1 U20946 ( .A(P1_P1_InstQueue_PTR5_PTR6), .B(P1_P1_InstQueue_PTR4_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR38) );
  MUX2_X1 U20947 ( .A(P1_P1_InstQueue_PTR5_PTR7), .B(P1_P1_InstQueue_PTR4_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR39) );
  MUX2_X1 U20948 ( .A(P1_P1_InstQueue_PTR7_PTR0), .B(P1_P1_InstQueue_PTR6_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR48) );
  MUX2_X1 U20949 ( .A(P1_P1_InstQueue_PTR7_PTR1), .B(P1_P1_InstQueue_PTR6_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR49) );
  MUX2_X1 U20950 ( .A(P1_P1_InstQueue_PTR7_PTR2), .B(P1_P1_InstQueue_PTR6_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR50) );
  MUX2_X1 U20951 ( .A(P1_P1_InstQueue_PTR7_PTR3), .B(P1_P1_InstQueue_PTR6_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR51) );
  MUX2_X1 U20952 ( .A(P1_P1_InstQueue_PTR7_PTR4), .B(P1_P1_InstQueue_PTR6_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR52) );
  MUX2_X1 U20953 ( .A(P1_P1_InstQueue_PTR7_PTR5), .B(P1_P1_InstQueue_PTR6_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR53) );
  MUX2_X1 U20954 ( .A(P1_P1_InstQueue_PTR7_PTR6), .B(P1_P1_InstQueue_PTR6_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR54) );
  MUX2_X1 U20955 ( .A(P1_P1_InstQueue_PTR7_PTR7), .B(P1_P1_InstQueue_PTR6_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR55) );
  MUX2_X1 U20956 ( .A(P1_P1_InstQueue_PTR9_PTR0), .B(P1_P1_InstQueue_PTR8_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR64) );
  MUX2_X1 U20957 ( .A(P1_P1_InstQueue_PTR9_PTR1), .B(P1_P1_InstQueue_PTR8_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR65) );
  MUX2_X1 U20958 ( .A(P1_P1_InstQueue_PTR9_PTR2), .B(P1_P1_InstQueue_PTR8_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR66) );
  MUX2_X1 U20959 ( .A(P1_P1_InstQueue_PTR9_PTR3), .B(P1_P1_InstQueue_PTR8_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR67) );
  MUX2_X1 U20960 ( .A(P1_P1_InstQueue_PTR9_PTR4), .B(P1_P1_InstQueue_PTR8_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR68) );
  MUX2_X1 U20961 ( .A(P1_P1_InstQueue_PTR9_PTR5), .B(P1_P1_InstQueue_PTR8_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR69) );
  MUX2_X1 U20962 ( .A(P1_P1_InstQueue_PTR9_PTR6), .B(P1_P1_InstQueue_PTR8_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR70) );
  MUX2_X1 U20963 ( .A(P1_P1_InstQueue_PTR9_PTR7), .B(P1_P1_InstQueue_PTR8_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR71) );
  MUX2_X1 U20964 ( .A(P1_P1_InstQueue_PTR11_PTR0), .B(P1_P1_InstQueue_PTR10_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR80) );
  MUX2_X1 U20965 ( .A(P1_P1_InstQueue_PTR11_PTR1), .B(P1_P1_InstQueue_PTR10_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR81) );
  MUX2_X1 U20966 ( .A(P1_P1_InstQueue_PTR11_PTR2), .B(P1_P1_InstQueue_PTR10_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR82) );
  MUX2_X1 U20967 ( .A(P1_P1_InstQueue_PTR11_PTR3), .B(P1_P1_InstQueue_PTR10_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR83) );
  MUX2_X1 U20968 ( .A(P1_P1_InstQueue_PTR11_PTR4), .B(P1_P1_InstQueue_PTR10_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR84) );
  MUX2_X1 U20969 ( .A(P1_P1_InstQueue_PTR11_PTR5), .B(P1_P1_InstQueue_PTR10_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR85) );
  MUX2_X1 U20970 ( .A(P1_P1_InstQueue_PTR11_PTR6), .B(P1_P1_InstQueue_PTR10_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR86) );
  MUX2_X1 U20971 ( .A(P1_P1_InstQueue_PTR11_PTR7), .B(P1_P1_InstQueue_PTR10_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR87) );
  MUX2_X1 U20972 ( .A(P1_P1_InstQueue_PTR13_PTR0), .B(P1_P1_InstQueue_PTR12_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR96) );
  MUX2_X1 U20973 ( .A(P1_P1_InstQueue_PTR13_PTR1), .B(P1_P1_InstQueue_PTR12_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR97) );
  MUX2_X1 U20974 ( .A(P1_P1_InstQueue_PTR13_PTR2), .B(P1_P1_InstQueue_PTR12_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR98) );
  MUX2_X1 U20975 ( .A(P1_P1_InstQueue_PTR13_PTR3), .B(P1_P1_InstQueue_PTR12_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR99) );
  MUX2_X1 U20976 ( .A(P1_P1_InstQueue_PTR13_PTR4), .B(P1_P1_InstQueue_PTR12_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR100) );
  MUX2_X1 U20977 ( .A(P1_P1_InstQueue_PTR13_PTR5), .B(P1_P1_InstQueue_PTR12_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR101) );
  MUX2_X1 U20978 ( .A(P1_P1_InstQueue_PTR13_PTR6), .B(P1_P1_InstQueue_PTR12_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR102) );
  MUX2_X1 U20979 ( .A(P1_P1_InstQueue_PTR13_PTR7), .B(P1_P1_InstQueue_PTR12_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR103) );
  MUX2_X1 U20980 ( .A(P1_P1_InstQueue_PTR15_PTR0), .B(P1_P1_InstQueue_PTR14_PTR0), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR112) );
  MUX2_X1 U20981 ( .A(P1_P1_InstQueue_PTR15_PTR1), .B(P1_P1_InstQueue_PTR14_PTR1), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR113) );
  MUX2_X1 U20982 ( .A(P1_P1_InstQueue_PTR15_PTR2), .B(P1_P1_InstQueue_PTR14_PTR2), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR114) );
  MUX2_X1 U20983 ( .A(P1_P1_InstQueue_PTR15_PTR3), .B(P1_P1_InstQueue_PTR14_PTR3), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR115) );
  MUX2_X1 U20984 ( .A(P1_P1_InstQueue_PTR15_PTR4), .B(P1_P1_InstQueue_PTR14_PTR4), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR116) );
  MUX2_X1 U20985 ( .A(P1_P1_InstQueue_PTR15_PTR5), .B(P1_P1_InstQueue_PTR14_PTR5), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR117) );
  MUX2_X1 U20986 ( .A(P1_P1_InstQueue_PTR15_PTR6), .B(P1_P1_InstQueue_PTR14_PTR6), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR118) );
  MUX2_X1 U20987 ( .A(P1_P1_InstQueue_PTR15_PTR7), .B(P1_P1_InstQueue_PTR14_PTR7), .S(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02843__PTR119) );
  MUX2_X1 U20988 ( .A(_02846__PTR0), .B(_02846__PTR64), .S(_01886__PTR6), .Z(_01887__PTR0) );
  MUX2_X1 U20989 ( .A(_02846__PTR1), .B(_02846__PTR65), .S(_01886__PTR6), .Z(_01887__PTR1) );
  MUX2_X1 U20990 ( .A(_02846__PTR2), .B(_02846__PTR66), .S(_01886__PTR6), .Z(_01887__PTR2) );
  MUX2_X1 U20991 ( .A(_02846__PTR3), .B(_02846__PTR67), .S(_01886__PTR6), .Z(_01887__PTR3) );
  MUX2_X1 U20992 ( .A(_02846__PTR4), .B(_02846__PTR68), .S(_01886__PTR6), .Z(_01887__PTR4) );
  MUX2_X1 U20993 ( .A(_02846__PTR5), .B(_02846__PTR69), .S(_01886__PTR6), .Z(_01887__PTR5) );
  MUX2_X1 U20994 ( .A(_02846__PTR6), .B(_02846__PTR70), .S(_01886__PTR6), .Z(_01887__PTR6) );
  MUX2_X1 U20995 ( .A(_02846__PTR7), .B(_02846__PTR71), .S(_01886__PTR6), .Z(_01887__PTR7) );
  MUX2_X1 U20996 ( .A(_02841__PTR32), .B(_02841__PTR0), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR0) );
  MUX2_X1 U20997 ( .A(_02841__PTR33), .B(_02841__PTR1), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR1) );
  MUX2_X1 U20998 ( .A(_02841__PTR34), .B(_02841__PTR2), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR2) );
  MUX2_X1 U20999 ( .A(_02841__PTR35), .B(_02841__PTR3), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR3) );
  MUX2_X1 U21000 ( .A(_02841__PTR36), .B(_02841__PTR4), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR4) );
  MUX2_X1 U21001 ( .A(_02841__PTR37), .B(_02841__PTR5), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR5) );
  MUX2_X1 U21002 ( .A(_02841__PTR38), .B(_02841__PTR6), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR6) );
  MUX2_X1 U21003 ( .A(_02841__PTR39), .B(_02841__PTR7), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR7) );
  MUX2_X1 U21004 ( .A(_02841__PTR96), .B(_02841__PTR64), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR64) );
  MUX2_X1 U21005 ( .A(_02841__PTR97), .B(_02841__PTR65), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR65) );
  MUX2_X1 U21006 ( .A(_02841__PTR98), .B(_02841__PTR66), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR66) );
  MUX2_X1 U21007 ( .A(_02841__PTR99), .B(_02841__PTR67), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR67) );
  MUX2_X1 U21008 ( .A(_02841__PTR100), .B(_02841__PTR68), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR68) );
  MUX2_X1 U21009 ( .A(_02841__PTR101), .B(_02841__PTR69), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR69) );
  MUX2_X1 U21010 ( .A(_02841__PTR102), .B(_02841__PTR70), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR70) );
  MUX2_X1 U21011 ( .A(_02841__PTR103), .B(_02841__PTR71), .S(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02846__PTR71) );
  MUX2_X1 U21012 ( .A(_02848__PTR0), .B(_02848__PTR64), .S(_01888__PTR6), .Z(_01889__PTR0) );
  MUX2_X1 U21013 ( .A(_02848__PTR1), .B(_02848__PTR65), .S(_01888__PTR6), .Z(_01889__PTR1) );
  MUX2_X1 U21014 ( .A(_02848__PTR2), .B(_02848__PTR66), .S(_01888__PTR6), .Z(_01889__PTR2) );
  MUX2_X1 U21015 ( .A(_02848__PTR3), .B(_02848__PTR67), .S(_01888__PTR6), .Z(_01889__PTR3) );
  MUX2_X1 U21016 ( .A(_02848__PTR4), .B(_02848__PTR68), .S(_01888__PTR6), .Z(_01889__PTR4) );
  MUX2_X1 U21017 ( .A(_02848__PTR5), .B(_02848__PTR69), .S(_01888__PTR6), .Z(_01889__PTR5) );
  MUX2_X1 U21018 ( .A(_02848__PTR6), .B(_02848__PTR70), .S(_01888__PTR6), .Z(_01889__PTR6) );
  MUX2_X1 U21019 ( .A(_02848__PTR7), .B(_02848__PTR71), .S(_01888__PTR6), .Z(_01889__PTR7) );
  MUX2_X1 U21020 ( .A(_02847__PTR0), .B(_02847__PTR32), .S(_01888__PTR5), .Z(_02848__PTR0) );
  MUX2_X1 U21021 ( .A(_02847__PTR1), .B(_02847__PTR33), .S(_01888__PTR5), .Z(_02848__PTR1) );
  MUX2_X1 U21022 ( .A(_02847__PTR2), .B(_02847__PTR34), .S(_01888__PTR5), .Z(_02848__PTR2) );
  MUX2_X1 U21023 ( .A(_02847__PTR3), .B(_02847__PTR35), .S(_01888__PTR5), .Z(_02848__PTR3) );
  MUX2_X1 U21024 ( .A(_02847__PTR4), .B(_02847__PTR36), .S(_01888__PTR5), .Z(_02848__PTR4) );
  MUX2_X1 U21025 ( .A(_02847__PTR5), .B(_02847__PTR37), .S(_01888__PTR5), .Z(_02848__PTR5) );
  MUX2_X1 U21026 ( .A(_02847__PTR6), .B(_02847__PTR38), .S(_01888__PTR5), .Z(_02848__PTR6) );
  MUX2_X1 U21027 ( .A(_02847__PTR7), .B(_02847__PTR39), .S(_01888__PTR5), .Z(_02848__PTR7) );
  MUX2_X1 U21028 ( .A(_02847__PTR64), .B(_02847__PTR96), .S(_01888__PTR5), .Z(_02848__PTR64) );
  MUX2_X1 U21029 ( .A(_02847__PTR65), .B(_02847__PTR97), .S(_01888__PTR5), .Z(_02848__PTR65) );
  MUX2_X1 U21030 ( .A(_02847__PTR66), .B(_02847__PTR98), .S(_01888__PTR5), .Z(_02848__PTR66) );
  MUX2_X1 U21031 ( .A(_02847__PTR67), .B(_02847__PTR99), .S(_01888__PTR5), .Z(_02848__PTR67) );
  MUX2_X1 U21032 ( .A(_02847__PTR68), .B(_02847__PTR100), .S(_01888__PTR5), .Z(_02848__PTR68) );
  MUX2_X1 U21033 ( .A(_02847__PTR69), .B(_02847__PTR101), .S(_01888__PTR5), .Z(_02848__PTR69) );
  MUX2_X1 U21034 ( .A(_02847__PTR70), .B(_02847__PTR102), .S(_01888__PTR5), .Z(_02848__PTR70) );
  MUX2_X1 U21035 ( .A(_02847__PTR71), .B(_02847__PTR103), .S(_01888__PTR5), .Z(_02848__PTR71) );
  MUX2_X1 U21036 ( .A(_02843__PTR0), .B(_02843__PTR16), .S(_01888__PTR4), .Z(_02847__PTR0) );
  MUX2_X1 U21037 ( .A(_02843__PTR1), .B(_02843__PTR17), .S(_01888__PTR4), .Z(_02847__PTR1) );
  MUX2_X1 U21038 ( .A(_02843__PTR2), .B(_02843__PTR18), .S(_01888__PTR4), .Z(_02847__PTR2) );
  MUX2_X1 U21039 ( .A(_02843__PTR3), .B(_02843__PTR19), .S(_01888__PTR4), .Z(_02847__PTR3) );
  MUX2_X1 U21040 ( .A(_02843__PTR4), .B(_02843__PTR20), .S(_01888__PTR4), .Z(_02847__PTR4) );
  MUX2_X1 U21041 ( .A(_02843__PTR5), .B(_02843__PTR21), .S(_01888__PTR4), .Z(_02847__PTR5) );
  MUX2_X1 U21042 ( .A(_02843__PTR6), .B(_02843__PTR22), .S(_01888__PTR4), .Z(_02847__PTR6) );
  MUX2_X1 U21043 ( .A(_02843__PTR7), .B(_02843__PTR23), .S(_01888__PTR4), .Z(_02847__PTR7) );
  MUX2_X1 U21044 ( .A(_02843__PTR32), .B(_02843__PTR48), .S(_01888__PTR4), .Z(_02847__PTR32) );
  MUX2_X1 U21045 ( .A(_02843__PTR33), .B(_02843__PTR49), .S(_01888__PTR4), .Z(_02847__PTR33) );
  MUX2_X1 U21046 ( .A(_02843__PTR34), .B(_02843__PTR50), .S(_01888__PTR4), .Z(_02847__PTR34) );
  MUX2_X1 U21047 ( .A(_02843__PTR35), .B(_02843__PTR51), .S(_01888__PTR4), .Z(_02847__PTR35) );
  MUX2_X1 U21048 ( .A(_02843__PTR36), .B(_02843__PTR52), .S(_01888__PTR4), .Z(_02847__PTR36) );
  MUX2_X1 U21049 ( .A(_02843__PTR37), .B(_02843__PTR53), .S(_01888__PTR4), .Z(_02847__PTR37) );
  MUX2_X1 U21050 ( .A(_02843__PTR38), .B(_02843__PTR54), .S(_01888__PTR4), .Z(_02847__PTR38) );
  MUX2_X1 U21051 ( .A(_02843__PTR39), .B(_02843__PTR55), .S(_01888__PTR4), .Z(_02847__PTR39) );
  MUX2_X1 U21052 ( .A(_02843__PTR64), .B(_02843__PTR80), .S(_01888__PTR4), .Z(_02847__PTR64) );
  MUX2_X1 U21053 ( .A(_02843__PTR65), .B(_02843__PTR81), .S(_01888__PTR4), .Z(_02847__PTR65) );
  MUX2_X1 U21054 ( .A(_02843__PTR66), .B(_02843__PTR82), .S(_01888__PTR4), .Z(_02847__PTR66) );
  MUX2_X1 U21055 ( .A(_02843__PTR67), .B(_02843__PTR83), .S(_01888__PTR4), .Z(_02847__PTR67) );
  MUX2_X1 U21056 ( .A(_02843__PTR68), .B(_02843__PTR84), .S(_01888__PTR4), .Z(_02847__PTR68) );
  MUX2_X1 U21057 ( .A(_02843__PTR69), .B(_02843__PTR85), .S(_01888__PTR4), .Z(_02847__PTR69) );
  MUX2_X1 U21058 ( .A(_02843__PTR70), .B(_02843__PTR86), .S(_01888__PTR4), .Z(_02847__PTR70) );
  MUX2_X1 U21059 ( .A(_02843__PTR71), .B(_02843__PTR87), .S(_01888__PTR4), .Z(_02847__PTR71) );
  MUX2_X1 U21060 ( .A(_02843__PTR96), .B(_02843__PTR112), .S(_01888__PTR4), .Z(_02847__PTR96) );
  MUX2_X1 U21061 ( .A(_02843__PTR97), .B(_02843__PTR113), .S(_01888__PTR4), .Z(_02847__PTR97) );
  MUX2_X1 U21062 ( .A(_02843__PTR98), .B(_02843__PTR114), .S(_01888__PTR4), .Z(_02847__PTR98) );
  MUX2_X1 U21063 ( .A(_02843__PTR99), .B(_02843__PTR115), .S(_01888__PTR4), .Z(_02847__PTR99) );
  MUX2_X1 U21064 ( .A(_02843__PTR100), .B(_02843__PTR116), .S(_01888__PTR4), .Z(_02847__PTR100) );
  MUX2_X1 U21065 ( .A(_02843__PTR101), .B(_02843__PTR117), .S(_01888__PTR4), .Z(_02847__PTR101) );
  MUX2_X1 U21066 ( .A(_02843__PTR102), .B(_02843__PTR118), .S(_01888__PTR4), .Z(_02847__PTR102) );
  MUX2_X1 U21067 ( .A(_02843__PTR103), .B(_02843__PTR119), .S(_01888__PTR4), .Z(_02847__PTR103) );
  MUX2_X1 U21068 ( .A(_02850__PTR0), .B(_02850__PTR64), .S(_01890__PTR6), .Z(_01891__PTR0) );
  MUX2_X1 U21069 ( .A(_02850__PTR1), .B(_02850__PTR65), .S(_01890__PTR6), .Z(_01891__PTR1) );
  MUX2_X1 U21070 ( .A(_02850__PTR2), .B(_02850__PTR66), .S(_01890__PTR6), .Z(_01891__PTR2) );
  MUX2_X1 U21071 ( .A(_02850__PTR3), .B(_02850__PTR67), .S(_01890__PTR6), .Z(_01891__PTR3) );
  MUX2_X1 U21072 ( .A(_02850__PTR4), .B(_02850__PTR68), .S(_01890__PTR6), .Z(_01891__PTR4) );
  MUX2_X1 U21073 ( .A(_02850__PTR5), .B(_02850__PTR69), .S(_01890__PTR6), .Z(_01891__PTR5) );
  MUX2_X1 U21074 ( .A(_02850__PTR6), .B(_02850__PTR70), .S(_01890__PTR6), .Z(_01891__PTR6) );
  MUX2_X1 U21075 ( .A(_02850__PTR7), .B(_02850__PTR71), .S(_01890__PTR6), .Z(_01891__PTR7) );
  MUX2_X1 U21076 ( .A(_02849__PTR0), .B(_02849__PTR32), .S(_01890__PTR5), .Z(_02850__PTR0) );
  MUX2_X1 U21077 ( .A(_02849__PTR1), .B(_02849__PTR33), .S(_01890__PTR5), .Z(_02850__PTR1) );
  MUX2_X1 U21078 ( .A(_02849__PTR2), .B(_02849__PTR34), .S(_01890__PTR5), .Z(_02850__PTR2) );
  MUX2_X1 U21079 ( .A(_02849__PTR3), .B(_02849__PTR35), .S(_01890__PTR5), .Z(_02850__PTR3) );
  MUX2_X1 U21080 ( .A(_02849__PTR4), .B(_02849__PTR36), .S(_01890__PTR5), .Z(_02850__PTR4) );
  MUX2_X1 U21081 ( .A(_02849__PTR5), .B(_02849__PTR37), .S(_01890__PTR5), .Z(_02850__PTR5) );
  MUX2_X1 U21082 ( .A(_02849__PTR6), .B(_02849__PTR38), .S(_01890__PTR5), .Z(_02850__PTR6) );
  MUX2_X1 U21083 ( .A(_02849__PTR7), .B(_02849__PTR39), .S(_01890__PTR5), .Z(_02850__PTR7) );
  MUX2_X1 U21084 ( .A(_02849__PTR64), .B(_02849__PTR96), .S(_01890__PTR5), .Z(_02850__PTR64) );
  MUX2_X1 U21085 ( .A(_02849__PTR65), .B(_02849__PTR97), .S(_01890__PTR5), .Z(_02850__PTR65) );
  MUX2_X1 U21086 ( .A(_02849__PTR66), .B(_02849__PTR98), .S(_01890__PTR5), .Z(_02850__PTR66) );
  MUX2_X1 U21087 ( .A(_02849__PTR67), .B(_02849__PTR99), .S(_01890__PTR5), .Z(_02850__PTR67) );
  MUX2_X1 U21088 ( .A(_02849__PTR68), .B(_02849__PTR100), .S(_01890__PTR5), .Z(_02850__PTR68) );
  MUX2_X1 U21089 ( .A(_02849__PTR69), .B(_02849__PTR101), .S(_01890__PTR5), .Z(_02850__PTR69) );
  MUX2_X1 U21090 ( .A(_02849__PTR70), .B(_02849__PTR102), .S(_01890__PTR5), .Z(_02850__PTR70) );
  MUX2_X1 U21091 ( .A(_02849__PTR71), .B(_02849__PTR103), .S(_01890__PTR5), .Z(_02850__PTR71) );
  MUX2_X1 U21092 ( .A(_02840__PTR16), .B(_02840__PTR0), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR0) );
  MUX2_X1 U21093 ( .A(_02840__PTR17), .B(_02840__PTR1), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR1) );
  MUX2_X1 U21094 ( .A(_02840__PTR18), .B(_02840__PTR2), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR2) );
  MUX2_X1 U21095 ( .A(_02840__PTR19), .B(_02840__PTR3), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR3) );
  MUX2_X1 U21096 ( .A(_02840__PTR20), .B(_02840__PTR4), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR4) );
  MUX2_X1 U21097 ( .A(_02840__PTR21), .B(_02840__PTR5), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR5) );
  MUX2_X1 U21098 ( .A(_02840__PTR22), .B(_02840__PTR6), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR6) );
  MUX2_X1 U21099 ( .A(_02840__PTR23), .B(_02840__PTR7), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR7) );
  MUX2_X1 U21100 ( .A(_02840__PTR48), .B(_02840__PTR32), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR32) );
  MUX2_X1 U21101 ( .A(_02840__PTR49), .B(_02840__PTR33), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR33) );
  MUX2_X1 U21102 ( .A(_02840__PTR50), .B(_02840__PTR34), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR34) );
  MUX2_X1 U21103 ( .A(_02840__PTR51), .B(_02840__PTR35), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR35) );
  MUX2_X1 U21104 ( .A(_02840__PTR52), .B(_02840__PTR36), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR36) );
  MUX2_X1 U21105 ( .A(_02840__PTR53), .B(_02840__PTR37), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR37) );
  MUX2_X1 U21106 ( .A(_02840__PTR54), .B(_02840__PTR38), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR38) );
  MUX2_X1 U21107 ( .A(_02840__PTR55), .B(_02840__PTR39), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR39) );
  MUX2_X1 U21108 ( .A(_02840__PTR80), .B(_02840__PTR64), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR64) );
  MUX2_X1 U21109 ( .A(_02840__PTR81), .B(_02840__PTR65), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR65) );
  MUX2_X1 U21110 ( .A(_02840__PTR82), .B(_02840__PTR66), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR66) );
  MUX2_X1 U21111 ( .A(_02840__PTR83), .B(_02840__PTR67), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR67) );
  MUX2_X1 U21112 ( .A(_02840__PTR84), .B(_02840__PTR68), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR68) );
  MUX2_X1 U21113 ( .A(_02840__PTR85), .B(_02840__PTR69), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR69) );
  MUX2_X1 U21114 ( .A(_02840__PTR86), .B(_02840__PTR70), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR70) );
  MUX2_X1 U21115 ( .A(_02840__PTR87), .B(_02840__PTR71), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR71) );
  MUX2_X1 U21116 ( .A(_02840__PTR112), .B(_02840__PTR96), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR96) );
  MUX2_X1 U21117 ( .A(_02840__PTR113), .B(_02840__PTR97), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR97) );
  MUX2_X1 U21118 ( .A(_02840__PTR114), .B(_02840__PTR98), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR98) );
  MUX2_X1 U21119 ( .A(_02840__PTR115), .B(_02840__PTR99), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR99) );
  MUX2_X1 U21120 ( .A(_02840__PTR116), .B(_02840__PTR100), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR100) );
  MUX2_X1 U21121 ( .A(_02840__PTR117), .B(_02840__PTR101), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR101) );
  MUX2_X1 U21122 ( .A(_02840__PTR118), .B(_02840__PTR102), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR102) );
  MUX2_X1 U21123 ( .A(_02840__PTR119), .B(_02840__PTR103), .S(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02849__PTR103) );
  MUX2_X1 U21124 ( .A(_02852__PTR0), .B(_02852__PTR128), .S(P1_P1_State2_PTR2), .Z(_02853__PTR0) );
  MUX2_X1 U21125 ( .A(_02852__PTR1), .B(_02852__PTR129), .S(P1_P1_State2_PTR2), .Z(_02853__PTR1) );
  MUX2_X1 U21126 ( .A(_02852__PTR2), .B(_02852__PTR130), .S(P1_P1_State2_PTR2), .Z(_02853__PTR2) );
  MUX2_X1 U21127 ( .A(_02852__PTR3), .B(_02852__PTR131), .S(P1_P1_State2_PTR2), .Z(_02853__PTR3) );
  MUX2_X1 U21128 ( .A(_02852__PTR4), .B(_02852__PTR132), .S(P1_P1_State2_PTR2), .Z(_02853__PTR4) );
  MUX2_X1 U21129 ( .A(_02852__PTR5), .B(_02852__PTR133), .S(P1_P1_State2_PTR2), .Z(_02853__PTR5) );
  MUX2_X1 U21130 ( .A(_02852__PTR6), .B(_02852__PTR134), .S(P1_P1_State2_PTR2), .Z(_02853__PTR6) );
  MUX2_X1 U21131 ( .A(_02852__PTR7), .B(_02852__PTR135), .S(P1_P1_State2_PTR2), .Z(_02853__PTR7) );
  MUX2_X1 U21132 ( .A(_02852__PTR8), .B(_02852__PTR136), .S(P1_P1_State2_PTR2), .Z(_02853__PTR8) );
  MUX2_X1 U21133 ( .A(_02852__PTR9), .B(_02852__PTR137), .S(P1_P1_State2_PTR2), .Z(_02853__PTR9) );
  MUX2_X1 U21134 ( .A(_02852__PTR10), .B(_02852__PTR138), .S(P1_P1_State2_PTR2), .Z(_02853__PTR10) );
  MUX2_X1 U21135 ( .A(_02852__PTR11), .B(_02852__PTR139), .S(P1_P1_State2_PTR2), .Z(_02853__PTR11) );
  MUX2_X1 U21136 ( .A(_02852__PTR12), .B(_02852__PTR140), .S(P1_P1_State2_PTR2), .Z(_02853__PTR12) );
  MUX2_X1 U21137 ( .A(_02852__PTR13), .B(_02852__PTR141), .S(P1_P1_State2_PTR2), .Z(_02853__PTR13) );
  MUX2_X1 U21138 ( .A(_02852__PTR14), .B(_02852__PTR142), .S(P1_P1_State2_PTR2), .Z(_02853__PTR14) );
  MUX2_X1 U21139 ( .A(_02852__PTR15), .B(_02852__PTR143), .S(P1_P1_State2_PTR2), .Z(_02853__PTR15) );
  MUX2_X1 U21140 ( .A(_02852__PTR16), .B(_02852__PTR144), .S(P1_P1_State2_PTR2), .Z(_02853__PTR16) );
  MUX2_X1 U21141 ( .A(_02852__PTR17), .B(_02852__PTR145), .S(P1_P1_State2_PTR2), .Z(_02853__PTR17) );
  MUX2_X1 U21142 ( .A(_02852__PTR18), .B(_02852__PTR146), .S(P1_P1_State2_PTR2), .Z(_02853__PTR18) );
  MUX2_X1 U21143 ( .A(_02852__PTR19), .B(_02852__PTR147), .S(P1_P1_State2_PTR2), .Z(_02853__PTR19) );
  MUX2_X1 U21144 ( .A(_02852__PTR20), .B(_02852__PTR148), .S(P1_P1_State2_PTR2), .Z(_02853__PTR20) );
  MUX2_X1 U21145 ( .A(_02852__PTR21), .B(_02852__PTR149), .S(P1_P1_State2_PTR2), .Z(_02853__PTR21) );
  MUX2_X1 U21146 ( .A(_02852__PTR22), .B(_02852__PTR150), .S(P1_P1_State2_PTR2), .Z(_02853__PTR22) );
  MUX2_X1 U21147 ( .A(_02852__PTR23), .B(_02852__PTR151), .S(P1_P1_State2_PTR2), .Z(_02853__PTR23) );
  MUX2_X1 U21148 ( .A(_02852__PTR24), .B(_02852__PTR152), .S(P1_P1_State2_PTR2), .Z(_02853__PTR24) );
  MUX2_X1 U21149 ( .A(_02852__PTR25), .B(_02852__PTR153), .S(P1_P1_State2_PTR2), .Z(_02853__PTR25) );
  MUX2_X1 U21150 ( .A(_02852__PTR26), .B(_02852__PTR154), .S(P1_P1_State2_PTR2), .Z(_02853__PTR26) );
  MUX2_X1 U21151 ( .A(_02852__PTR27), .B(_02852__PTR155), .S(P1_P1_State2_PTR2), .Z(_02853__PTR27) );
  MUX2_X1 U21152 ( .A(_02852__PTR28), .B(_02852__PTR156), .S(P1_P1_State2_PTR2), .Z(_02853__PTR28) );
  MUX2_X1 U21153 ( .A(_02852__PTR29), .B(_02852__PTR157), .S(P1_P1_State2_PTR2), .Z(_02853__PTR29) );
  MUX2_X1 U21154 ( .A(_02852__PTR30), .B(_02852__PTR158), .S(P1_P1_State2_PTR2), .Z(_02853__PTR30) );
  MUX2_X1 U21155 ( .A(_02852__PTR31), .B(_02852__PTR159), .S(P1_P1_State2_PTR2), .Z(_02853__PTR31) );
  MUX2_X1 U21156 ( .A(_02851__PTR0), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR0) );
  MUX2_X1 U21157 ( .A(_02851__PTR1), .B(_02851__PTR65), .S(P1_P1_State2_PTR1), .Z(_02852__PTR1) );
  MUX2_X1 U21158 ( .A(_02851__PTR2), .B(_02851__PTR66), .S(P1_P1_State2_PTR1), .Z(_02852__PTR2) );
  MUX2_X1 U21159 ( .A(_02851__PTR3), .B(_02851__PTR67), .S(P1_P1_State2_PTR1), .Z(_02852__PTR3) );
  MUX2_X1 U21160 ( .A(_02851__PTR4), .B(_02851__PTR68), .S(P1_P1_State2_PTR1), .Z(_02852__PTR4) );
  MUX2_X1 U21161 ( .A(_02851__PTR5), .B(_02851__PTR69), .S(P1_P1_State2_PTR1), .Z(_02852__PTR5) );
  MUX2_X1 U21162 ( .A(_02851__PTR6), .B(_02851__PTR70), .S(P1_P1_State2_PTR1), .Z(_02852__PTR6) );
  MUX2_X1 U21163 ( .A(_02851__PTR7), .B(_02851__PTR71), .S(P1_P1_State2_PTR1), .Z(_02852__PTR7) );
  MUX2_X1 U21164 ( .A(_02851__PTR8), .B(_02851__PTR72), .S(P1_P1_State2_PTR1), .Z(_02852__PTR8) );
  MUX2_X1 U21165 ( .A(_02851__PTR9), .B(_02851__PTR73), .S(P1_P1_State2_PTR1), .Z(_02852__PTR9) );
  MUX2_X1 U21166 ( .A(_02851__PTR10), .B(_02851__PTR74), .S(P1_P1_State2_PTR1), .Z(_02852__PTR10) );
  MUX2_X1 U21167 ( .A(_02851__PTR11), .B(_02851__PTR75), .S(P1_P1_State2_PTR1), .Z(_02852__PTR11) );
  MUX2_X1 U21168 ( .A(_02851__PTR12), .B(_02851__PTR76), .S(P1_P1_State2_PTR1), .Z(_02852__PTR12) );
  MUX2_X1 U21169 ( .A(_02851__PTR13), .B(_02851__PTR77), .S(P1_P1_State2_PTR1), .Z(_02852__PTR13) );
  MUX2_X1 U21170 ( .A(_02851__PTR14), .B(_02851__PTR78), .S(P1_P1_State2_PTR1), .Z(_02852__PTR14) );
  MUX2_X1 U21171 ( .A(_02851__PTR15), .B(_02851__PTR79), .S(P1_P1_State2_PTR1), .Z(_02852__PTR15) );
  MUX2_X1 U21172 ( .A(_02851__PTR16), .B(_02851__PTR80), .S(P1_P1_State2_PTR1), .Z(_02852__PTR16) );
  MUX2_X1 U21173 ( .A(_02851__PTR17), .B(_02851__PTR81), .S(P1_P1_State2_PTR1), .Z(_02852__PTR17) );
  MUX2_X1 U21174 ( .A(_02851__PTR18), .B(_02851__PTR82), .S(P1_P1_State2_PTR1), .Z(_02852__PTR18) );
  MUX2_X1 U21175 ( .A(_02851__PTR19), .B(_02851__PTR83), .S(P1_P1_State2_PTR1), .Z(_02852__PTR19) );
  MUX2_X1 U21176 ( .A(_02851__PTR20), .B(_02851__PTR84), .S(P1_P1_State2_PTR1), .Z(_02852__PTR20) );
  MUX2_X1 U21177 ( .A(_02851__PTR21), .B(_02851__PTR85), .S(P1_P1_State2_PTR1), .Z(_02852__PTR21) );
  MUX2_X1 U21178 ( .A(_02851__PTR22), .B(_02851__PTR86), .S(P1_P1_State2_PTR1), .Z(_02852__PTR22) );
  MUX2_X1 U21179 ( .A(_02851__PTR23), .B(_02851__PTR87), .S(P1_P1_State2_PTR1), .Z(_02852__PTR23) );
  MUX2_X1 U21180 ( .A(_02851__PTR24), .B(_02851__PTR88), .S(P1_P1_State2_PTR1), .Z(_02852__PTR24) );
  MUX2_X1 U21181 ( .A(_02851__PTR25), .B(_02851__PTR89), .S(P1_P1_State2_PTR1), .Z(_02852__PTR25) );
  MUX2_X1 U21182 ( .A(_02851__PTR26), .B(_02851__PTR90), .S(P1_P1_State2_PTR1), .Z(_02852__PTR26) );
  MUX2_X1 U21183 ( .A(_02851__PTR27), .B(_02851__PTR91), .S(P1_P1_State2_PTR1), .Z(_02852__PTR27) );
  MUX2_X1 U21184 ( .A(_02851__PTR28), .B(_02851__PTR92), .S(P1_P1_State2_PTR1), .Z(_02852__PTR28) );
  MUX2_X1 U21185 ( .A(_02851__PTR29), .B(_02851__PTR93), .S(P1_P1_State2_PTR1), .Z(_02852__PTR29) );
  MUX2_X1 U21186 ( .A(_02851__PTR30), .B(_02851__PTR94), .S(P1_P1_State2_PTR1), .Z(_02852__PTR30) );
  MUX2_X1 U21187 ( .A(_02851__PTR31), .B(_02851__PTR95), .S(P1_P1_State2_PTR1), .Z(_02852__PTR31) );
  MUX2_X1 U21188 ( .A(_02851__PTR128), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR128) );
  MUX2_X1 U21189 ( .A(_02851__PTR129), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR129) );
  MUX2_X1 U21190 ( .A(_02851__PTR130), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR130) );
  MUX2_X1 U21191 ( .A(_02851__PTR131), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR131) );
  MUX2_X1 U21192 ( .A(_02851__PTR132), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR132) );
  MUX2_X1 U21193 ( .A(_02851__PTR133), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR133) );
  MUX2_X1 U21194 ( .A(_02851__PTR134), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR134) );
  MUX2_X1 U21195 ( .A(_02851__PTR135), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR135) );
  MUX2_X1 U21196 ( .A(_02851__PTR136), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR136) );
  MUX2_X1 U21197 ( .A(_02851__PTR137), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR137) );
  MUX2_X1 U21198 ( .A(_02851__PTR138), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR138) );
  MUX2_X1 U21199 ( .A(_02851__PTR139), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR139) );
  MUX2_X1 U21200 ( .A(_02851__PTR140), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR140) );
  MUX2_X1 U21201 ( .A(_02851__PTR141), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR141) );
  MUX2_X1 U21202 ( .A(_02851__PTR142), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR142) );
  MUX2_X1 U21203 ( .A(_02851__PTR143), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR143) );
  MUX2_X1 U21204 ( .A(_02851__PTR144), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR144) );
  MUX2_X1 U21205 ( .A(_02851__PTR145), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR145) );
  MUX2_X1 U21206 ( .A(_02851__PTR146), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR146) );
  MUX2_X1 U21207 ( .A(_02851__PTR147), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR147) );
  MUX2_X1 U21208 ( .A(_02851__PTR148), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR148) );
  MUX2_X1 U21209 ( .A(_02851__PTR149), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR149) );
  MUX2_X1 U21210 ( .A(_02851__PTR150), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR150) );
  MUX2_X1 U21211 ( .A(_02851__PTR151), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR151) );
  MUX2_X1 U21212 ( .A(_02851__PTR152), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR152) );
  MUX2_X1 U21213 ( .A(_02851__PTR153), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR153) );
  MUX2_X1 U21214 ( .A(_02851__PTR154), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR154) );
  MUX2_X1 U21215 ( .A(_02851__PTR155), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR155) );
  MUX2_X1 U21216 ( .A(_02851__PTR156), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR156) );
  MUX2_X1 U21217 ( .A(_02851__PTR157), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR157) );
  MUX2_X1 U21218 ( .A(_02851__PTR158), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR158) );
  MUX2_X1 U21219 ( .A(_02851__PTR159), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02852__PTR159) );
  MUX2_X1 U21220 ( .A(P1_rEIP_PTR0), .B(P1_P1_PhyAddrPointer_PTR0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR0) );
  MUX2_X1 U21221 ( .A(P1_rEIP_PTR1), .B(P1_P1_PhyAddrPointer_PTR1), .S(P1_P1_State2_PTR0), .Z(_02851__PTR1) );
  MUX2_X1 U21222 ( .A(P1_rEIP_PTR2), .B(P1_P1_PhyAddrPointer_PTR2), .S(P1_P1_State2_PTR0), .Z(_02851__PTR2) );
  MUX2_X1 U21223 ( .A(P1_rEIP_PTR3), .B(P1_P1_PhyAddrPointer_PTR3), .S(P1_P1_State2_PTR0), .Z(_02851__PTR3) );
  MUX2_X1 U21224 ( .A(P1_rEIP_PTR4), .B(P1_P1_PhyAddrPointer_PTR4), .S(P1_P1_State2_PTR0), .Z(_02851__PTR4) );
  MUX2_X1 U21225 ( .A(P1_rEIP_PTR5), .B(P1_P1_PhyAddrPointer_PTR5), .S(P1_P1_State2_PTR0), .Z(_02851__PTR5) );
  MUX2_X1 U21226 ( .A(P1_rEIP_PTR6), .B(P1_P1_PhyAddrPointer_PTR6), .S(P1_P1_State2_PTR0), .Z(_02851__PTR6) );
  MUX2_X1 U21227 ( .A(P1_rEIP_PTR7), .B(P1_P1_PhyAddrPointer_PTR7), .S(P1_P1_State2_PTR0), .Z(_02851__PTR7) );
  MUX2_X1 U21228 ( .A(P1_rEIP_PTR8), .B(P1_P1_PhyAddrPointer_PTR8), .S(P1_P1_State2_PTR0), .Z(_02851__PTR8) );
  MUX2_X1 U21229 ( .A(P1_rEIP_PTR9), .B(P1_P1_PhyAddrPointer_PTR9), .S(P1_P1_State2_PTR0), .Z(_02851__PTR9) );
  MUX2_X1 U21230 ( .A(P1_rEIP_PTR10), .B(P1_P1_PhyAddrPointer_PTR10), .S(P1_P1_State2_PTR0), .Z(_02851__PTR10) );
  MUX2_X1 U21231 ( .A(P1_rEIP_PTR11), .B(P1_P1_PhyAddrPointer_PTR11), .S(P1_P1_State2_PTR0), .Z(_02851__PTR11) );
  MUX2_X1 U21232 ( .A(P1_rEIP_PTR12), .B(P1_P1_PhyAddrPointer_PTR12), .S(P1_P1_State2_PTR0), .Z(_02851__PTR12) );
  MUX2_X1 U21233 ( .A(P1_rEIP_PTR13), .B(P1_P1_PhyAddrPointer_PTR13), .S(P1_P1_State2_PTR0), .Z(_02851__PTR13) );
  MUX2_X1 U21234 ( .A(P1_rEIP_PTR14), .B(P1_P1_PhyAddrPointer_PTR14), .S(P1_P1_State2_PTR0), .Z(_02851__PTR14) );
  MUX2_X1 U21235 ( .A(P1_rEIP_PTR15), .B(P1_P1_PhyAddrPointer_PTR15), .S(P1_P1_State2_PTR0), .Z(_02851__PTR15) );
  MUX2_X1 U21236 ( .A(P1_rEIP_PTR16), .B(P1_P1_PhyAddrPointer_PTR16), .S(P1_P1_State2_PTR0), .Z(_02851__PTR16) );
  MUX2_X1 U21237 ( .A(P1_rEIP_PTR17), .B(P1_P1_PhyAddrPointer_PTR17), .S(P1_P1_State2_PTR0), .Z(_02851__PTR17) );
  MUX2_X1 U21238 ( .A(P1_rEIP_PTR18), .B(P1_P1_PhyAddrPointer_PTR18), .S(P1_P1_State2_PTR0), .Z(_02851__PTR18) );
  MUX2_X1 U21239 ( .A(P1_rEIP_PTR19), .B(P1_P1_PhyAddrPointer_PTR19), .S(P1_P1_State2_PTR0), .Z(_02851__PTR19) );
  MUX2_X1 U21240 ( .A(P1_rEIP_PTR20), .B(P1_P1_PhyAddrPointer_PTR20), .S(P1_P1_State2_PTR0), .Z(_02851__PTR20) );
  MUX2_X1 U21241 ( .A(P1_rEIP_PTR21), .B(P1_P1_PhyAddrPointer_PTR21), .S(P1_P1_State2_PTR0), .Z(_02851__PTR21) );
  MUX2_X1 U21242 ( .A(P1_rEIP_PTR22), .B(P1_P1_PhyAddrPointer_PTR22), .S(P1_P1_State2_PTR0), .Z(_02851__PTR22) );
  MUX2_X1 U21243 ( .A(P1_rEIP_PTR23), .B(P1_P1_PhyAddrPointer_PTR23), .S(P1_P1_State2_PTR0), .Z(_02851__PTR23) );
  MUX2_X1 U21244 ( .A(P1_rEIP_PTR24), .B(P1_P1_PhyAddrPointer_PTR24), .S(P1_P1_State2_PTR0), .Z(_02851__PTR24) );
  MUX2_X1 U21245 ( .A(P1_rEIP_PTR25), .B(P1_P1_PhyAddrPointer_PTR25), .S(P1_P1_State2_PTR0), .Z(_02851__PTR25) );
  MUX2_X1 U21246 ( .A(P1_rEIP_PTR26), .B(P1_P1_PhyAddrPointer_PTR26), .S(P1_P1_State2_PTR0), .Z(_02851__PTR26) );
  MUX2_X1 U21247 ( .A(P1_rEIP_PTR27), .B(P1_P1_PhyAddrPointer_PTR27), .S(P1_P1_State2_PTR0), .Z(_02851__PTR27) );
  MUX2_X1 U21248 ( .A(P1_rEIP_PTR28), .B(P1_P1_PhyAddrPointer_PTR28), .S(P1_P1_State2_PTR0), .Z(_02851__PTR28) );
  MUX2_X1 U21249 ( .A(P1_rEIP_PTR29), .B(P1_P1_PhyAddrPointer_PTR29), .S(P1_P1_State2_PTR0), .Z(_02851__PTR29) );
  MUX2_X1 U21250 ( .A(P1_rEIP_PTR30), .B(P1_P1_PhyAddrPointer_PTR30), .S(P1_P1_State2_PTR0), .Z(_02851__PTR30) );
  MUX2_X1 U21251 ( .A(P1_rEIP_PTR31), .B(P1_P1_PhyAddrPointer_PTR31), .S(P1_P1_State2_PTR0), .Z(_02851__PTR31) );
  MUX2_X1 U21252 ( .A(_01892__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR65) );
  MUX2_X1 U21253 ( .A(_01892__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR66) );
  MUX2_X1 U21254 ( .A(_01892__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR67) );
  MUX2_X1 U21255 ( .A(_01892__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR68) );
  MUX2_X1 U21256 ( .A(_01892__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR69) );
  MUX2_X1 U21257 ( .A(_01892__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR70) );
  MUX2_X1 U21258 ( .A(_01892__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR71) );
  MUX2_X1 U21259 ( .A(_01892__PTR72), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR72) );
  MUX2_X1 U21260 ( .A(_01892__PTR73), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR73) );
  MUX2_X1 U21261 ( .A(_01892__PTR74), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR74) );
  MUX2_X1 U21262 ( .A(_01892__PTR75), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR75) );
  MUX2_X1 U21263 ( .A(_01892__PTR76), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR76) );
  MUX2_X1 U21264 ( .A(_01892__PTR77), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR77) );
  MUX2_X1 U21265 ( .A(_01892__PTR78), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR78) );
  MUX2_X1 U21266 ( .A(_01892__PTR79), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR79) );
  MUX2_X1 U21267 ( .A(_01892__PTR80), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR80) );
  MUX2_X1 U21268 ( .A(_01892__PTR81), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR81) );
  MUX2_X1 U21269 ( .A(_01892__PTR82), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR82) );
  MUX2_X1 U21270 ( .A(_01892__PTR83), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR83) );
  MUX2_X1 U21271 ( .A(_01892__PTR84), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR84) );
  MUX2_X1 U21272 ( .A(_01892__PTR85), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR85) );
  MUX2_X1 U21273 ( .A(_01892__PTR86), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR86) );
  MUX2_X1 U21274 ( .A(_01892__PTR87), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR87) );
  MUX2_X1 U21275 ( .A(_01892__PTR88), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR88) );
  MUX2_X1 U21276 ( .A(_01892__PTR89), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR89) );
  MUX2_X1 U21277 ( .A(_01892__PTR90), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR90) );
  MUX2_X1 U21278 ( .A(_01892__PTR91), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR91) );
  MUX2_X1 U21279 ( .A(_01892__PTR92), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR92) );
  MUX2_X1 U21280 ( .A(_01892__PTR93), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR93) );
  MUX2_X1 U21281 ( .A(_01892__PTR94), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR94) );
  MUX2_X1 U21282 ( .A(_01892__PTR95), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02851__PTR95) );
  MUX2_X1 U21283 ( .A(1'b0), .B(_01892__PTR160), .S(P1_P1_State2_PTR0), .Z(_02851__PTR128) );
  MUX2_X1 U21284 ( .A(_01892__PTR129), .B(_01892__PTR161), .S(P1_P1_State2_PTR0), .Z(_02851__PTR129) );
  MUX2_X1 U21285 ( .A(_01892__PTR130), .B(_01892__PTR162), .S(P1_P1_State2_PTR0), .Z(_02851__PTR130) );
  MUX2_X1 U21286 ( .A(_01892__PTR131), .B(_01892__PTR163), .S(P1_P1_State2_PTR0), .Z(_02851__PTR131) );
  MUX2_X1 U21287 ( .A(_01892__PTR132), .B(_01892__PTR164), .S(P1_P1_State2_PTR0), .Z(_02851__PTR132) );
  MUX2_X1 U21288 ( .A(_01892__PTR133), .B(_01892__PTR165), .S(P1_P1_State2_PTR0), .Z(_02851__PTR133) );
  MUX2_X1 U21289 ( .A(_01892__PTR134), .B(_01892__PTR166), .S(P1_P1_State2_PTR0), .Z(_02851__PTR134) );
  MUX2_X1 U21290 ( .A(_01892__PTR135), .B(_01892__PTR167), .S(P1_P1_State2_PTR0), .Z(_02851__PTR135) );
  MUX2_X1 U21291 ( .A(_01892__PTR136), .B(_01892__PTR168), .S(P1_P1_State2_PTR0), .Z(_02851__PTR136) );
  MUX2_X1 U21292 ( .A(_01892__PTR137), .B(_01892__PTR169), .S(P1_P1_State2_PTR0), .Z(_02851__PTR137) );
  MUX2_X1 U21293 ( .A(_01892__PTR138), .B(_01892__PTR170), .S(P1_P1_State2_PTR0), .Z(_02851__PTR138) );
  MUX2_X1 U21294 ( .A(_01892__PTR139), .B(_01892__PTR171), .S(P1_P1_State2_PTR0), .Z(_02851__PTR139) );
  MUX2_X1 U21295 ( .A(_01892__PTR140), .B(_01892__PTR172), .S(P1_P1_State2_PTR0), .Z(_02851__PTR140) );
  MUX2_X1 U21296 ( .A(_01892__PTR141), .B(_01892__PTR173), .S(P1_P1_State2_PTR0), .Z(_02851__PTR141) );
  MUX2_X1 U21297 ( .A(_01892__PTR142), .B(_01892__PTR174), .S(P1_P1_State2_PTR0), .Z(_02851__PTR142) );
  MUX2_X1 U21298 ( .A(_01892__PTR143), .B(_01892__PTR175), .S(P1_P1_State2_PTR0), .Z(_02851__PTR143) );
  MUX2_X1 U21299 ( .A(_01892__PTR144), .B(_01892__PTR176), .S(P1_P1_State2_PTR0), .Z(_02851__PTR144) );
  MUX2_X1 U21300 ( .A(_01892__PTR145), .B(_01892__PTR177), .S(P1_P1_State2_PTR0), .Z(_02851__PTR145) );
  MUX2_X1 U21301 ( .A(_01892__PTR146), .B(_01892__PTR178), .S(P1_P1_State2_PTR0), .Z(_02851__PTR146) );
  MUX2_X1 U21302 ( .A(_01892__PTR147), .B(_01892__PTR179), .S(P1_P1_State2_PTR0), .Z(_02851__PTR147) );
  MUX2_X1 U21303 ( .A(_01892__PTR148), .B(_01892__PTR180), .S(P1_P1_State2_PTR0), .Z(_02851__PTR148) );
  MUX2_X1 U21304 ( .A(_01892__PTR149), .B(_01892__PTR181), .S(P1_P1_State2_PTR0), .Z(_02851__PTR149) );
  MUX2_X1 U21305 ( .A(_01892__PTR150), .B(_01892__PTR182), .S(P1_P1_State2_PTR0), .Z(_02851__PTR150) );
  MUX2_X1 U21306 ( .A(_01892__PTR151), .B(_01892__PTR183), .S(P1_P1_State2_PTR0), .Z(_02851__PTR151) );
  MUX2_X1 U21307 ( .A(_01892__PTR152), .B(_01892__PTR184), .S(P1_P1_State2_PTR0), .Z(_02851__PTR152) );
  MUX2_X1 U21308 ( .A(_01892__PTR153), .B(_01892__PTR185), .S(P1_P1_State2_PTR0), .Z(_02851__PTR153) );
  MUX2_X1 U21309 ( .A(_01892__PTR154), .B(_01892__PTR186), .S(P1_P1_State2_PTR0), .Z(_02851__PTR154) );
  MUX2_X1 U21310 ( .A(_01892__PTR155), .B(_01892__PTR187), .S(P1_P1_State2_PTR0), .Z(_02851__PTR155) );
  MUX2_X1 U21311 ( .A(_01892__PTR156), .B(_01892__PTR188), .S(P1_P1_State2_PTR0), .Z(_02851__PTR156) );
  MUX2_X1 U21312 ( .A(_01892__PTR157), .B(_01892__PTR189), .S(P1_P1_State2_PTR0), .Z(_02851__PTR157) );
  MUX2_X1 U21313 ( .A(_01892__PTR158), .B(_01892__PTR190), .S(P1_P1_State2_PTR0), .Z(_02851__PTR158) );
  MUX2_X1 U21314 ( .A(_01892__PTR159), .B(_01892__PTR191), .S(P1_P1_State2_PTR0), .Z(_02851__PTR159) );
  MUX2_X1 U21315 ( .A(_02855__PTR0), .B(_02855__PTR128), .S(P1_P1_State2_PTR2), .Z(_02856__PTR0) );
  MUX2_X1 U21316 ( .A(_02855__PTR1), .B(_02855__PTR129), .S(P1_P1_State2_PTR2), .Z(_02856__PTR1) );
  MUX2_X1 U21317 ( .A(_02855__PTR2), .B(_02855__PTR130), .S(P1_P1_State2_PTR2), .Z(_02856__PTR2) );
  MUX2_X1 U21318 ( .A(_02855__PTR3), .B(_02855__PTR131), .S(P1_P1_State2_PTR2), .Z(_02856__PTR3) );
  MUX2_X1 U21319 ( .A(_02855__PTR4), .B(_02855__PTR132), .S(P1_P1_State2_PTR2), .Z(_02856__PTR4) );
  MUX2_X1 U21320 ( .A(_02855__PTR5), .B(_02855__PTR133), .S(P1_P1_State2_PTR2), .Z(_02856__PTR5) );
  MUX2_X1 U21321 ( .A(_02855__PTR6), .B(_02855__PTR134), .S(P1_P1_State2_PTR2), .Z(_02856__PTR6) );
  MUX2_X1 U21322 ( .A(_02855__PTR7), .B(_02855__PTR135), .S(P1_P1_State2_PTR2), .Z(_02856__PTR7) );
  MUX2_X1 U21323 ( .A(_02855__PTR8), .B(_02855__PTR136), .S(P1_P1_State2_PTR2), .Z(_02856__PTR8) );
  MUX2_X1 U21324 ( .A(_02855__PTR9), .B(_02855__PTR137), .S(P1_P1_State2_PTR2), .Z(_02856__PTR9) );
  MUX2_X1 U21325 ( .A(_02855__PTR10), .B(_02855__PTR138), .S(P1_P1_State2_PTR2), .Z(_02856__PTR10) );
  MUX2_X1 U21326 ( .A(_02855__PTR11), .B(_02855__PTR139), .S(P1_P1_State2_PTR2), .Z(_02856__PTR11) );
  MUX2_X1 U21327 ( .A(_02855__PTR12), .B(_02855__PTR140), .S(P1_P1_State2_PTR2), .Z(_02856__PTR12) );
  MUX2_X1 U21328 ( .A(_02855__PTR13), .B(_02855__PTR141), .S(P1_P1_State2_PTR2), .Z(_02856__PTR13) );
  MUX2_X1 U21329 ( .A(_02855__PTR14), .B(_02855__PTR142), .S(P1_P1_State2_PTR2), .Z(_02856__PTR14) );
  MUX2_X1 U21330 ( .A(_02855__PTR15), .B(_02855__PTR143), .S(P1_P1_State2_PTR2), .Z(_02856__PTR15) );
  MUX2_X1 U21331 ( .A(_02855__PTR16), .B(_02855__PTR144), .S(P1_P1_State2_PTR2), .Z(_02856__PTR16) );
  MUX2_X1 U21332 ( .A(_02855__PTR17), .B(_02855__PTR145), .S(P1_P1_State2_PTR2), .Z(_02856__PTR17) );
  MUX2_X1 U21333 ( .A(_02855__PTR18), .B(_02855__PTR146), .S(P1_P1_State2_PTR2), .Z(_02856__PTR18) );
  MUX2_X1 U21334 ( .A(_02855__PTR19), .B(_02855__PTR147), .S(P1_P1_State2_PTR2), .Z(_02856__PTR19) );
  MUX2_X1 U21335 ( .A(_02855__PTR20), .B(_02855__PTR148), .S(P1_P1_State2_PTR2), .Z(_02856__PTR20) );
  MUX2_X1 U21336 ( .A(_02855__PTR21), .B(_02855__PTR149), .S(P1_P1_State2_PTR2), .Z(_02856__PTR21) );
  MUX2_X1 U21337 ( .A(_02855__PTR22), .B(_02855__PTR150), .S(P1_P1_State2_PTR2), .Z(_02856__PTR22) );
  MUX2_X1 U21338 ( .A(_02855__PTR23), .B(_02855__PTR151), .S(P1_P1_State2_PTR2), .Z(_02856__PTR23) );
  MUX2_X1 U21339 ( .A(_02855__PTR24), .B(_02855__PTR152), .S(P1_P1_State2_PTR2), .Z(_02856__PTR24) );
  MUX2_X1 U21340 ( .A(_02855__PTR25), .B(_02855__PTR153), .S(P1_P1_State2_PTR2), .Z(_02856__PTR25) );
  MUX2_X1 U21341 ( .A(_02855__PTR26), .B(_02855__PTR154), .S(P1_P1_State2_PTR2), .Z(_02856__PTR26) );
  MUX2_X1 U21342 ( .A(_02855__PTR27), .B(_02855__PTR155), .S(P1_P1_State2_PTR2), .Z(_02856__PTR27) );
  MUX2_X1 U21343 ( .A(_02855__PTR28), .B(_02855__PTR156), .S(P1_P1_State2_PTR2), .Z(_02856__PTR28) );
  MUX2_X1 U21344 ( .A(_02855__PTR29), .B(_02855__PTR157), .S(P1_P1_State2_PTR2), .Z(_02856__PTR29) );
  MUX2_X1 U21345 ( .A(_02855__PTR30), .B(_02855__PTR158), .S(P1_P1_State2_PTR2), .Z(_02856__PTR30) );
  MUX2_X1 U21346 ( .A(_02855__PTR31), .B(_02855__PTR159), .S(P1_P1_State2_PTR2), .Z(_02856__PTR31) );
  MUX2_X1 U21347 ( .A(_02854__PTR0), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR0) );
  MUX2_X1 U21348 ( .A(_02854__PTR1), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR1) );
  MUX2_X1 U21349 ( .A(_02854__PTR2), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR2) );
  MUX2_X1 U21350 ( .A(_02854__PTR3), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR3) );
  MUX2_X1 U21351 ( .A(_02854__PTR4), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR4) );
  MUX2_X1 U21352 ( .A(_02854__PTR5), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR5) );
  MUX2_X1 U21353 ( .A(_02854__PTR6), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR6) );
  MUX2_X1 U21354 ( .A(_02854__PTR7), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR7) );
  MUX2_X1 U21355 ( .A(_02854__PTR8), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR8) );
  MUX2_X1 U21356 ( .A(_02854__PTR9), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR9) );
  MUX2_X1 U21357 ( .A(_02854__PTR10), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR10) );
  MUX2_X1 U21358 ( .A(_02854__PTR11), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR11) );
  MUX2_X1 U21359 ( .A(_02854__PTR12), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR12) );
  MUX2_X1 U21360 ( .A(_02854__PTR13), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR13) );
  MUX2_X1 U21361 ( .A(_02854__PTR14), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR14) );
  MUX2_X1 U21362 ( .A(_02854__PTR15), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR15) );
  MUX2_X1 U21363 ( .A(_02854__PTR16), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR16) );
  MUX2_X1 U21364 ( .A(_02854__PTR17), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR17) );
  MUX2_X1 U21365 ( .A(_02854__PTR18), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR18) );
  MUX2_X1 U21366 ( .A(_02854__PTR19), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR19) );
  MUX2_X1 U21367 ( .A(_02854__PTR20), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR20) );
  MUX2_X1 U21368 ( .A(_02854__PTR21), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR21) );
  MUX2_X1 U21369 ( .A(_02854__PTR22), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR22) );
  MUX2_X1 U21370 ( .A(_02854__PTR23), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR23) );
  MUX2_X1 U21371 ( .A(_02854__PTR24), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR24) );
  MUX2_X1 U21372 ( .A(_02854__PTR25), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR25) );
  MUX2_X1 U21373 ( .A(_02854__PTR26), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR26) );
  MUX2_X1 U21374 ( .A(_02854__PTR27), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR27) );
  MUX2_X1 U21375 ( .A(_02854__PTR28), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR28) );
  MUX2_X1 U21376 ( .A(_02854__PTR29), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR29) );
  MUX2_X1 U21377 ( .A(_02854__PTR30), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR30) );
  MUX2_X1 U21378 ( .A(_02854__PTR31), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR31) );
  MUX2_X1 U21379 ( .A(_02854__PTR128), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR128) );
  MUX2_X1 U21380 ( .A(_02854__PTR129), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR129) );
  MUX2_X1 U21381 ( .A(_02854__PTR130), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR130) );
  MUX2_X1 U21382 ( .A(_02854__PTR131), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR131) );
  MUX2_X1 U21383 ( .A(_02854__PTR132), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR132) );
  MUX2_X1 U21384 ( .A(_02854__PTR133), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR133) );
  MUX2_X1 U21385 ( .A(_02854__PTR134), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR134) );
  MUX2_X1 U21386 ( .A(_02854__PTR135), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR135) );
  MUX2_X1 U21387 ( .A(_02854__PTR136), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR136) );
  MUX2_X1 U21388 ( .A(_02854__PTR137), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR137) );
  MUX2_X1 U21389 ( .A(_02854__PTR138), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR138) );
  MUX2_X1 U21390 ( .A(_02854__PTR139), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR139) );
  MUX2_X1 U21391 ( .A(_02854__PTR140), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR140) );
  MUX2_X1 U21392 ( .A(_02854__PTR141), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR141) );
  MUX2_X1 U21393 ( .A(_02854__PTR142), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR142) );
  MUX2_X1 U21394 ( .A(_02854__PTR143), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR143) );
  MUX2_X1 U21395 ( .A(_02854__PTR144), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR144) );
  MUX2_X1 U21396 ( .A(_02854__PTR145), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR145) );
  MUX2_X1 U21397 ( .A(_02854__PTR146), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR146) );
  MUX2_X1 U21398 ( .A(_02854__PTR147), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR147) );
  MUX2_X1 U21399 ( .A(_02854__PTR148), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR148) );
  MUX2_X1 U21400 ( .A(_02854__PTR149), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR149) );
  MUX2_X1 U21401 ( .A(_02854__PTR150), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR150) );
  MUX2_X1 U21402 ( .A(_02854__PTR151), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR151) );
  MUX2_X1 U21403 ( .A(_02854__PTR152), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR152) );
  MUX2_X1 U21404 ( .A(_02854__PTR153), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR153) );
  MUX2_X1 U21405 ( .A(_02854__PTR154), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR154) );
  MUX2_X1 U21406 ( .A(_02854__PTR155), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR155) );
  MUX2_X1 U21407 ( .A(_02854__PTR156), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR156) );
  MUX2_X1 U21408 ( .A(_02854__PTR157), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR157) );
  MUX2_X1 U21409 ( .A(_02854__PTR158), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR158) );
  MUX2_X1 U21410 ( .A(_02854__PTR159), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02855__PTR159) );
  MUX2_X1 U21411 ( .A(P1_rEIP_PTR0), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR0) );
  MUX2_X1 U21412 ( .A(P1_rEIP_PTR1), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR1) );
  MUX2_X1 U21413 ( .A(P1_rEIP_PTR2), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR2) );
  MUX2_X1 U21414 ( .A(P1_rEIP_PTR3), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR3) );
  MUX2_X1 U21415 ( .A(P1_rEIP_PTR4), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR4) );
  MUX2_X1 U21416 ( .A(P1_rEIP_PTR5), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR5) );
  MUX2_X1 U21417 ( .A(P1_rEIP_PTR6), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR6) );
  MUX2_X1 U21418 ( .A(P1_rEIP_PTR7), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR7) );
  MUX2_X1 U21419 ( .A(P1_rEIP_PTR8), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR8) );
  MUX2_X1 U21420 ( .A(P1_rEIP_PTR9), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR9) );
  MUX2_X1 U21421 ( .A(P1_rEIP_PTR10), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR10) );
  MUX2_X1 U21422 ( .A(P1_rEIP_PTR11), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR11) );
  MUX2_X1 U21423 ( .A(P1_rEIP_PTR12), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR12) );
  MUX2_X1 U21424 ( .A(P1_rEIP_PTR13), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR13) );
  MUX2_X1 U21425 ( .A(P1_rEIP_PTR14), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR14) );
  MUX2_X1 U21426 ( .A(P1_rEIP_PTR15), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR15) );
  MUX2_X1 U21427 ( .A(P1_rEIP_PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR16) );
  MUX2_X1 U21428 ( .A(P1_rEIP_PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR17) );
  MUX2_X1 U21429 ( .A(P1_rEIP_PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR18) );
  MUX2_X1 U21430 ( .A(P1_rEIP_PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR19) );
  MUX2_X1 U21431 ( .A(P1_rEIP_PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR20) );
  MUX2_X1 U21432 ( .A(P1_rEIP_PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR21) );
  MUX2_X1 U21433 ( .A(P1_rEIP_PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR22) );
  MUX2_X1 U21434 ( .A(P1_rEIP_PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR23) );
  MUX2_X1 U21435 ( .A(P1_rEIP_PTR24), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR24) );
  MUX2_X1 U21436 ( .A(P1_rEIP_PTR25), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR25) );
  MUX2_X1 U21437 ( .A(P1_rEIP_PTR26), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR26) );
  MUX2_X1 U21438 ( .A(P1_rEIP_PTR27), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR27) );
  MUX2_X1 U21439 ( .A(P1_rEIP_PTR28), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR28) );
  MUX2_X1 U21440 ( .A(P1_rEIP_PTR29), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR29) );
  MUX2_X1 U21441 ( .A(P1_rEIP_PTR30), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR30) );
  MUX2_X1 U21442 ( .A(P1_rEIP_PTR31), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02854__PTR31) );
  MUX2_X1 U21443 ( .A(1'b0), .B(_01893__PTR160), .S(P1_P1_State2_PTR0), .Z(_02854__PTR128) );
  MUX2_X1 U21444 ( .A(1'b0), .B(_01893__PTR161), .S(P1_P1_State2_PTR0), .Z(_02854__PTR129) );
  MUX2_X1 U21445 ( .A(1'b0), .B(_01893__PTR162), .S(P1_P1_State2_PTR0), .Z(_02854__PTR130) );
  MUX2_X1 U21446 ( .A(1'b0), .B(_01893__PTR163), .S(P1_P1_State2_PTR0), .Z(_02854__PTR131) );
  MUX2_X1 U21447 ( .A(1'b0), .B(_01893__PTR164), .S(P1_P1_State2_PTR0), .Z(_02854__PTR132) );
  MUX2_X1 U21448 ( .A(1'b0), .B(_01893__PTR165), .S(P1_P1_State2_PTR0), .Z(_02854__PTR133) );
  MUX2_X1 U21449 ( .A(1'b0), .B(_01893__PTR166), .S(P1_P1_State2_PTR0), .Z(_02854__PTR134) );
  MUX2_X1 U21450 ( .A(1'b0), .B(_01893__PTR167), .S(P1_P1_State2_PTR0), .Z(_02854__PTR135) );
  MUX2_X1 U21451 ( .A(1'b0), .B(_01893__PTR168), .S(P1_P1_State2_PTR0), .Z(_02854__PTR136) );
  MUX2_X1 U21452 ( .A(1'b0), .B(_01893__PTR169), .S(P1_P1_State2_PTR0), .Z(_02854__PTR137) );
  MUX2_X1 U21453 ( .A(1'b0), .B(_01893__PTR170), .S(P1_P1_State2_PTR0), .Z(_02854__PTR138) );
  MUX2_X1 U21454 ( .A(1'b0), .B(_01893__PTR171), .S(P1_P1_State2_PTR0), .Z(_02854__PTR139) );
  MUX2_X1 U21455 ( .A(1'b0), .B(_01893__PTR172), .S(P1_P1_State2_PTR0), .Z(_02854__PTR140) );
  MUX2_X1 U21456 ( .A(1'b0), .B(_01893__PTR173), .S(P1_P1_State2_PTR0), .Z(_02854__PTR141) );
  MUX2_X1 U21457 ( .A(1'b0), .B(_01893__PTR174), .S(P1_P1_State2_PTR0), .Z(_02854__PTR142) );
  MUX2_X1 U21458 ( .A(1'b0), .B(_01893__PTR175), .S(P1_P1_State2_PTR0), .Z(_02854__PTR143) );
  MUX2_X1 U21459 ( .A(1'b0), .B(_01893__PTR176), .S(P1_P1_State2_PTR0), .Z(_02854__PTR144) );
  MUX2_X1 U21460 ( .A(1'b0), .B(_01893__PTR177), .S(P1_P1_State2_PTR0), .Z(_02854__PTR145) );
  MUX2_X1 U21461 ( .A(1'b0), .B(_01893__PTR178), .S(P1_P1_State2_PTR0), .Z(_02854__PTR146) );
  MUX2_X1 U21462 ( .A(1'b0), .B(_01893__PTR179), .S(P1_P1_State2_PTR0), .Z(_02854__PTR147) );
  MUX2_X1 U21463 ( .A(1'b0), .B(_01893__PTR180), .S(P1_P1_State2_PTR0), .Z(_02854__PTR148) );
  MUX2_X1 U21464 ( .A(1'b0), .B(_01893__PTR181), .S(P1_P1_State2_PTR0), .Z(_02854__PTR149) );
  MUX2_X1 U21465 ( .A(1'b0), .B(_01893__PTR182), .S(P1_P1_State2_PTR0), .Z(_02854__PTR150) );
  MUX2_X1 U21466 ( .A(1'b0), .B(_01893__PTR183), .S(P1_P1_State2_PTR0), .Z(_02854__PTR151) );
  MUX2_X1 U21467 ( .A(1'b0), .B(_01893__PTR184), .S(P1_P1_State2_PTR0), .Z(_02854__PTR152) );
  MUX2_X1 U21468 ( .A(1'b0), .B(_01893__PTR185), .S(P1_P1_State2_PTR0), .Z(_02854__PTR153) );
  MUX2_X1 U21469 ( .A(1'b0), .B(_01893__PTR186), .S(P1_P1_State2_PTR0), .Z(_02854__PTR154) );
  MUX2_X1 U21470 ( .A(1'b0), .B(_01893__PTR187), .S(P1_P1_State2_PTR0), .Z(_02854__PTR155) );
  MUX2_X1 U21471 ( .A(1'b0), .B(_01893__PTR188), .S(P1_P1_State2_PTR0), .Z(_02854__PTR156) );
  MUX2_X1 U21472 ( .A(1'b0), .B(_01893__PTR189), .S(P1_P1_State2_PTR0), .Z(_02854__PTR157) );
  MUX2_X1 U21473 ( .A(1'b0), .B(_01893__PTR190), .S(P1_P1_State2_PTR0), .Z(_02854__PTR158) );
  MUX2_X1 U21474 ( .A(1'b0), .B(_01893__PTR191), .S(P1_P1_State2_PTR0), .Z(_02854__PTR159) );
  MUX2_X1 U21475 ( .A(_02859__PTR0), .B(_02857__PTR32), .S(P1_P1_State2_PTR3), .Z(_01895__PTR0) );
  MUX2_X1 U21476 ( .A(_02859__PTR1), .B(1'b0), .S(P1_P1_State2_PTR3), .Z(_01895__PTR1) );
  MUX2_X1 U21477 ( .A(_02859__PTR2), .B(1'b0), .S(P1_P1_State2_PTR3), .Z(_01895__PTR2) );
  MUX2_X1 U21478 ( .A(_02859__PTR3), .B(_00302_), .S(P1_P1_State2_PTR3), .Z(_01895__PTR3) );
  MUX2_X1 U21479 ( .A(_02857__PTR0), .B(_02857__PTR16), .S(P1_P1_State2_PTR2), .Z(_02859__PTR0) );
  MUX2_X1 U21480 ( .A(_02857__PTR1), .B(_02857__PTR17), .S(P1_P1_State2_PTR2), .Z(_02859__PTR1) );
  MUX2_X1 U21481 ( .A(_02857__PTR2), .B(_02857__PTR18), .S(P1_P1_State2_PTR2), .Z(_02859__PTR2) );
  MUX2_X1 U21482 ( .A(1'b0), .B(_02857__PTR19), .S(P1_P1_State2_PTR2), .Z(_02859__PTR3) );
  MUX2_X1 U21483 ( .A(_02860__PTR1), .B(_02858__PTR1), .S(P1_P1_State2_PTR1), .Z(_02857__PTR1) );
  MUX2_X1 U21484 ( .A(1'b0), .B(_02858__PTR2), .S(P1_P1_State2_PTR1), .Z(_02857__PTR2) );
  MUX2_X1 U21485 ( .A(_02858__PTR8), .B(_02858__PTR16), .S(P1_P1_State2_PTR1), .Z(_02857__PTR16) );
  MUX2_X1 U21486 ( .A(_02858__PTR9), .B(_02858__PTR17), .S(P1_P1_State2_PTR1), .Z(_02857__PTR17) );
  MUX2_X1 U21487 ( .A(_02858__PTR10), .B(_02858__PTR18), .S(P1_P1_State2_PTR1), .Z(_02857__PTR18) );
  MUX2_X1 U21488 ( .A(_02858__PTR11), .B(_02858__PTR19), .S(P1_P1_State2_PTR1), .Z(_02857__PTR19) );
  MUX2_X1 U21489 ( .A(1'b0), .B(_01894__PTR14), .S(P1_P1_State2_PTR0), .Z(_02860__PTR1) );
  MUX2_X1 U21490 ( .A(1'b1), .B(P1_READY_n), .S(P1_P1_State2_PTR0), .Z(_02857__PTR0) );
  MUX2_X1 U21491 ( .A(_01894__PTR9), .B(P1_READY_n), .S(P1_P1_State2_PTR0), .Z(_02858__PTR1) );
  MUX2_X1 U21492 ( .A(P1_StateBS16), .B(_01894__PTR14), .S(P1_P1_State2_PTR0), .Z(_02858__PTR2) );
  MUX2_X1 U21493 ( .A(1'b1), .B(_01894__PTR20), .S(P1_P1_State2_PTR0), .Z(_02858__PTR8) );
  MUX2_X1 U21494 ( .A(1'b0), .B(_01894__PTR21), .S(P1_P1_State2_PTR0), .Z(_02858__PTR9) );
  MUX2_X1 U21495 ( .A(1'b1), .B(_01894__PTR22), .S(P1_P1_State2_PTR0), .Z(_02858__PTR10) );
  MUX2_X1 U21496 ( .A(1'b0), .B(_01894__PTR23), .S(P1_P1_State2_PTR0), .Z(_02858__PTR11) );
  MUX2_X1 U21497 ( .A(_01894__PTR26), .B(_01894__PTR28), .S(P1_P1_State2_PTR0), .Z(_02858__PTR16) );
  MUX2_X1 U21498 ( .A(_01849__PTR6), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02858__PTR17) );
  MUX2_X1 U21499 ( .A(_01894__PTR26), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02858__PTR18) );
  MUX2_X1 U21500 ( .A(_01849__PTR6), .B(1'b1), .S(P1_P1_State2_PTR0), .Z(_02858__PTR19) );
  MUX2_X1 U21501 ( .A(_01894__PTR32), .B(1'b1), .S(P1_P1_State2_PTR0), .Z(_02857__PTR32) );
  MUX2_X1 U21502 ( .A(_02861__PTR32), .B(_02861__PTR128), .S(P1_P1_State2_PTR1), .Z(_02862__PTR0) );
  MUX2_X1 U21503 ( .A(_02861__PTR32), .B(_02861__PTR129), .S(P1_P1_State2_PTR1), .Z(_02862__PTR1) );
  MUX2_X1 U21504 ( .A(_02861__PTR32), .B(_02861__PTR130), .S(P1_P1_State2_PTR1), .Z(_02862__PTR2) );
  MUX2_X1 U21505 ( .A(_02861__PTR32), .B(_02861__PTR131), .S(P1_P1_State2_PTR1), .Z(_02862__PTR3) );
  MUX2_X1 U21506 ( .A(_02861__PTR19), .B(_02861__PTR132), .S(P1_P1_State2_PTR1), .Z(_02862__PTR4) );
  MUX2_X1 U21507 ( .A(_02861__PTR19), .B(_02861__PTR133), .S(P1_P1_State2_PTR1), .Z(_02862__PTR5) );
  MUX2_X1 U21508 ( .A(_02861__PTR19), .B(_02861__PTR134), .S(P1_P1_State2_PTR1), .Z(_02862__PTR6) );
  MUX2_X1 U21509 ( .A(_02861__PTR19), .B(_02861__PTR135), .S(P1_P1_State2_PTR1), .Z(_02862__PTR7) );
  MUX2_X1 U21510 ( .A(_02861__PTR19), .B(_02861__PTR136), .S(P1_P1_State2_PTR1), .Z(_02862__PTR8) );
  MUX2_X1 U21511 ( .A(_02861__PTR19), .B(_02861__PTR137), .S(P1_P1_State2_PTR1), .Z(_02862__PTR9) );
  MUX2_X1 U21512 ( .A(_02861__PTR19), .B(_02861__PTR138), .S(P1_P1_State2_PTR1), .Z(_02862__PTR10) );
  MUX2_X1 U21513 ( .A(_02861__PTR19), .B(_02861__PTR139), .S(P1_P1_State2_PTR1), .Z(_02862__PTR11) );
  MUX2_X1 U21514 ( .A(_02861__PTR19), .B(_02861__PTR140), .S(P1_P1_State2_PTR1), .Z(_02862__PTR12) );
  MUX2_X1 U21515 ( .A(_02861__PTR19), .B(_02861__PTR141), .S(P1_P1_State2_PTR1), .Z(_02862__PTR13) );
  MUX2_X1 U21516 ( .A(_02861__PTR19), .B(_02861__PTR142), .S(P1_P1_State2_PTR1), .Z(_02862__PTR14) );
  MUX2_X1 U21517 ( .A(_02861__PTR19), .B(_02861__PTR143), .S(P1_P1_State2_PTR1), .Z(_02862__PTR15) );
  MUX2_X1 U21518 ( .A(_02861__PTR19), .B(_02861__PTR144), .S(P1_P1_State2_PTR1), .Z(_02862__PTR16) );
  MUX2_X1 U21519 ( .A(_02861__PTR19), .B(_02861__PTR145), .S(P1_P1_State2_PTR1), .Z(_02862__PTR17) );
  MUX2_X1 U21520 ( .A(_02861__PTR19), .B(_02861__PTR146), .S(P1_P1_State2_PTR1), .Z(_02862__PTR18) );
  MUX2_X1 U21521 ( .A(_02861__PTR19), .B(_02861__PTR147), .S(P1_P1_State2_PTR1), .Z(_02862__PTR19) );
  MUX2_X1 U21522 ( .A(_02861__PTR32), .B(_02861__PTR148), .S(P1_P1_State2_PTR1), .Z(_02862__PTR20) );
  MUX2_X1 U21523 ( .A(_02861__PTR32), .B(_02861__PTR149), .S(P1_P1_State2_PTR1), .Z(_02862__PTR21) );
  MUX2_X1 U21524 ( .A(_02861__PTR32), .B(_02861__PTR150), .S(P1_P1_State2_PTR1), .Z(_02862__PTR22) );
  MUX2_X1 U21525 ( .A(_02861__PTR32), .B(_02861__PTR151), .S(P1_P1_State2_PTR1), .Z(_02862__PTR23) );
  MUX2_X1 U21526 ( .A(_02861__PTR32), .B(_02861__PTR152), .S(P1_P1_State2_PTR1), .Z(_02862__PTR24) );
  MUX2_X1 U21527 ( .A(_02861__PTR32), .B(_02861__PTR153), .S(P1_P1_State2_PTR1), .Z(_02862__PTR25) );
  MUX2_X1 U21528 ( .A(_02861__PTR32), .B(_02861__PTR154), .S(P1_P1_State2_PTR1), .Z(_02862__PTR26) );
  MUX2_X1 U21529 ( .A(_02861__PTR32), .B(_02861__PTR155), .S(P1_P1_State2_PTR1), .Z(_02862__PTR27) );
  MUX2_X1 U21530 ( .A(_02861__PTR32), .B(_02861__PTR156), .S(P1_P1_State2_PTR1), .Z(_02862__PTR28) );
  MUX2_X1 U21531 ( .A(_02861__PTR32), .B(_02861__PTR157), .S(P1_P1_State2_PTR1), .Z(_02862__PTR29) );
  MUX2_X1 U21532 ( .A(_02861__PTR32), .B(_02861__PTR158), .S(P1_P1_State2_PTR1), .Z(_02862__PTR30) );
  MUX2_X1 U21533 ( .A(_02861__PTR32), .B(_02861__PTR160), .S(P1_P1_State2_PTR1), .Z(_02862__PTR32) );
  MUX2_X1 U21534 ( .A(_02861__PTR256), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR256) );
  MUX2_X1 U21535 ( .A(_02861__PTR257), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR257) );
  MUX2_X1 U21536 ( .A(_02861__PTR258), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR258) );
  MUX2_X1 U21537 ( .A(_02861__PTR259), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR259) );
  MUX2_X1 U21538 ( .A(_02861__PTR260), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR260) );
  MUX2_X1 U21539 ( .A(_02861__PTR261), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR261) );
  MUX2_X1 U21540 ( .A(_02861__PTR262), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR262) );
  MUX2_X1 U21541 ( .A(_02861__PTR263), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR263) );
  MUX2_X1 U21542 ( .A(_02861__PTR264), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR264) );
  MUX2_X1 U21543 ( .A(_02861__PTR265), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR265) );
  MUX2_X1 U21544 ( .A(_02861__PTR266), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR266) );
  MUX2_X1 U21545 ( .A(_02861__PTR267), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR267) );
  MUX2_X1 U21546 ( .A(_02861__PTR268), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR268) );
  MUX2_X1 U21547 ( .A(_02861__PTR269), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR269) );
  MUX2_X1 U21548 ( .A(_02861__PTR270), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR270) );
  MUX2_X1 U21549 ( .A(_02861__PTR271), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR271) );
  MUX2_X1 U21550 ( .A(_02861__PTR272), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR272) );
  MUX2_X1 U21551 ( .A(_02861__PTR273), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR273) );
  MUX2_X1 U21552 ( .A(_02861__PTR274), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR274) );
  MUX2_X1 U21553 ( .A(_02861__PTR275), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR275) );
  MUX2_X1 U21554 ( .A(_02861__PTR276), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR276) );
  MUX2_X1 U21555 ( .A(_02861__PTR277), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR277) );
  MUX2_X1 U21556 ( .A(_02861__PTR278), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR278) );
  MUX2_X1 U21557 ( .A(_02861__PTR279), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR279) );
  MUX2_X1 U21558 ( .A(_02861__PTR280), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR280) );
  MUX2_X1 U21559 ( .A(_02861__PTR281), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR281) );
  MUX2_X1 U21560 ( .A(_02861__PTR282), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR282) );
  MUX2_X1 U21561 ( .A(_02861__PTR283), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR283) );
  MUX2_X1 U21562 ( .A(_02861__PTR284), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR284) );
  MUX2_X1 U21563 ( .A(_02861__PTR285), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR285) );
  MUX2_X1 U21564 ( .A(_02861__PTR286), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR286) );
  MUX2_X1 U21565 ( .A(_02861__PTR288), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02862__PTR288) );
  MUX2_X1 U21566 ( .A(1'b0), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR32) );
  MUX2_X1 U21567 ( .A(1'b1), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR19) );
  MUX2_X1 U21568 ( .A(_01896__PTR128), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR128) );
  MUX2_X1 U21569 ( .A(_01896__PTR129), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR129) );
  MUX2_X1 U21570 ( .A(_01896__PTR130), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR130) );
  MUX2_X1 U21571 ( .A(_01896__PTR131), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR131) );
  MUX2_X1 U21572 ( .A(_01896__PTR132), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR132) );
  MUX2_X1 U21573 ( .A(_01896__PTR133), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR133) );
  MUX2_X1 U21574 ( .A(_01896__PTR134), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR134) );
  MUX2_X1 U21575 ( .A(_01896__PTR135), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR135) );
  MUX2_X1 U21576 ( .A(_01896__PTR136), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR136) );
  MUX2_X1 U21577 ( .A(_01896__PTR137), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR137) );
  MUX2_X1 U21578 ( .A(_01896__PTR138), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR138) );
  MUX2_X1 U21579 ( .A(_01896__PTR139), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR139) );
  MUX2_X1 U21580 ( .A(_01896__PTR140), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR140) );
  MUX2_X1 U21581 ( .A(_01896__PTR141), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR141) );
  MUX2_X1 U21582 ( .A(_01896__PTR142), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR142) );
  MUX2_X1 U21583 ( .A(_01896__PTR143), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR143) );
  MUX2_X1 U21584 ( .A(_01896__PTR144), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR144) );
  MUX2_X1 U21585 ( .A(_01896__PTR145), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR145) );
  MUX2_X1 U21586 ( .A(_01896__PTR146), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR146) );
  MUX2_X1 U21587 ( .A(_01896__PTR147), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR147) );
  MUX2_X1 U21588 ( .A(_01896__PTR148), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR148) );
  MUX2_X1 U21589 ( .A(_01896__PTR149), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR149) );
  MUX2_X1 U21590 ( .A(_01896__PTR150), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR150) );
  MUX2_X1 U21591 ( .A(_01896__PTR151), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR151) );
  MUX2_X1 U21592 ( .A(_01896__PTR152), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR152) );
  MUX2_X1 U21593 ( .A(_01896__PTR153), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR153) );
  MUX2_X1 U21594 ( .A(_01896__PTR154), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR154) );
  MUX2_X1 U21595 ( .A(_01896__PTR155), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR155) );
  MUX2_X1 U21596 ( .A(_01896__PTR156), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR156) );
  MUX2_X1 U21597 ( .A(_01896__PTR157), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR157) );
  MUX2_X1 U21598 ( .A(_01896__PTR158), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR158) );
  MUX2_X1 U21599 ( .A(_01896__PTR160), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02861__PTR160) );
  MUX2_X1 U21600 ( .A(1'b0), .B(_01896__PTR320), .S(P1_P1_State2_PTR0), .Z(_02861__PTR256) );
  MUX2_X1 U21601 ( .A(1'b0), .B(_01896__PTR321), .S(P1_P1_State2_PTR0), .Z(_02861__PTR257) );
  MUX2_X1 U21602 ( .A(1'b0), .B(_01896__PTR322), .S(P1_P1_State2_PTR0), .Z(_02861__PTR258) );
  MUX2_X1 U21603 ( .A(1'b0), .B(_01896__PTR323), .S(P1_P1_State2_PTR0), .Z(_02861__PTR259) );
  MUX2_X1 U21604 ( .A(1'b0), .B(_01896__PTR324), .S(P1_P1_State2_PTR0), .Z(_02861__PTR260) );
  MUX2_X1 U21605 ( .A(1'b0), .B(_01896__PTR325), .S(P1_P1_State2_PTR0), .Z(_02861__PTR261) );
  MUX2_X1 U21606 ( .A(1'b0), .B(_01896__PTR326), .S(P1_P1_State2_PTR0), .Z(_02861__PTR262) );
  MUX2_X1 U21607 ( .A(1'b0), .B(_01896__PTR327), .S(P1_P1_State2_PTR0), .Z(_02861__PTR263) );
  MUX2_X1 U21608 ( .A(1'b0), .B(_01896__PTR328), .S(P1_P1_State2_PTR0), .Z(_02861__PTR264) );
  MUX2_X1 U21609 ( .A(1'b0), .B(_01896__PTR329), .S(P1_P1_State2_PTR0), .Z(_02861__PTR265) );
  MUX2_X1 U21610 ( .A(1'b0), .B(_01896__PTR330), .S(P1_P1_State2_PTR0), .Z(_02861__PTR266) );
  MUX2_X1 U21611 ( .A(1'b0), .B(_01896__PTR331), .S(P1_P1_State2_PTR0), .Z(_02861__PTR267) );
  MUX2_X1 U21612 ( .A(1'b0), .B(_01896__PTR332), .S(P1_P1_State2_PTR0), .Z(_02861__PTR268) );
  MUX2_X1 U21613 ( .A(1'b0), .B(_01896__PTR333), .S(P1_P1_State2_PTR0), .Z(_02861__PTR269) );
  MUX2_X1 U21614 ( .A(1'b0), .B(_01896__PTR334), .S(P1_P1_State2_PTR0), .Z(_02861__PTR270) );
  MUX2_X1 U21615 ( .A(1'b0), .B(_01896__PTR335), .S(P1_P1_State2_PTR0), .Z(_02861__PTR271) );
  MUX2_X1 U21616 ( .A(1'b0), .B(_01896__PTR336), .S(P1_P1_State2_PTR0), .Z(_02861__PTR272) );
  MUX2_X1 U21617 ( .A(1'b0), .B(_01896__PTR337), .S(P1_P1_State2_PTR0), .Z(_02861__PTR273) );
  MUX2_X1 U21618 ( .A(1'b0), .B(_01896__PTR338), .S(P1_P1_State2_PTR0), .Z(_02861__PTR274) );
  MUX2_X1 U21619 ( .A(1'b0), .B(_01896__PTR339), .S(P1_P1_State2_PTR0), .Z(_02861__PTR275) );
  MUX2_X1 U21620 ( .A(1'b0), .B(_01896__PTR340), .S(P1_P1_State2_PTR0), .Z(_02861__PTR276) );
  MUX2_X1 U21621 ( .A(1'b0), .B(_01896__PTR341), .S(P1_P1_State2_PTR0), .Z(_02861__PTR277) );
  MUX2_X1 U21622 ( .A(1'b0), .B(_01896__PTR342), .S(P1_P1_State2_PTR0), .Z(_02861__PTR278) );
  MUX2_X1 U21623 ( .A(1'b0), .B(_01896__PTR343), .S(P1_P1_State2_PTR0), .Z(_02861__PTR279) );
  MUX2_X1 U21624 ( .A(1'b0), .B(_01896__PTR344), .S(P1_P1_State2_PTR0), .Z(_02861__PTR280) );
  MUX2_X1 U21625 ( .A(1'b0), .B(_01896__PTR345), .S(P1_P1_State2_PTR0), .Z(_02861__PTR281) );
  MUX2_X1 U21626 ( .A(1'b0), .B(_01896__PTR346), .S(P1_P1_State2_PTR0), .Z(_02861__PTR282) );
  MUX2_X1 U21627 ( .A(1'b0), .B(_01896__PTR347), .S(P1_P1_State2_PTR0), .Z(_02861__PTR283) );
  MUX2_X1 U21628 ( .A(1'b0), .B(_01896__PTR348), .S(P1_P1_State2_PTR0), .Z(_02861__PTR284) );
  MUX2_X1 U21629 ( .A(1'b0), .B(_01896__PTR349), .S(P1_P1_State2_PTR0), .Z(_02861__PTR285) );
  MUX2_X1 U21630 ( .A(1'b0), .B(_01896__PTR350), .S(P1_P1_State2_PTR0), .Z(_02861__PTR286) );
  MUX2_X1 U21631 ( .A(1'b0), .B(_01896__PTR352), .S(P1_P1_State2_PTR0), .Z(_02861__PTR288) );
  MUX2_X1 U21632 ( .A(_02863__PTR0), .B(_02851__PTR0), .S(P1_P1_State2_PTR3), .Z(_01897__PTR0) );
  MUX2_X1 U21633 ( .A(_02863__PTR1), .B(_02851__PTR1), .S(P1_P1_State2_PTR3), .Z(_01897__PTR1) );
  MUX2_X1 U21634 ( .A(_02863__PTR2), .B(_02851__PTR2), .S(P1_P1_State2_PTR3), .Z(_01897__PTR2) );
  MUX2_X1 U21635 ( .A(_02863__PTR3), .B(_02851__PTR3), .S(P1_P1_State2_PTR3), .Z(_01897__PTR3) );
  MUX2_X1 U21636 ( .A(_02863__PTR4), .B(_02851__PTR4), .S(P1_P1_State2_PTR3), .Z(_01897__PTR4) );
  MUX2_X1 U21637 ( .A(_02863__PTR5), .B(_02851__PTR5), .S(P1_P1_State2_PTR3), .Z(_01897__PTR5) );
  MUX2_X1 U21638 ( .A(_02863__PTR6), .B(_02851__PTR6), .S(P1_P1_State2_PTR3), .Z(_01897__PTR6) );
  MUX2_X1 U21639 ( .A(_02863__PTR7), .B(_02851__PTR7), .S(P1_P1_State2_PTR3), .Z(_01897__PTR7) );
  MUX2_X1 U21640 ( .A(_02863__PTR8), .B(_02851__PTR8), .S(P1_P1_State2_PTR3), .Z(_01897__PTR8) );
  MUX2_X1 U21641 ( .A(_02863__PTR9), .B(_02851__PTR9), .S(P1_P1_State2_PTR3), .Z(_01897__PTR9) );
  MUX2_X1 U21642 ( .A(_02863__PTR10), .B(_02851__PTR10), .S(P1_P1_State2_PTR3), .Z(_01897__PTR10) );
  MUX2_X1 U21643 ( .A(_02863__PTR11), .B(_02851__PTR11), .S(P1_P1_State2_PTR3), .Z(_01897__PTR11) );
  MUX2_X1 U21644 ( .A(_02863__PTR12), .B(_02851__PTR12), .S(P1_P1_State2_PTR3), .Z(_01897__PTR12) );
  MUX2_X1 U21645 ( .A(_02863__PTR13), .B(_02851__PTR13), .S(P1_P1_State2_PTR3), .Z(_01897__PTR13) );
  MUX2_X1 U21646 ( .A(_02863__PTR14), .B(_02851__PTR14), .S(P1_P1_State2_PTR3), .Z(_01897__PTR14) );
  MUX2_X1 U21647 ( .A(_02863__PTR15), .B(_02851__PTR15), .S(P1_P1_State2_PTR3), .Z(_01897__PTR15) );
  MUX2_X1 U21648 ( .A(_02863__PTR16), .B(_02851__PTR16), .S(P1_P1_State2_PTR3), .Z(_01897__PTR16) );
  MUX2_X1 U21649 ( .A(_02863__PTR17), .B(_02851__PTR17), .S(P1_P1_State2_PTR3), .Z(_01897__PTR17) );
  MUX2_X1 U21650 ( .A(_02863__PTR18), .B(_02851__PTR18), .S(P1_P1_State2_PTR3), .Z(_01897__PTR18) );
  MUX2_X1 U21651 ( .A(_02863__PTR19), .B(_02851__PTR19), .S(P1_P1_State2_PTR3), .Z(_01897__PTR19) );
  MUX2_X1 U21652 ( .A(_02863__PTR20), .B(_02851__PTR20), .S(P1_P1_State2_PTR3), .Z(_01897__PTR20) );
  MUX2_X1 U21653 ( .A(_02863__PTR21), .B(_02851__PTR21), .S(P1_P1_State2_PTR3), .Z(_01897__PTR21) );
  MUX2_X1 U21654 ( .A(_02863__PTR22), .B(_02851__PTR22), .S(P1_P1_State2_PTR3), .Z(_01897__PTR22) );
  MUX2_X1 U21655 ( .A(_02863__PTR23), .B(_02851__PTR23), .S(P1_P1_State2_PTR3), .Z(_01897__PTR23) );
  MUX2_X1 U21656 ( .A(_02863__PTR24), .B(_02851__PTR24), .S(P1_P1_State2_PTR3), .Z(_01897__PTR24) );
  MUX2_X1 U21657 ( .A(_02863__PTR25), .B(_02851__PTR25), .S(P1_P1_State2_PTR3), .Z(_01897__PTR25) );
  MUX2_X1 U21658 ( .A(_02863__PTR26), .B(_02851__PTR26), .S(P1_P1_State2_PTR3), .Z(_01897__PTR26) );
  MUX2_X1 U21659 ( .A(_02863__PTR27), .B(_02851__PTR27), .S(P1_P1_State2_PTR3), .Z(_01897__PTR27) );
  MUX2_X1 U21660 ( .A(_02863__PTR28), .B(_02851__PTR28), .S(P1_P1_State2_PTR3), .Z(_01897__PTR28) );
  MUX2_X1 U21661 ( .A(_02863__PTR29), .B(_02851__PTR29), .S(P1_P1_State2_PTR3), .Z(_01897__PTR29) );
  MUX2_X1 U21662 ( .A(_02863__PTR30), .B(_02851__PTR30), .S(P1_P1_State2_PTR3), .Z(_01897__PTR30) );
  MUX2_X1 U21663 ( .A(_02863__PTR32), .B(_02851__PTR31), .S(P1_P1_State2_PTR3), .Z(_01897__PTR32) );
  MUX2_X1 U21664 ( .A(_02862__PTR0), .B(_02862__PTR256), .S(P1_P1_State2_PTR2), .Z(_02863__PTR0) );
  MUX2_X1 U21665 ( .A(_02862__PTR1), .B(_02862__PTR257), .S(P1_P1_State2_PTR2), .Z(_02863__PTR1) );
  MUX2_X1 U21666 ( .A(_02862__PTR2), .B(_02862__PTR258), .S(P1_P1_State2_PTR2), .Z(_02863__PTR2) );
  MUX2_X1 U21667 ( .A(_02862__PTR3), .B(_02862__PTR259), .S(P1_P1_State2_PTR2), .Z(_02863__PTR3) );
  MUX2_X1 U21668 ( .A(_02862__PTR4), .B(_02862__PTR260), .S(P1_P1_State2_PTR2), .Z(_02863__PTR4) );
  MUX2_X1 U21669 ( .A(_02862__PTR5), .B(_02862__PTR261), .S(P1_P1_State2_PTR2), .Z(_02863__PTR5) );
  MUX2_X1 U21670 ( .A(_02862__PTR6), .B(_02862__PTR262), .S(P1_P1_State2_PTR2), .Z(_02863__PTR6) );
  MUX2_X1 U21671 ( .A(_02862__PTR7), .B(_02862__PTR263), .S(P1_P1_State2_PTR2), .Z(_02863__PTR7) );
  MUX2_X1 U21672 ( .A(_02862__PTR8), .B(_02862__PTR264), .S(P1_P1_State2_PTR2), .Z(_02863__PTR8) );
  MUX2_X1 U21673 ( .A(_02862__PTR9), .B(_02862__PTR265), .S(P1_P1_State2_PTR2), .Z(_02863__PTR9) );
  MUX2_X1 U21674 ( .A(_02862__PTR10), .B(_02862__PTR266), .S(P1_P1_State2_PTR2), .Z(_02863__PTR10) );
  MUX2_X1 U21675 ( .A(_02862__PTR11), .B(_02862__PTR267), .S(P1_P1_State2_PTR2), .Z(_02863__PTR11) );
  MUX2_X1 U21676 ( .A(_02862__PTR12), .B(_02862__PTR268), .S(P1_P1_State2_PTR2), .Z(_02863__PTR12) );
  MUX2_X1 U21677 ( .A(_02862__PTR13), .B(_02862__PTR269), .S(P1_P1_State2_PTR2), .Z(_02863__PTR13) );
  MUX2_X1 U21678 ( .A(_02862__PTR14), .B(_02862__PTR270), .S(P1_P1_State2_PTR2), .Z(_02863__PTR14) );
  MUX2_X1 U21679 ( .A(_02862__PTR15), .B(_02862__PTR271), .S(P1_P1_State2_PTR2), .Z(_02863__PTR15) );
  MUX2_X1 U21680 ( .A(_02862__PTR16), .B(_02862__PTR272), .S(P1_P1_State2_PTR2), .Z(_02863__PTR16) );
  MUX2_X1 U21681 ( .A(_02862__PTR17), .B(_02862__PTR273), .S(P1_P1_State2_PTR2), .Z(_02863__PTR17) );
  MUX2_X1 U21682 ( .A(_02862__PTR18), .B(_02862__PTR274), .S(P1_P1_State2_PTR2), .Z(_02863__PTR18) );
  MUX2_X1 U21683 ( .A(_02862__PTR19), .B(_02862__PTR275), .S(P1_P1_State2_PTR2), .Z(_02863__PTR19) );
  MUX2_X1 U21684 ( .A(_02862__PTR20), .B(_02862__PTR276), .S(P1_P1_State2_PTR2), .Z(_02863__PTR20) );
  MUX2_X1 U21685 ( .A(_02862__PTR21), .B(_02862__PTR277), .S(P1_P1_State2_PTR2), .Z(_02863__PTR21) );
  MUX2_X1 U21686 ( .A(_02862__PTR22), .B(_02862__PTR278), .S(P1_P1_State2_PTR2), .Z(_02863__PTR22) );
  MUX2_X1 U21687 ( .A(_02862__PTR23), .B(_02862__PTR279), .S(P1_P1_State2_PTR2), .Z(_02863__PTR23) );
  MUX2_X1 U21688 ( .A(_02862__PTR24), .B(_02862__PTR280), .S(P1_P1_State2_PTR2), .Z(_02863__PTR24) );
  MUX2_X1 U21689 ( .A(_02862__PTR25), .B(_02862__PTR281), .S(P1_P1_State2_PTR2), .Z(_02863__PTR25) );
  MUX2_X1 U21690 ( .A(_02862__PTR26), .B(_02862__PTR282), .S(P1_P1_State2_PTR2), .Z(_02863__PTR26) );
  MUX2_X1 U21691 ( .A(_02862__PTR27), .B(_02862__PTR283), .S(P1_P1_State2_PTR2), .Z(_02863__PTR27) );
  MUX2_X1 U21692 ( .A(_02862__PTR28), .B(_02862__PTR284), .S(P1_P1_State2_PTR2), .Z(_02863__PTR28) );
  MUX2_X1 U21693 ( .A(_02862__PTR29), .B(_02862__PTR285), .S(P1_P1_State2_PTR2), .Z(_02863__PTR29) );
  MUX2_X1 U21694 ( .A(_02862__PTR30), .B(_02862__PTR286), .S(P1_P1_State2_PTR2), .Z(_02863__PTR30) );
  MUX2_X1 U21695 ( .A(_02862__PTR32), .B(_02862__PTR288), .S(P1_P1_State2_PTR2), .Z(_02863__PTR32) );
  MUX2_X1 U21696 ( .A(_02866__PTR0), .B(_02864__PTR64), .S(P1_P1_State2_PTR3), .Z(_01899__PTR0) );
  MUX2_X1 U21697 ( .A(_02866__PTR1), .B(_02864__PTR65), .S(P1_P1_State2_PTR3), .Z(_01899__PTR1) );
  MUX2_X1 U21698 ( .A(_02866__PTR2), .B(_02864__PTR66), .S(P1_P1_State2_PTR3), .Z(_01899__PTR2) );
  MUX2_X1 U21699 ( .A(_02866__PTR3), .B(_02864__PTR67), .S(P1_P1_State2_PTR3), .Z(_01899__PTR3) );
  MUX2_X1 U21700 ( .A(_02866__PTR4), .B(_02864__PTR68), .S(P1_P1_State2_PTR3), .Z(_01899__PTR4) );
  MUX2_X1 U21701 ( .A(_02866__PTR5), .B(_02864__PTR69), .S(P1_P1_State2_PTR3), .Z(_01899__PTR5) );
  MUX2_X1 U21702 ( .A(_02866__PTR6), .B(_02864__PTR70), .S(P1_P1_State2_PTR3), .Z(_01899__PTR6) );
  MUX2_X1 U21703 ( .A(_02866__PTR7), .B(_02864__PTR71), .S(P1_P1_State2_PTR3), .Z(_01899__PTR7) );
  MUX2_X1 U21704 ( .A(_02865__PTR0), .B(_02865__PTR32), .S(P1_P1_State2_PTR2), .Z(_02866__PTR0) );
  MUX2_X1 U21705 ( .A(_02865__PTR1), .B(_02865__PTR33), .S(P1_P1_State2_PTR2), .Z(_02866__PTR1) );
  MUX2_X1 U21706 ( .A(_02865__PTR2), .B(_02865__PTR34), .S(P1_P1_State2_PTR2), .Z(_02866__PTR2) );
  MUX2_X1 U21707 ( .A(_02865__PTR3), .B(_02865__PTR35), .S(P1_P1_State2_PTR2), .Z(_02866__PTR3) );
  MUX2_X1 U21708 ( .A(_02865__PTR4), .B(_02865__PTR36), .S(P1_P1_State2_PTR2), .Z(_02866__PTR4) );
  MUX2_X1 U21709 ( .A(_02865__PTR5), .B(_02865__PTR37), .S(P1_P1_State2_PTR2), .Z(_02866__PTR5) );
  MUX2_X1 U21710 ( .A(_02865__PTR6), .B(_02865__PTR38), .S(P1_P1_State2_PTR2), .Z(_02866__PTR6) );
  MUX2_X1 U21711 ( .A(_02865__PTR7), .B(_02865__PTR39), .S(P1_P1_State2_PTR2), .Z(_02866__PTR7) );
  MUX2_X1 U21712 ( .A(1'b0), .B(_02864__PTR16), .S(P1_P1_State2_PTR1), .Z(_02865__PTR0) );
  MUX2_X1 U21713 ( .A(1'b0), .B(_02864__PTR17), .S(P1_P1_State2_PTR1), .Z(_02865__PTR1) );
  MUX2_X1 U21714 ( .A(1'b0), .B(_02864__PTR18), .S(P1_P1_State2_PTR1), .Z(_02865__PTR2) );
  MUX2_X1 U21715 ( .A(1'b0), .B(_02864__PTR19), .S(P1_P1_State2_PTR1), .Z(_02865__PTR3) );
  MUX2_X1 U21716 ( .A(1'b0), .B(_02864__PTR20), .S(P1_P1_State2_PTR1), .Z(_02865__PTR4) );
  MUX2_X1 U21717 ( .A(1'b0), .B(_02864__PTR21), .S(P1_P1_State2_PTR1), .Z(_02865__PTR5) );
  MUX2_X1 U21718 ( .A(1'b0), .B(_02864__PTR22), .S(P1_P1_State2_PTR1), .Z(_02865__PTR6) );
  MUX2_X1 U21719 ( .A(1'b0), .B(_02864__PTR23), .S(P1_P1_State2_PTR1), .Z(_02865__PTR7) );
  MUX2_X1 U21720 ( .A(_02864__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02865__PTR32) );
  MUX2_X1 U21721 ( .A(_02864__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02865__PTR33) );
  MUX2_X1 U21722 ( .A(_02864__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02865__PTR34) );
  MUX2_X1 U21723 ( .A(_02864__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02865__PTR35) );
  MUX2_X1 U21724 ( .A(_02864__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02865__PTR36) );
  MUX2_X1 U21725 ( .A(_02864__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02865__PTR37) );
  MUX2_X1 U21726 ( .A(_02864__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02865__PTR38) );
  MUX2_X1 U21727 ( .A(_02864__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02865__PTR39) );
  MUX2_X1 U21728 ( .A(_01898__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR16) );
  MUX2_X1 U21729 ( .A(_01898__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR17) );
  MUX2_X1 U21730 ( .A(_01898__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR18) );
  MUX2_X1 U21731 ( .A(_01898__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR19) );
  MUX2_X1 U21732 ( .A(_01898__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR20) );
  MUX2_X1 U21733 ( .A(_01898__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR21) );
  MUX2_X1 U21734 ( .A(_01898__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR22) );
  MUX2_X1 U21735 ( .A(_01898__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR23) );
  MUX2_X1 U21736 ( .A(_01898__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR32) );
  MUX2_X1 U21737 ( .A(_01898__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR33) );
  MUX2_X1 U21738 ( .A(_01898__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR34) );
  MUX2_X1 U21739 ( .A(_01898__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR35) );
  MUX2_X1 U21740 ( .A(_01898__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR36) );
  MUX2_X1 U21741 ( .A(_01898__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR37) );
  MUX2_X1 U21742 ( .A(_01898__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR38) );
  MUX2_X1 U21743 ( .A(_01898__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR39) );
  MUX2_X1 U21744 ( .A(_01898__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR64) );
  MUX2_X1 U21745 ( .A(_01898__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR65) );
  MUX2_X1 U21746 ( .A(_01898__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR66) );
  MUX2_X1 U21747 ( .A(_01898__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR67) );
  MUX2_X1 U21748 ( .A(_01898__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR68) );
  MUX2_X1 U21749 ( .A(_01898__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR69) );
  MUX2_X1 U21750 ( .A(_01898__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR70) );
  MUX2_X1 U21751 ( .A(_01898__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02864__PTR71) );
  MUX2_X1 U21752 ( .A(_02869__PTR0), .B(_02867__PTR64), .S(P1_P1_State2_PTR3), .Z(_01901__PTR0) );
  MUX2_X1 U21753 ( .A(_02869__PTR1), .B(_02867__PTR65), .S(P1_P1_State2_PTR3), .Z(_01901__PTR1) );
  MUX2_X1 U21754 ( .A(_02869__PTR2), .B(_02867__PTR66), .S(P1_P1_State2_PTR3), .Z(_01901__PTR2) );
  MUX2_X1 U21755 ( .A(_02869__PTR3), .B(_02867__PTR67), .S(P1_P1_State2_PTR3), .Z(_01901__PTR3) );
  MUX2_X1 U21756 ( .A(_02869__PTR4), .B(_02867__PTR68), .S(P1_P1_State2_PTR3), .Z(_01901__PTR4) );
  MUX2_X1 U21757 ( .A(_02869__PTR5), .B(_02867__PTR69), .S(P1_P1_State2_PTR3), .Z(_01901__PTR5) );
  MUX2_X1 U21758 ( .A(_02869__PTR6), .B(_02867__PTR70), .S(P1_P1_State2_PTR3), .Z(_01901__PTR6) );
  MUX2_X1 U21759 ( .A(_02869__PTR7), .B(_02867__PTR71), .S(P1_P1_State2_PTR3), .Z(_01901__PTR7) );
  MUX2_X1 U21760 ( .A(_02868__PTR0), .B(_02868__PTR32), .S(P1_P1_State2_PTR2), .Z(_02869__PTR0) );
  MUX2_X1 U21761 ( .A(_02868__PTR1), .B(_02868__PTR33), .S(P1_P1_State2_PTR2), .Z(_02869__PTR1) );
  MUX2_X1 U21762 ( .A(_02868__PTR2), .B(_02868__PTR34), .S(P1_P1_State2_PTR2), .Z(_02869__PTR2) );
  MUX2_X1 U21763 ( .A(_02868__PTR3), .B(_02868__PTR35), .S(P1_P1_State2_PTR2), .Z(_02869__PTR3) );
  MUX2_X1 U21764 ( .A(_02868__PTR4), .B(_02868__PTR36), .S(P1_P1_State2_PTR2), .Z(_02869__PTR4) );
  MUX2_X1 U21765 ( .A(_02868__PTR5), .B(_02868__PTR37), .S(P1_P1_State2_PTR2), .Z(_02869__PTR5) );
  MUX2_X1 U21766 ( .A(_02868__PTR6), .B(_02868__PTR38), .S(P1_P1_State2_PTR2), .Z(_02869__PTR6) );
  MUX2_X1 U21767 ( .A(_02868__PTR7), .B(_02868__PTR39), .S(P1_P1_State2_PTR2), .Z(_02869__PTR7) );
  MUX2_X1 U21768 ( .A(1'b0), .B(_02867__PTR16), .S(P1_P1_State2_PTR1), .Z(_02868__PTR0) );
  MUX2_X1 U21769 ( .A(1'b0), .B(_02867__PTR17), .S(P1_P1_State2_PTR1), .Z(_02868__PTR1) );
  MUX2_X1 U21770 ( .A(1'b0), .B(_02867__PTR18), .S(P1_P1_State2_PTR1), .Z(_02868__PTR2) );
  MUX2_X1 U21771 ( .A(1'b0), .B(_02867__PTR19), .S(P1_P1_State2_PTR1), .Z(_02868__PTR3) );
  MUX2_X1 U21772 ( .A(1'b0), .B(_02867__PTR20), .S(P1_P1_State2_PTR1), .Z(_02868__PTR4) );
  MUX2_X1 U21773 ( .A(1'b0), .B(_02867__PTR21), .S(P1_P1_State2_PTR1), .Z(_02868__PTR5) );
  MUX2_X1 U21774 ( .A(1'b0), .B(_02867__PTR22), .S(P1_P1_State2_PTR1), .Z(_02868__PTR6) );
  MUX2_X1 U21775 ( .A(1'b0), .B(_02867__PTR23), .S(P1_P1_State2_PTR1), .Z(_02868__PTR7) );
  MUX2_X1 U21776 ( .A(_02867__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02868__PTR32) );
  MUX2_X1 U21777 ( .A(_02867__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02868__PTR33) );
  MUX2_X1 U21778 ( .A(_02867__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02868__PTR34) );
  MUX2_X1 U21779 ( .A(_02867__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02868__PTR35) );
  MUX2_X1 U21780 ( .A(_02867__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02868__PTR36) );
  MUX2_X1 U21781 ( .A(_02867__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02868__PTR37) );
  MUX2_X1 U21782 ( .A(_02867__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02868__PTR38) );
  MUX2_X1 U21783 ( .A(_02867__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02868__PTR39) );
  MUX2_X1 U21784 ( .A(_01900__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR16) );
  MUX2_X1 U21785 ( .A(_01900__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR17) );
  MUX2_X1 U21786 ( .A(_01900__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR18) );
  MUX2_X1 U21787 ( .A(_01900__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR19) );
  MUX2_X1 U21788 ( .A(_01900__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR20) );
  MUX2_X1 U21789 ( .A(_01900__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR21) );
  MUX2_X1 U21790 ( .A(_01900__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR22) );
  MUX2_X1 U21791 ( .A(_01900__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR23) );
  MUX2_X1 U21792 ( .A(_01900__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR32) );
  MUX2_X1 U21793 ( .A(_01900__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR33) );
  MUX2_X1 U21794 ( .A(_01900__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR34) );
  MUX2_X1 U21795 ( .A(_01900__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR35) );
  MUX2_X1 U21796 ( .A(_01900__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR36) );
  MUX2_X1 U21797 ( .A(_01900__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR37) );
  MUX2_X1 U21798 ( .A(_01900__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR38) );
  MUX2_X1 U21799 ( .A(_01900__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR39) );
  MUX2_X1 U21800 ( .A(_01900__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR64) );
  MUX2_X1 U21801 ( .A(_01900__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR65) );
  MUX2_X1 U21802 ( .A(_01900__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR66) );
  MUX2_X1 U21803 ( .A(_01900__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR67) );
  MUX2_X1 U21804 ( .A(_01900__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR68) );
  MUX2_X1 U21805 ( .A(_01900__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR69) );
  MUX2_X1 U21806 ( .A(_01900__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR70) );
  MUX2_X1 U21807 ( .A(_01900__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02867__PTR71) );
  MUX2_X1 U21808 ( .A(_02872__PTR0), .B(_02870__PTR64), .S(P1_P1_State2_PTR3), .Z(_01903__PTR0) );
  MUX2_X1 U21809 ( .A(_02872__PTR1), .B(_02870__PTR65), .S(P1_P1_State2_PTR3), .Z(_01903__PTR1) );
  MUX2_X1 U21810 ( .A(_02872__PTR2), .B(_02870__PTR66), .S(P1_P1_State2_PTR3), .Z(_01903__PTR2) );
  MUX2_X1 U21811 ( .A(_02872__PTR3), .B(_02870__PTR67), .S(P1_P1_State2_PTR3), .Z(_01903__PTR3) );
  MUX2_X1 U21812 ( .A(_02872__PTR4), .B(_02870__PTR68), .S(P1_P1_State2_PTR3), .Z(_01903__PTR4) );
  MUX2_X1 U21813 ( .A(_02872__PTR5), .B(_02870__PTR69), .S(P1_P1_State2_PTR3), .Z(_01903__PTR5) );
  MUX2_X1 U21814 ( .A(_02872__PTR6), .B(_02870__PTR70), .S(P1_P1_State2_PTR3), .Z(_01903__PTR6) );
  MUX2_X1 U21815 ( .A(_02872__PTR7), .B(_02870__PTR71), .S(P1_P1_State2_PTR3), .Z(_01903__PTR7) );
  MUX2_X1 U21816 ( .A(_02871__PTR0), .B(_02871__PTR32), .S(P1_P1_State2_PTR2), .Z(_02872__PTR0) );
  MUX2_X1 U21817 ( .A(_02871__PTR1), .B(_02871__PTR33), .S(P1_P1_State2_PTR2), .Z(_02872__PTR1) );
  MUX2_X1 U21818 ( .A(_02871__PTR2), .B(_02871__PTR34), .S(P1_P1_State2_PTR2), .Z(_02872__PTR2) );
  MUX2_X1 U21819 ( .A(_02871__PTR3), .B(_02871__PTR35), .S(P1_P1_State2_PTR2), .Z(_02872__PTR3) );
  MUX2_X1 U21820 ( .A(_02871__PTR4), .B(_02871__PTR36), .S(P1_P1_State2_PTR2), .Z(_02872__PTR4) );
  MUX2_X1 U21821 ( .A(_02871__PTR5), .B(_02871__PTR37), .S(P1_P1_State2_PTR2), .Z(_02872__PTR5) );
  MUX2_X1 U21822 ( .A(_02871__PTR6), .B(_02871__PTR38), .S(P1_P1_State2_PTR2), .Z(_02872__PTR6) );
  MUX2_X1 U21823 ( .A(_02871__PTR7), .B(_02871__PTR39), .S(P1_P1_State2_PTR2), .Z(_02872__PTR7) );
  MUX2_X1 U21824 ( .A(1'b0), .B(_02870__PTR16), .S(P1_P1_State2_PTR1), .Z(_02871__PTR0) );
  MUX2_X1 U21825 ( .A(1'b0), .B(_02870__PTR17), .S(P1_P1_State2_PTR1), .Z(_02871__PTR1) );
  MUX2_X1 U21826 ( .A(1'b0), .B(_02870__PTR18), .S(P1_P1_State2_PTR1), .Z(_02871__PTR2) );
  MUX2_X1 U21827 ( .A(1'b0), .B(_02870__PTR19), .S(P1_P1_State2_PTR1), .Z(_02871__PTR3) );
  MUX2_X1 U21828 ( .A(1'b0), .B(_02870__PTR20), .S(P1_P1_State2_PTR1), .Z(_02871__PTR4) );
  MUX2_X1 U21829 ( .A(1'b0), .B(_02870__PTR21), .S(P1_P1_State2_PTR1), .Z(_02871__PTR5) );
  MUX2_X1 U21830 ( .A(1'b0), .B(_02870__PTR22), .S(P1_P1_State2_PTR1), .Z(_02871__PTR6) );
  MUX2_X1 U21831 ( .A(1'b0), .B(_02870__PTR23), .S(P1_P1_State2_PTR1), .Z(_02871__PTR7) );
  MUX2_X1 U21832 ( .A(_02870__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02871__PTR32) );
  MUX2_X1 U21833 ( .A(_02870__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02871__PTR33) );
  MUX2_X1 U21834 ( .A(_02870__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02871__PTR34) );
  MUX2_X1 U21835 ( .A(_02870__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02871__PTR35) );
  MUX2_X1 U21836 ( .A(_02870__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02871__PTR36) );
  MUX2_X1 U21837 ( .A(_02870__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02871__PTR37) );
  MUX2_X1 U21838 ( .A(_02870__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02871__PTR38) );
  MUX2_X1 U21839 ( .A(_02870__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02871__PTR39) );
  MUX2_X1 U21840 ( .A(_01902__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR16) );
  MUX2_X1 U21841 ( .A(_01902__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR17) );
  MUX2_X1 U21842 ( .A(_01902__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR18) );
  MUX2_X1 U21843 ( .A(_01902__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR19) );
  MUX2_X1 U21844 ( .A(_01902__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR20) );
  MUX2_X1 U21845 ( .A(_01902__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR21) );
  MUX2_X1 U21846 ( .A(_01902__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR22) );
  MUX2_X1 U21847 ( .A(_01902__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR23) );
  MUX2_X1 U21848 ( .A(_01902__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR32) );
  MUX2_X1 U21849 ( .A(_01902__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR33) );
  MUX2_X1 U21850 ( .A(_01902__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR34) );
  MUX2_X1 U21851 ( .A(_01902__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR35) );
  MUX2_X1 U21852 ( .A(_01902__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR36) );
  MUX2_X1 U21853 ( .A(_01902__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR37) );
  MUX2_X1 U21854 ( .A(_01902__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR38) );
  MUX2_X1 U21855 ( .A(_01902__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR39) );
  MUX2_X1 U21856 ( .A(_01902__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR64) );
  MUX2_X1 U21857 ( .A(_01902__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR65) );
  MUX2_X1 U21858 ( .A(_01902__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR66) );
  MUX2_X1 U21859 ( .A(_01902__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR67) );
  MUX2_X1 U21860 ( .A(_01902__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR68) );
  MUX2_X1 U21861 ( .A(_01902__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR69) );
  MUX2_X1 U21862 ( .A(_01902__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR70) );
  MUX2_X1 U21863 ( .A(_01902__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02870__PTR71) );
  MUX2_X1 U21864 ( .A(_02875__PTR0), .B(_02873__PTR64), .S(P1_P1_State2_PTR3), .Z(_01905__PTR0) );
  MUX2_X1 U21865 ( .A(_02875__PTR1), .B(_02873__PTR65), .S(P1_P1_State2_PTR3), .Z(_01905__PTR1) );
  MUX2_X1 U21866 ( .A(_02875__PTR2), .B(_02873__PTR66), .S(P1_P1_State2_PTR3), .Z(_01905__PTR2) );
  MUX2_X1 U21867 ( .A(_02875__PTR3), .B(_02873__PTR67), .S(P1_P1_State2_PTR3), .Z(_01905__PTR3) );
  MUX2_X1 U21868 ( .A(_02875__PTR4), .B(_02873__PTR68), .S(P1_P1_State2_PTR3), .Z(_01905__PTR4) );
  MUX2_X1 U21869 ( .A(_02875__PTR5), .B(_02873__PTR69), .S(P1_P1_State2_PTR3), .Z(_01905__PTR5) );
  MUX2_X1 U21870 ( .A(_02875__PTR6), .B(_02873__PTR70), .S(P1_P1_State2_PTR3), .Z(_01905__PTR6) );
  MUX2_X1 U21871 ( .A(_02875__PTR7), .B(_02873__PTR71), .S(P1_P1_State2_PTR3), .Z(_01905__PTR7) );
  MUX2_X1 U21872 ( .A(_02874__PTR0), .B(_02874__PTR32), .S(P1_P1_State2_PTR2), .Z(_02875__PTR0) );
  MUX2_X1 U21873 ( .A(_02874__PTR1), .B(_02874__PTR33), .S(P1_P1_State2_PTR2), .Z(_02875__PTR1) );
  MUX2_X1 U21874 ( .A(_02874__PTR2), .B(_02874__PTR34), .S(P1_P1_State2_PTR2), .Z(_02875__PTR2) );
  MUX2_X1 U21875 ( .A(_02874__PTR3), .B(_02874__PTR35), .S(P1_P1_State2_PTR2), .Z(_02875__PTR3) );
  MUX2_X1 U21876 ( .A(_02874__PTR4), .B(_02874__PTR36), .S(P1_P1_State2_PTR2), .Z(_02875__PTR4) );
  MUX2_X1 U21877 ( .A(_02874__PTR5), .B(_02874__PTR37), .S(P1_P1_State2_PTR2), .Z(_02875__PTR5) );
  MUX2_X1 U21878 ( .A(_02874__PTR6), .B(_02874__PTR38), .S(P1_P1_State2_PTR2), .Z(_02875__PTR6) );
  MUX2_X1 U21879 ( .A(_02874__PTR7), .B(_02874__PTR39), .S(P1_P1_State2_PTR2), .Z(_02875__PTR7) );
  MUX2_X1 U21880 ( .A(1'b0), .B(_02873__PTR16), .S(P1_P1_State2_PTR1), .Z(_02874__PTR0) );
  MUX2_X1 U21881 ( .A(1'b0), .B(_02873__PTR17), .S(P1_P1_State2_PTR1), .Z(_02874__PTR1) );
  MUX2_X1 U21882 ( .A(1'b0), .B(_02873__PTR18), .S(P1_P1_State2_PTR1), .Z(_02874__PTR2) );
  MUX2_X1 U21883 ( .A(1'b0), .B(_02873__PTR19), .S(P1_P1_State2_PTR1), .Z(_02874__PTR3) );
  MUX2_X1 U21884 ( .A(1'b0), .B(_02873__PTR20), .S(P1_P1_State2_PTR1), .Z(_02874__PTR4) );
  MUX2_X1 U21885 ( .A(1'b0), .B(_02873__PTR21), .S(P1_P1_State2_PTR1), .Z(_02874__PTR5) );
  MUX2_X1 U21886 ( .A(1'b0), .B(_02873__PTR22), .S(P1_P1_State2_PTR1), .Z(_02874__PTR6) );
  MUX2_X1 U21887 ( .A(1'b0), .B(_02873__PTR23), .S(P1_P1_State2_PTR1), .Z(_02874__PTR7) );
  MUX2_X1 U21888 ( .A(_02873__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02874__PTR32) );
  MUX2_X1 U21889 ( .A(_02873__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02874__PTR33) );
  MUX2_X1 U21890 ( .A(_02873__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02874__PTR34) );
  MUX2_X1 U21891 ( .A(_02873__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02874__PTR35) );
  MUX2_X1 U21892 ( .A(_02873__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02874__PTR36) );
  MUX2_X1 U21893 ( .A(_02873__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02874__PTR37) );
  MUX2_X1 U21894 ( .A(_02873__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02874__PTR38) );
  MUX2_X1 U21895 ( .A(_02873__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02874__PTR39) );
  MUX2_X1 U21896 ( .A(_01904__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR16) );
  MUX2_X1 U21897 ( .A(_01904__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR17) );
  MUX2_X1 U21898 ( .A(_01904__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR18) );
  MUX2_X1 U21899 ( .A(_01904__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR19) );
  MUX2_X1 U21900 ( .A(_01904__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR20) );
  MUX2_X1 U21901 ( .A(_01904__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR21) );
  MUX2_X1 U21902 ( .A(_01904__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR22) );
  MUX2_X1 U21903 ( .A(_01904__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR23) );
  MUX2_X1 U21904 ( .A(_01904__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR32) );
  MUX2_X1 U21905 ( .A(_01904__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR33) );
  MUX2_X1 U21906 ( .A(_01904__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR34) );
  MUX2_X1 U21907 ( .A(_01904__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR35) );
  MUX2_X1 U21908 ( .A(_01904__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR36) );
  MUX2_X1 U21909 ( .A(_01904__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR37) );
  MUX2_X1 U21910 ( .A(_01904__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR38) );
  MUX2_X1 U21911 ( .A(_01904__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR39) );
  MUX2_X1 U21912 ( .A(_01904__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR64) );
  MUX2_X1 U21913 ( .A(_01904__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR65) );
  MUX2_X1 U21914 ( .A(_01904__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR66) );
  MUX2_X1 U21915 ( .A(_01904__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR67) );
  MUX2_X1 U21916 ( .A(_01904__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR68) );
  MUX2_X1 U21917 ( .A(_01904__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR69) );
  MUX2_X1 U21918 ( .A(_01904__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR70) );
  MUX2_X1 U21919 ( .A(_01904__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02873__PTR71) );
  MUX2_X1 U21920 ( .A(_02878__PTR0), .B(_02876__PTR64), .S(P1_P1_State2_PTR3), .Z(_01907__PTR0) );
  MUX2_X1 U21921 ( .A(_02878__PTR1), .B(_02876__PTR65), .S(P1_P1_State2_PTR3), .Z(_01907__PTR1) );
  MUX2_X1 U21922 ( .A(_02878__PTR2), .B(_02876__PTR66), .S(P1_P1_State2_PTR3), .Z(_01907__PTR2) );
  MUX2_X1 U21923 ( .A(_02878__PTR3), .B(_02876__PTR67), .S(P1_P1_State2_PTR3), .Z(_01907__PTR3) );
  MUX2_X1 U21924 ( .A(_02878__PTR4), .B(_02876__PTR68), .S(P1_P1_State2_PTR3), .Z(_01907__PTR4) );
  MUX2_X1 U21925 ( .A(_02878__PTR5), .B(_02876__PTR69), .S(P1_P1_State2_PTR3), .Z(_01907__PTR5) );
  MUX2_X1 U21926 ( .A(_02878__PTR6), .B(_02876__PTR70), .S(P1_P1_State2_PTR3), .Z(_01907__PTR6) );
  MUX2_X1 U21927 ( .A(_02878__PTR7), .B(_02876__PTR71), .S(P1_P1_State2_PTR3), .Z(_01907__PTR7) );
  MUX2_X1 U21928 ( .A(_02877__PTR0), .B(_02877__PTR32), .S(P1_P1_State2_PTR2), .Z(_02878__PTR0) );
  MUX2_X1 U21929 ( .A(_02877__PTR1), .B(_02877__PTR33), .S(P1_P1_State2_PTR2), .Z(_02878__PTR1) );
  MUX2_X1 U21930 ( .A(_02877__PTR2), .B(_02877__PTR34), .S(P1_P1_State2_PTR2), .Z(_02878__PTR2) );
  MUX2_X1 U21931 ( .A(_02877__PTR3), .B(_02877__PTR35), .S(P1_P1_State2_PTR2), .Z(_02878__PTR3) );
  MUX2_X1 U21932 ( .A(_02877__PTR4), .B(_02877__PTR36), .S(P1_P1_State2_PTR2), .Z(_02878__PTR4) );
  MUX2_X1 U21933 ( .A(_02877__PTR5), .B(_02877__PTR37), .S(P1_P1_State2_PTR2), .Z(_02878__PTR5) );
  MUX2_X1 U21934 ( .A(_02877__PTR6), .B(_02877__PTR38), .S(P1_P1_State2_PTR2), .Z(_02878__PTR6) );
  MUX2_X1 U21935 ( .A(_02877__PTR7), .B(_02877__PTR39), .S(P1_P1_State2_PTR2), .Z(_02878__PTR7) );
  MUX2_X1 U21936 ( .A(1'b0), .B(_02876__PTR16), .S(P1_P1_State2_PTR1), .Z(_02877__PTR0) );
  MUX2_X1 U21937 ( .A(1'b0), .B(_02876__PTR17), .S(P1_P1_State2_PTR1), .Z(_02877__PTR1) );
  MUX2_X1 U21938 ( .A(1'b0), .B(_02876__PTR18), .S(P1_P1_State2_PTR1), .Z(_02877__PTR2) );
  MUX2_X1 U21939 ( .A(1'b0), .B(_02876__PTR19), .S(P1_P1_State2_PTR1), .Z(_02877__PTR3) );
  MUX2_X1 U21940 ( .A(1'b0), .B(_02876__PTR20), .S(P1_P1_State2_PTR1), .Z(_02877__PTR4) );
  MUX2_X1 U21941 ( .A(1'b0), .B(_02876__PTR21), .S(P1_P1_State2_PTR1), .Z(_02877__PTR5) );
  MUX2_X1 U21942 ( .A(1'b0), .B(_02876__PTR22), .S(P1_P1_State2_PTR1), .Z(_02877__PTR6) );
  MUX2_X1 U21943 ( .A(1'b0), .B(_02876__PTR23), .S(P1_P1_State2_PTR1), .Z(_02877__PTR7) );
  MUX2_X1 U21944 ( .A(_02876__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02877__PTR32) );
  MUX2_X1 U21945 ( .A(_02876__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02877__PTR33) );
  MUX2_X1 U21946 ( .A(_02876__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02877__PTR34) );
  MUX2_X1 U21947 ( .A(_02876__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02877__PTR35) );
  MUX2_X1 U21948 ( .A(_02876__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02877__PTR36) );
  MUX2_X1 U21949 ( .A(_02876__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02877__PTR37) );
  MUX2_X1 U21950 ( .A(_02876__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02877__PTR38) );
  MUX2_X1 U21951 ( .A(_02876__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02877__PTR39) );
  MUX2_X1 U21952 ( .A(_01906__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR16) );
  MUX2_X1 U21953 ( .A(_01906__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR17) );
  MUX2_X1 U21954 ( .A(_01906__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR18) );
  MUX2_X1 U21955 ( .A(_01906__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR19) );
  MUX2_X1 U21956 ( .A(_01906__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR20) );
  MUX2_X1 U21957 ( .A(_01906__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR21) );
  MUX2_X1 U21958 ( .A(_01906__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR22) );
  MUX2_X1 U21959 ( .A(_01906__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR23) );
  MUX2_X1 U21960 ( .A(_01906__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR32) );
  MUX2_X1 U21961 ( .A(_01906__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR33) );
  MUX2_X1 U21962 ( .A(_01906__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR34) );
  MUX2_X1 U21963 ( .A(_01906__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR35) );
  MUX2_X1 U21964 ( .A(_01906__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR36) );
  MUX2_X1 U21965 ( .A(_01906__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR37) );
  MUX2_X1 U21966 ( .A(_01906__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR38) );
  MUX2_X1 U21967 ( .A(_01906__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR39) );
  MUX2_X1 U21968 ( .A(_01906__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR64) );
  MUX2_X1 U21969 ( .A(_01906__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR65) );
  MUX2_X1 U21970 ( .A(_01906__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR66) );
  MUX2_X1 U21971 ( .A(_01906__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR67) );
  MUX2_X1 U21972 ( .A(_01906__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR68) );
  MUX2_X1 U21973 ( .A(_01906__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR69) );
  MUX2_X1 U21974 ( .A(_01906__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR70) );
  MUX2_X1 U21975 ( .A(_01906__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02876__PTR71) );
  MUX2_X1 U21976 ( .A(_02881__PTR0), .B(_02879__PTR64), .S(P1_P1_State2_PTR3), .Z(_01909__PTR0) );
  MUX2_X1 U21977 ( .A(_02881__PTR1), .B(_02879__PTR65), .S(P1_P1_State2_PTR3), .Z(_01909__PTR1) );
  MUX2_X1 U21978 ( .A(_02881__PTR2), .B(_02879__PTR66), .S(P1_P1_State2_PTR3), .Z(_01909__PTR2) );
  MUX2_X1 U21979 ( .A(_02881__PTR3), .B(_02879__PTR67), .S(P1_P1_State2_PTR3), .Z(_01909__PTR3) );
  MUX2_X1 U21980 ( .A(_02881__PTR4), .B(_02879__PTR68), .S(P1_P1_State2_PTR3), .Z(_01909__PTR4) );
  MUX2_X1 U21981 ( .A(_02881__PTR5), .B(_02879__PTR69), .S(P1_P1_State2_PTR3), .Z(_01909__PTR5) );
  MUX2_X1 U21982 ( .A(_02881__PTR6), .B(_02879__PTR70), .S(P1_P1_State2_PTR3), .Z(_01909__PTR6) );
  MUX2_X1 U21983 ( .A(_02881__PTR7), .B(_02879__PTR71), .S(P1_P1_State2_PTR3), .Z(_01909__PTR7) );
  MUX2_X1 U21984 ( .A(_02880__PTR0), .B(_02880__PTR32), .S(P1_P1_State2_PTR2), .Z(_02881__PTR0) );
  MUX2_X1 U21985 ( .A(_02880__PTR1), .B(_02880__PTR33), .S(P1_P1_State2_PTR2), .Z(_02881__PTR1) );
  MUX2_X1 U21986 ( .A(_02880__PTR2), .B(_02880__PTR34), .S(P1_P1_State2_PTR2), .Z(_02881__PTR2) );
  MUX2_X1 U21987 ( .A(_02880__PTR3), .B(_02880__PTR35), .S(P1_P1_State2_PTR2), .Z(_02881__PTR3) );
  MUX2_X1 U21988 ( .A(_02880__PTR4), .B(_02880__PTR36), .S(P1_P1_State2_PTR2), .Z(_02881__PTR4) );
  MUX2_X1 U21989 ( .A(_02880__PTR5), .B(_02880__PTR37), .S(P1_P1_State2_PTR2), .Z(_02881__PTR5) );
  MUX2_X1 U21990 ( .A(_02880__PTR6), .B(_02880__PTR38), .S(P1_P1_State2_PTR2), .Z(_02881__PTR6) );
  MUX2_X1 U21991 ( .A(_02880__PTR7), .B(_02880__PTR39), .S(P1_P1_State2_PTR2), .Z(_02881__PTR7) );
  MUX2_X1 U21992 ( .A(1'b0), .B(_02879__PTR16), .S(P1_P1_State2_PTR1), .Z(_02880__PTR0) );
  MUX2_X1 U21993 ( .A(1'b0), .B(_02879__PTR17), .S(P1_P1_State2_PTR1), .Z(_02880__PTR1) );
  MUX2_X1 U21994 ( .A(1'b0), .B(_02879__PTR18), .S(P1_P1_State2_PTR1), .Z(_02880__PTR2) );
  MUX2_X1 U21995 ( .A(1'b0), .B(_02879__PTR19), .S(P1_P1_State2_PTR1), .Z(_02880__PTR3) );
  MUX2_X1 U21996 ( .A(1'b0), .B(_02879__PTR20), .S(P1_P1_State2_PTR1), .Z(_02880__PTR4) );
  MUX2_X1 U21997 ( .A(1'b0), .B(_02879__PTR21), .S(P1_P1_State2_PTR1), .Z(_02880__PTR5) );
  MUX2_X1 U21998 ( .A(1'b0), .B(_02879__PTR22), .S(P1_P1_State2_PTR1), .Z(_02880__PTR6) );
  MUX2_X1 U21999 ( .A(1'b0), .B(_02879__PTR23), .S(P1_P1_State2_PTR1), .Z(_02880__PTR7) );
  MUX2_X1 U22000 ( .A(_02879__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02880__PTR32) );
  MUX2_X1 U22001 ( .A(_02879__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02880__PTR33) );
  MUX2_X1 U22002 ( .A(_02879__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02880__PTR34) );
  MUX2_X1 U22003 ( .A(_02879__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02880__PTR35) );
  MUX2_X1 U22004 ( .A(_02879__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02880__PTR36) );
  MUX2_X1 U22005 ( .A(_02879__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02880__PTR37) );
  MUX2_X1 U22006 ( .A(_02879__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02880__PTR38) );
  MUX2_X1 U22007 ( .A(_02879__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02880__PTR39) );
  MUX2_X1 U22008 ( .A(_01908__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR16) );
  MUX2_X1 U22009 ( .A(_01908__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR17) );
  MUX2_X1 U22010 ( .A(_01908__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR18) );
  MUX2_X1 U22011 ( .A(_01908__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR19) );
  MUX2_X1 U22012 ( .A(_01908__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR20) );
  MUX2_X1 U22013 ( .A(_01908__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR21) );
  MUX2_X1 U22014 ( .A(_01908__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR22) );
  MUX2_X1 U22015 ( .A(_01908__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR23) );
  MUX2_X1 U22016 ( .A(_01908__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR32) );
  MUX2_X1 U22017 ( .A(_01908__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR33) );
  MUX2_X1 U22018 ( .A(_01908__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR34) );
  MUX2_X1 U22019 ( .A(_01908__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR35) );
  MUX2_X1 U22020 ( .A(_01908__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR36) );
  MUX2_X1 U22021 ( .A(_01908__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR37) );
  MUX2_X1 U22022 ( .A(_01908__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR38) );
  MUX2_X1 U22023 ( .A(_01908__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR39) );
  MUX2_X1 U22024 ( .A(_01908__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR64) );
  MUX2_X1 U22025 ( .A(_01908__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR65) );
  MUX2_X1 U22026 ( .A(_01908__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR66) );
  MUX2_X1 U22027 ( .A(_01908__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR67) );
  MUX2_X1 U22028 ( .A(_01908__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR68) );
  MUX2_X1 U22029 ( .A(_01908__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR69) );
  MUX2_X1 U22030 ( .A(_01908__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR70) );
  MUX2_X1 U22031 ( .A(_01908__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02879__PTR71) );
  MUX2_X1 U22032 ( .A(_02884__PTR0), .B(_02882__PTR64), .S(P1_P1_State2_PTR3), .Z(_01911__PTR0) );
  MUX2_X1 U22033 ( .A(_02884__PTR1), .B(_02882__PTR65), .S(P1_P1_State2_PTR3), .Z(_01911__PTR1) );
  MUX2_X1 U22034 ( .A(_02884__PTR2), .B(_02882__PTR66), .S(P1_P1_State2_PTR3), .Z(_01911__PTR2) );
  MUX2_X1 U22035 ( .A(_02884__PTR3), .B(_02882__PTR67), .S(P1_P1_State2_PTR3), .Z(_01911__PTR3) );
  MUX2_X1 U22036 ( .A(_02884__PTR4), .B(_02882__PTR68), .S(P1_P1_State2_PTR3), .Z(_01911__PTR4) );
  MUX2_X1 U22037 ( .A(_02884__PTR5), .B(_02882__PTR69), .S(P1_P1_State2_PTR3), .Z(_01911__PTR5) );
  MUX2_X1 U22038 ( .A(_02884__PTR6), .B(_02882__PTR70), .S(P1_P1_State2_PTR3), .Z(_01911__PTR6) );
  MUX2_X1 U22039 ( .A(_02884__PTR7), .B(_02882__PTR71), .S(P1_P1_State2_PTR3), .Z(_01911__PTR7) );
  MUX2_X1 U22040 ( .A(_02883__PTR0), .B(_02883__PTR32), .S(P1_P1_State2_PTR2), .Z(_02884__PTR0) );
  MUX2_X1 U22041 ( .A(_02883__PTR1), .B(_02883__PTR33), .S(P1_P1_State2_PTR2), .Z(_02884__PTR1) );
  MUX2_X1 U22042 ( .A(_02883__PTR2), .B(_02883__PTR34), .S(P1_P1_State2_PTR2), .Z(_02884__PTR2) );
  MUX2_X1 U22043 ( .A(_02883__PTR3), .B(_02883__PTR35), .S(P1_P1_State2_PTR2), .Z(_02884__PTR3) );
  MUX2_X1 U22044 ( .A(_02883__PTR4), .B(_02883__PTR36), .S(P1_P1_State2_PTR2), .Z(_02884__PTR4) );
  MUX2_X1 U22045 ( .A(_02883__PTR5), .B(_02883__PTR37), .S(P1_P1_State2_PTR2), .Z(_02884__PTR5) );
  MUX2_X1 U22046 ( .A(_02883__PTR6), .B(_02883__PTR38), .S(P1_P1_State2_PTR2), .Z(_02884__PTR6) );
  MUX2_X1 U22047 ( .A(_02883__PTR7), .B(_02883__PTR39), .S(P1_P1_State2_PTR2), .Z(_02884__PTR7) );
  MUX2_X1 U22048 ( .A(1'b0), .B(_02882__PTR16), .S(P1_P1_State2_PTR1), .Z(_02883__PTR0) );
  MUX2_X1 U22049 ( .A(1'b0), .B(_02882__PTR17), .S(P1_P1_State2_PTR1), .Z(_02883__PTR1) );
  MUX2_X1 U22050 ( .A(1'b0), .B(_02882__PTR18), .S(P1_P1_State2_PTR1), .Z(_02883__PTR2) );
  MUX2_X1 U22051 ( .A(1'b0), .B(_02882__PTR19), .S(P1_P1_State2_PTR1), .Z(_02883__PTR3) );
  MUX2_X1 U22052 ( .A(1'b0), .B(_02882__PTR20), .S(P1_P1_State2_PTR1), .Z(_02883__PTR4) );
  MUX2_X1 U22053 ( .A(1'b0), .B(_02882__PTR21), .S(P1_P1_State2_PTR1), .Z(_02883__PTR5) );
  MUX2_X1 U22054 ( .A(1'b0), .B(_02882__PTR22), .S(P1_P1_State2_PTR1), .Z(_02883__PTR6) );
  MUX2_X1 U22055 ( .A(1'b0), .B(_02882__PTR23), .S(P1_P1_State2_PTR1), .Z(_02883__PTR7) );
  MUX2_X1 U22056 ( .A(_02882__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02883__PTR32) );
  MUX2_X1 U22057 ( .A(_02882__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02883__PTR33) );
  MUX2_X1 U22058 ( .A(_02882__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02883__PTR34) );
  MUX2_X1 U22059 ( .A(_02882__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02883__PTR35) );
  MUX2_X1 U22060 ( .A(_02882__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02883__PTR36) );
  MUX2_X1 U22061 ( .A(_02882__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02883__PTR37) );
  MUX2_X1 U22062 ( .A(_02882__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02883__PTR38) );
  MUX2_X1 U22063 ( .A(_02882__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02883__PTR39) );
  MUX2_X1 U22064 ( .A(_01910__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR16) );
  MUX2_X1 U22065 ( .A(_01910__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR17) );
  MUX2_X1 U22066 ( .A(_01910__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR18) );
  MUX2_X1 U22067 ( .A(_01910__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR19) );
  MUX2_X1 U22068 ( .A(_01910__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR20) );
  MUX2_X1 U22069 ( .A(_01910__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR21) );
  MUX2_X1 U22070 ( .A(_01910__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR22) );
  MUX2_X1 U22071 ( .A(_01910__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR23) );
  MUX2_X1 U22072 ( .A(_01910__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR32) );
  MUX2_X1 U22073 ( .A(_01910__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR33) );
  MUX2_X1 U22074 ( .A(_01910__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR34) );
  MUX2_X1 U22075 ( .A(_01910__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR35) );
  MUX2_X1 U22076 ( .A(_01910__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR36) );
  MUX2_X1 U22077 ( .A(_01910__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR37) );
  MUX2_X1 U22078 ( .A(_01910__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR38) );
  MUX2_X1 U22079 ( .A(_01910__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR39) );
  MUX2_X1 U22080 ( .A(_01910__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR64) );
  MUX2_X1 U22081 ( .A(_01910__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR65) );
  MUX2_X1 U22082 ( .A(_01910__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR66) );
  MUX2_X1 U22083 ( .A(_01910__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR67) );
  MUX2_X1 U22084 ( .A(_01910__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR68) );
  MUX2_X1 U22085 ( .A(_01910__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR69) );
  MUX2_X1 U22086 ( .A(_01910__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR70) );
  MUX2_X1 U22087 ( .A(_01910__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02882__PTR71) );
  MUX2_X1 U22088 ( .A(_02887__PTR0), .B(_02885__PTR64), .S(P1_P1_State2_PTR3), .Z(_01913__PTR0) );
  MUX2_X1 U22089 ( .A(_02887__PTR1), .B(_02885__PTR65), .S(P1_P1_State2_PTR3), .Z(_01913__PTR1) );
  MUX2_X1 U22090 ( .A(_02887__PTR2), .B(_02885__PTR66), .S(P1_P1_State2_PTR3), .Z(_01913__PTR2) );
  MUX2_X1 U22091 ( .A(_02887__PTR3), .B(_02885__PTR67), .S(P1_P1_State2_PTR3), .Z(_01913__PTR3) );
  MUX2_X1 U22092 ( .A(_02887__PTR4), .B(_02885__PTR68), .S(P1_P1_State2_PTR3), .Z(_01913__PTR4) );
  MUX2_X1 U22093 ( .A(_02887__PTR5), .B(_02885__PTR69), .S(P1_P1_State2_PTR3), .Z(_01913__PTR5) );
  MUX2_X1 U22094 ( .A(_02887__PTR6), .B(_02885__PTR70), .S(P1_P1_State2_PTR3), .Z(_01913__PTR6) );
  MUX2_X1 U22095 ( .A(_02887__PTR7), .B(_02885__PTR71), .S(P1_P1_State2_PTR3), .Z(_01913__PTR7) );
  MUX2_X1 U22096 ( .A(_02886__PTR0), .B(_02886__PTR32), .S(P1_P1_State2_PTR2), .Z(_02887__PTR0) );
  MUX2_X1 U22097 ( .A(_02886__PTR1), .B(_02886__PTR33), .S(P1_P1_State2_PTR2), .Z(_02887__PTR1) );
  MUX2_X1 U22098 ( .A(_02886__PTR2), .B(_02886__PTR34), .S(P1_P1_State2_PTR2), .Z(_02887__PTR2) );
  MUX2_X1 U22099 ( .A(_02886__PTR3), .B(_02886__PTR35), .S(P1_P1_State2_PTR2), .Z(_02887__PTR3) );
  MUX2_X1 U22100 ( .A(_02886__PTR4), .B(_02886__PTR36), .S(P1_P1_State2_PTR2), .Z(_02887__PTR4) );
  MUX2_X1 U22101 ( .A(_02886__PTR5), .B(_02886__PTR37), .S(P1_P1_State2_PTR2), .Z(_02887__PTR5) );
  MUX2_X1 U22102 ( .A(_02886__PTR6), .B(_02886__PTR38), .S(P1_P1_State2_PTR2), .Z(_02887__PTR6) );
  MUX2_X1 U22103 ( .A(_02886__PTR7), .B(_02886__PTR39), .S(P1_P1_State2_PTR2), .Z(_02887__PTR7) );
  MUX2_X1 U22104 ( .A(1'b0), .B(_02885__PTR16), .S(P1_P1_State2_PTR1), .Z(_02886__PTR0) );
  MUX2_X1 U22105 ( .A(1'b0), .B(_02885__PTR17), .S(P1_P1_State2_PTR1), .Z(_02886__PTR1) );
  MUX2_X1 U22106 ( .A(1'b0), .B(_02885__PTR18), .S(P1_P1_State2_PTR1), .Z(_02886__PTR2) );
  MUX2_X1 U22107 ( .A(1'b0), .B(_02885__PTR19), .S(P1_P1_State2_PTR1), .Z(_02886__PTR3) );
  MUX2_X1 U22108 ( .A(1'b0), .B(_02885__PTR20), .S(P1_P1_State2_PTR1), .Z(_02886__PTR4) );
  MUX2_X1 U22109 ( .A(1'b0), .B(_02885__PTR21), .S(P1_P1_State2_PTR1), .Z(_02886__PTR5) );
  MUX2_X1 U22110 ( .A(1'b0), .B(_02885__PTR22), .S(P1_P1_State2_PTR1), .Z(_02886__PTR6) );
  MUX2_X1 U22111 ( .A(1'b0), .B(_02885__PTR23), .S(P1_P1_State2_PTR1), .Z(_02886__PTR7) );
  MUX2_X1 U22112 ( .A(_02885__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02886__PTR32) );
  MUX2_X1 U22113 ( .A(_02885__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02886__PTR33) );
  MUX2_X1 U22114 ( .A(_02885__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02886__PTR34) );
  MUX2_X1 U22115 ( .A(_02885__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02886__PTR35) );
  MUX2_X1 U22116 ( .A(_02885__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02886__PTR36) );
  MUX2_X1 U22117 ( .A(_02885__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02886__PTR37) );
  MUX2_X1 U22118 ( .A(_02885__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02886__PTR38) );
  MUX2_X1 U22119 ( .A(_02885__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02886__PTR39) );
  MUX2_X1 U22120 ( .A(_01912__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR16) );
  MUX2_X1 U22121 ( .A(_01912__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR17) );
  MUX2_X1 U22122 ( .A(_01912__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR18) );
  MUX2_X1 U22123 ( .A(_01912__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR19) );
  MUX2_X1 U22124 ( .A(_01912__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR20) );
  MUX2_X1 U22125 ( .A(_01912__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR21) );
  MUX2_X1 U22126 ( .A(_01912__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR22) );
  MUX2_X1 U22127 ( .A(_01912__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR23) );
  MUX2_X1 U22128 ( .A(_01912__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR32) );
  MUX2_X1 U22129 ( .A(_01912__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR33) );
  MUX2_X1 U22130 ( .A(_01912__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR34) );
  MUX2_X1 U22131 ( .A(_01912__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR35) );
  MUX2_X1 U22132 ( .A(_01912__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR36) );
  MUX2_X1 U22133 ( .A(_01912__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR37) );
  MUX2_X1 U22134 ( .A(_01912__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR38) );
  MUX2_X1 U22135 ( .A(_01912__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR39) );
  MUX2_X1 U22136 ( .A(_01912__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR64) );
  MUX2_X1 U22137 ( .A(_01912__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR65) );
  MUX2_X1 U22138 ( .A(_01912__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR66) );
  MUX2_X1 U22139 ( .A(_01912__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR67) );
  MUX2_X1 U22140 ( .A(_01912__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR68) );
  MUX2_X1 U22141 ( .A(_01912__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR69) );
  MUX2_X1 U22142 ( .A(_01912__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR70) );
  MUX2_X1 U22143 ( .A(_01912__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02885__PTR71) );
  MUX2_X1 U22144 ( .A(_02890__PTR0), .B(_02888__PTR64), .S(P1_P1_State2_PTR3), .Z(_01915__PTR0) );
  MUX2_X1 U22145 ( .A(_02890__PTR1), .B(_02888__PTR65), .S(P1_P1_State2_PTR3), .Z(_01915__PTR1) );
  MUX2_X1 U22146 ( .A(_02890__PTR2), .B(_02888__PTR66), .S(P1_P1_State2_PTR3), .Z(_01915__PTR2) );
  MUX2_X1 U22147 ( .A(_02890__PTR3), .B(_02888__PTR67), .S(P1_P1_State2_PTR3), .Z(_01915__PTR3) );
  MUX2_X1 U22148 ( .A(_02890__PTR4), .B(_02888__PTR68), .S(P1_P1_State2_PTR3), .Z(_01915__PTR4) );
  MUX2_X1 U22149 ( .A(_02890__PTR5), .B(_02888__PTR69), .S(P1_P1_State2_PTR3), .Z(_01915__PTR5) );
  MUX2_X1 U22150 ( .A(_02890__PTR6), .B(_02888__PTR70), .S(P1_P1_State2_PTR3), .Z(_01915__PTR6) );
  MUX2_X1 U22151 ( .A(_02890__PTR7), .B(_02888__PTR71), .S(P1_P1_State2_PTR3), .Z(_01915__PTR7) );
  MUX2_X1 U22152 ( .A(_02889__PTR0), .B(_02889__PTR32), .S(P1_P1_State2_PTR2), .Z(_02890__PTR0) );
  MUX2_X1 U22153 ( .A(_02889__PTR1), .B(_02889__PTR33), .S(P1_P1_State2_PTR2), .Z(_02890__PTR1) );
  MUX2_X1 U22154 ( .A(_02889__PTR2), .B(_02889__PTR34), .S(P1_P1_State2_PTR2), .Z(_02890__PTR2) );
  MUX2_X1 U22155 ( .A(_02889__PTR3), .B(_02889__PTR35), .S(P1_P1_State2_PTR2), .Z(_02890__PTR3) );
  MUX2_X1 U22156 ( .A(_02889__PTR4), .B(_02889__PTR36), .S(P1_P1_State2_PTR2), .Z(_02890__PTR4) );
  MUX2_X1 U22157 ( .A(_02889__PTR5), .B(_02889__PTR37), .S(P1_P1_State2_PTR2), .Z(_02890__PTR5) );
  MUX2_X1 U22158 ( .A(_02889__PTR6), .B(_02889__PTR38), .S(P1_P1_State2_PTR2), .Z(_02890__PTR6) );
  MUX2_X1 U22159 ( .A(_02889__PTR7), .B(_02889__PTR39), .S(P1_P1_State2_PTR2), .Z(_02890__PTR7) );
  MUX2_X1 U22160 ( .A(1'b0), .B(_02888__PTR16), .S(P1_P1_State2_PTR1), .Z(_02889__PTR0) );
  MUX2_X1 U22161 ( .A(1'b0), .B(_02888__PTR17), .S(P1_P1_State2_PTR1), .Z(_02889__PTR1) );
  MUX2_X1 U22162 ( .A(1'b0), .B(_02888__PTR18), .S(P1_P1_State2_PTR1), .Z(_02889__PTR2) );
  MUX2_X1 U22163 ( .A(1'b0), .B(_02888__PTR19), .S(P1_P1_State2_PTR1), .Z(_02889__PTR3) );
  MUX2_X1 U22164 ( .A(1'b0), .B(_02888__PTR20), .S(P1_P1_State2_PTR1), .Z(_02889__PTR4) );
  MUX2_X1 U22165 ( .A(1'b0), .B(_02888__PTR21), .S(P1_P1_State2_PTR1), .Z(_02889__PTR5) );
  MUX2_X1 U22166 ( .A(1'b0), .B(_02888__PTR22), .S(P1_P1_State2_PTR1), .Z(_02889__PTR6) );
  MUX2_X1 U22167 ( .A(1'b0), .B(_02888__PTR23), .S(P1_P1_State2_PTR1), .Z(_02889__PTR7) );
  MUX2_X1 U22168 ( .A(_02888__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02889__PTR32) );
  MUX2_X1 U22169 ( .A(_02888__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02889__PTR33) );
  MUX2_X1 U22170 ( .A(_02888__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02889__PTR34) );
  MUX2_X1 U22171 ( .A(_02888__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02889__PTR35) );
  MUX2_X1 U22172 ( .A(_02888__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02889__PTR36) );
  MUX2_X1 U22173 ( .A(_02888__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02889__PTR37) );
  MUX2_X1 U22174 ( .A(_02888__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02889__PTR38) );
  MUX2_X1 U22175 ( .A(_02888__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02889__PTR39) );
  MUX2_X1 U22176 ( .A(_01914__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR16) );
  MUX2_X1 U22177 ( .A(_01914__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR17) );
  MUX2_X1 U22178 ( .A(_01914__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR18) );
  MUX2_X1 U22179 ( .A(_01914__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR19) );
  MUX2_X1 U22180 ( .A(_01914__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR20) );
  MUX2_X1 U22181 ( .A(_01914__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR21) );
  MUX2_X1 U22182 ( .A(_01914__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR22) );
  MUX2_X1 U22183 ( .A(_01914__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR23) );
  MUX2_X1 U22184 ( .A(_01914__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR32) );
  MUX2_X1 U22185 ( .A(_01914__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR33) );
  MUX2_X1 U22186 ( .A(_01914__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR34) );
  MUX2_X1 U22187 ( .A(_01914__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR35) );
  MUX2_X1 U22188 ( .A(_01914__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR36) );
  MUX2_X1 U22189 ( .A(_01914__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR37) );
  MUX2_X1 U22190 ( .A(_01914__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR38) );
  MUX2_X1 U22191 ( .A(_01914__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR39) );
  MUX2_X1 U22192 ( .A(_01914__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR64) );
  MUX2_X1 U22193 ( .A(_01914__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR65) );
  MUX2_X1 U22194 ( .A(_01914__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR66) );
  MUX2_X1 U22195 ( .A(_01914__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR67) );
  MUX2_X1 U22196 ( .A(_01914__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR68) );
  MUX2_X1 U22197 ( .A(_01914__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR69) );
  MUX2_X1 U22198 ( .A(_01914__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR70) );
  MUX2_X1 U22199 ( .A(_01914__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02888__PTR71) );
  MUX2_X1 U22200 ( .A(_02893__PTR0), .B(_02891__PTR64), .S(P1_P1_State2_PTR3), .Z(_01917__PTR0) );
  MUX2_X1 U22201 ( .A(_02893__PTR1), .B(_02891__PTR65), .S(P1_P1_State2_PTR3), .Z(_01917__PTR1) );
  MUX2_X1 U22202 ( .A(_02893__PTR2), .B(_02891__PTR66), .S(P1_P1_State2_PTR3), .Z(_01917__PTR2) );
  MUX2_X1 U22203 ( .A(_02893__PTR3), .B(_02891__PTR67), .S(P1_P1_State2_PTR3), .Z(_01917__PTR3) );
  MUX2_X1 U22204 ( .A(_02893__PTR4), .B(_02891__PTR68), .S(P1_P1_State2_PTR3), .Z(_01917__PTR4) );
  MUX2_X1 U22205 ( .A(_02893__PTR5), .B(_02891__PTR69), .S(P1_P1_State2_PTR3), .Z(_01917__PTR5) );
  MUX2_X1 U22206 ( .A(_02893__PTR6), .B(_02891__PTR70), .S(P1_P1_State2_PTR3), .Z(_01917__PTR6) );
  MUX2_X1 U22207 ( .A(_02893__PTR7), .B(_02891__PTR71), .S(P1_P1_State2_PTR3), .Z(_01917__PTR7) );
  MUX2_X1 U22208 ( .A(_02892__PTR0), .B(_02892__PTR32), .S(P1_P1_State2_PTR2), .Z(_02893__PTR0) );
  MUX2_X1 U22209 ( .A(_02892__PTR1), .B(_02892__PTR33), .S(P1_P1_State2_PTR2), .Z(_02893__PTR1) );
  MUX2_X1 U22210 ( .A(_02892__PTR2), .B(_02892__PTR34), .S(P1_P1_State2_PTR2), .Z(_02893__PTR2) );
  MUX2_X1 U22211 ( .A(_02892__PTR3), .B(_02892__PTR35), .S(P1_P1_State2_PTR2), .Z(_02893__PTR3) );
  MUX2_X1 U22212 ( .A(_02892__PTR4), .B(_02892__PTR36), .S(P1_P1_State2_PTR2), .Z(_02893__PTR4) );
  MUX2_X1 U22213 ( .A(_02892__PTR5), .B(_02892__PTR37), .S(P1_P1_State2_PTR2), .Z(_02893__PTR5) );
  MUX2_X1 U22214 ( .A(_02892__PTR6), .B(_02892__PTR38), .S(P1_P1_State2_PTR2), .Z(_02893__PTR6) );
  MUX2_X1 U22215 ( .A(_02892__PTR7), .B(_02892__PTR39), .S(P1_P1_State2_PTR2), .Z(_02893__PTR7) );
  MUX2_X1 U22216 ( .A(1'b0), .B(_02891__PTR16), .S(P1_P1_State2_PTR1), .Z(_02892__PTR0) );
  MUX2_X1 U22217 ( .A(1'b0), .B(_02891__PTR17), .S(P1_P1_State2_PTR1), .Z(_02892__PTR1) );
  MUX2_X1 U22218 ( .A(1'b0), .B(_02891__PTR18), .S(P1_P1_State2_PTR1), .Z(_02892__PTR2) );
  MUX2_X1 U22219 ( .A(1'b0), .B(_02891__PTR19), .S(P1_P1_State2_PTR1), .Z(_02892__PTR3) );
  MUX2_X1 U22220 ( .A(1'b0), .B(_02891__PTR20), .S(P1_P1_State2_PTR1), .Z(_02892__PTR4) );
  MUX2_X1 U22221 ( .A(1'b0), .B(_02891__PTR21), .S(P1_P1_State2_PTR1), .Z(_02892__PTR5) );
  MUX2_X1 U22222 ( .A(1'b0), .B(_02891__PTR22), .S(P1_P1_State2_PTR1), .Z(_02892__PTR6) );
  MUX2_X1 U22223 ( .A(1'b0), .B(_02891__PTR23), .S(P1_P1_State2_PTR1), .Z(_02892__PTR7) );
  MUX2_X1 U22224 ( .A(_02891__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02892__PTR32) );
  MUX2_X1 U22225 ( .A(_02891__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02892__PTR33) );
  MUX2_X1 U22226 ( .A(_02891__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02892__PTR34) );
  MUX2_X1 U22227 ( .A(_02891__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02892__PTR35) );
  MUX2_X1 U22228 ( .A(_02891__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02892__PTR36) );
  MUX2_X1 U22229 ( .A(_02891__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02892__PTR37) );
  MUX2_X1 U22230 ( .A(_02891__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02892__PTR38) );
  MUX2_X1 U22231 ( .A(_02891__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02892__PTR39) );
  MUX2_X1 U22232 ( .A(_01916__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR16) );
  MUX2_X1 U22233 ( .A(_01916__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR17) );
  MUX2_X1 U22234 ( .A(_01916__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR18) );
  MUX2_X1 U22235 ( .A(_01916__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR19) );
  MUX2_X1 U22236 ( .A(_01916__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR20) );
  MUX2_X1 U22237 ( .A(_01916__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR21) );
  MUX2_X1 U22238 ( .A(_01916__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR22) );
  MUX2_X1 U22239 ( .A(_01916__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR23) );
  MUX2_X1 U22240 ( .A(_01916__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR32) );
  MUX2_X1 U22241 ( .A(_01916__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR33) );
  MUX2_X1 U22242 ( .A(_01916__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR34) );
  MUX2_X1 U22243 ( .A(_01916__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR35) );
  MUX2_X1 U22244 ( .A(_01916__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR36) );
  MUX2_X1 U22245 ( .A(_01916__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR37) );
  MUX2_X1 U22246 ( .A(_01916__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR38) );
  MUX2_X1 U22247 ( .A(_01916__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR39) );
  MUX2_X1 U22248 ( .A(_01916__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR64) );
  MUX2_X1 U22249 ( .A(_01916__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR65) );
  MUX2_X1 U22250 ( .A(_01916__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR66) );
  MUX2_X1 U22251 ( .A(_01916__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR67) );
  MUX2_X1 U22252 ( .A(_01916__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR68) );
  MUX2_X1 U22253 ( .A(_01916__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR69) );
  MUX2_X1 U22254 ( .A(_01916__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR70) );
  MUX2_X1 U22255 ( .A(_01916__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02891__PTR71) );
  MUX2_X1 U22256 ( .A(_02896__PTR0), .B(_02894__PTR64), .S(P1_P1_State2_PTR3), .Z(_01919__PTR0) );
  MUX2_X1 U22257 ( .A(_02896__PTR1), .B(_02894__PTR65), .S(P1_P1_State2_PTR3), .Z(_01919__PTR1) );
  MUX2_X1 U22258 ( .A(_02896__PTR2), .B(_02894__PTR66), .S(P1_P1_State2_PTR3), .Z(_01919__PTR2) );
  MUX2_X1 U22259 ( .A(_02896__PTR3), .B(_02894__PTR67), .S(P1_P1_State2_PTR3), .Z(_01919__PTR3) );
  MUX2_X1 U22260 ( .A(_02896__PTR4), .B(_02894__PTR68), .S(P1_P1_State2_PTR3), .Z(_01919__PTR4) );
  MUX2_X1 U22261 ( .A(_02896__PTR5), .B(_02894__PTR69), .S(P1_P1_State2_PTR3), .Z(_01919__PTR5) );
  MUX2_X1 U22262 ( .A(_02896__PTR6), .B(_02894__PTR70), .S(P1_P1_State2_PTR3), .Z(_01919__PTR6) );
  MUX2_X1 U22263 ( .A(_02896__PTR7), .B(_02894__PTR71), .S(P1_P1_State2_PTR3), .Z(_01919__PTR7) );
  MUX2_X1 U22264 ( .A(_02895__PTR0), .B(_02895__PTR32), .S(P1_P1_State2_PTR2), .Z(_02896__PTR0) );
  MUX2_X1 U22265 ( .A(_02895__PTR1), .B(_02895__PTR33), .S(P1_P1_State2_PTR2), .Z(_02896__PTR1) );
  MUX2_X1 U22266 ( .A(_02895__PTR2), .B(_02895__PTR34), .S(P1_P1_State2_PTR2), .Z(_02896__PTR2) );
  MUX2_X1 U22267 ( .A(_02895__PTR3), .B(_02895__PTR35), .S(P1_P1_State2_PTR2), .Z(_02896__PTR3) );
  MUX2_X1 U22268 ( .A(_02895__PTR4), .B(_02895__PTR36), .S(P1_P1_State2_PTR2), .Z(_02896__PTR4) );
  MUX2_X1 U22269 ( .A(_02895__PTR5), .B(_02895__PTR37), .S(P1_P1_State2_PTR2), .Z(_02896__PTR5) );
  MUX2_X1 U22270 ( .A(_02895__PTR6), .B(_02895__PTR38), .S(P1_P1_State2_PTR2), .Z(_02896__PTR6) );
  MUX2_X1 U22271 ( .A(_02895__PTR7), .B(_02895__PTR39), .S(P1_P1_State2_PTR2), .Z(_02896__PTR7) );
  MUX2_X1 U22272 ( .A(1'b0), .B(_02894__PTR16), .S(P1_P1_State2_PTR1), .Z(_02895__PTR0) );
  MUX2_X1 U22273 ( .A(1'b0), .B(_02894__PTR17), .S(P1_P1_State2_PTR1), .Z(_02895__PTR1) );
  MUX2_X1 U22274 ( .A(1'b0), .B(_02894__PTR18), .S(P1_P1_State2_PTR1), .Z(_02895__PTR2) );
  MUX2_X1 U22275 ( .A(1'b0), .B(_02894__PTR19), .S(P1_P1_State2_PTR1), .Z(_02895__PTR3) );
  MUX2_X1 U22276 ( .A(1'b0), .B(_02894__PTR20), .S(P1_P1_State2_PTR1), .Z(_02895__PTR4) );
  MUX2_X1 U22277 ( .A(1'b0), .B(_02894__PTR21), .S(P1_P1_State2_PTR1), .Z(_02895__PTR5) );
  MUX2_X1 U22278 ( .A(1'b0), .B(_02894__PTR22), .S(P1_P1_State2_PTR1), .Z(_02895__PTR6) );
  MUX2_X1 U22279 ( .A(1'b0), .B(_02894__PTR23), .S(P1_P1_State2_PTR1), .Z(_02895__PTR7) );
  MUX2_X1 U22280 ( .A(_02894__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02895__PTR32) );
  MUX2_X1 U22281 ( .A(_02894__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02895__PTR33) );
  MUX2_X1 U22282 ( .A(_02894__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02895__PTR34) );
  MUX2_X1 U22283 ( .A(_02894__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02895__PTR35) );
  MUX2_X1 U22284 ( .A(_02894__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02895__PTR36) );
  MUX2_X1 U22285 ( .A(_02894__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02895__PTR37) );
  MUX2_X1 U22286 ( .A(_02894__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02895__PTR38) );
  MUX2_X1 U22287 ( .A(_02894__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02895__PTR39) );
  MUX2_X1 U22288 ( .A(_01918__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR16) );
  MUX2_X1 U22289 ( .A(_01918__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR17) );
  MUX2_X1 U22290 ( .A(_01918__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR18) );
  MUX2_X1 U22291 ( .A(_01918__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR19) );
  MUX2_X1 U22292 ( .A(_01918__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR20) );
  MUX2_X1 U22293 ( .A(_01918__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR21) );
  MUX2_X1 U22294 ( .A(_01918__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR22) );
  MUX2_X1 U22295 ( .A(_01918__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR23) );
  MUX2_X1 U22296 ( .A(_01918__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR32) );
  MUX2_X1 U22297 ( .A(_01918__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR33) );
  MUX2_X1 U22298 ( .A(_01918__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR34) );
  MUX2_X1 U22299 ( .A(_01918__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR35) );
  MUX2_X1 U22300 ( .A(_01918__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR36) );
  MUX2_X1 U22301 ( .A(_01918__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR37) );
  MUX2_X1 U22302 ( .A(_01918__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR38) );
  MUX2_X1 U22303 ( .A(_01918__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR39) );
  MUX2_X1 U22304 ( .A(_01918__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR64) );
  MUX2_X1 U22305 ( .A(_01918__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR65) );
  MUX2_X1 U22306 ( .A(_01918__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR66) );
  MUX2_X1 U22307 ( .A(_01918__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR67) );
  MUX2_X1 U22308 ( .A(_01918__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR68) );
  MUX2_X1 U22309 ( .A(_01918__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR69) );
  MUX2_X1 U22310 ( .A(_01918__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR70) );
  MUX2_X1 U22311 ( .A(_01918__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02894__PTR71) );
  MUX2_X1 U22312 ( .A(_02899__PTR0), .B(_02897__PTR64), .S(P1_P1_State2_PTR3), .Z(_01921__PTR0) );
  MUX2_X1 U22313 ( .A(_02899__PTR1), .B(_02897__PTR65), .S(P1_P1_State2_PTR3), .Z(_01921__PTR1) );
  MUX2_X1 U22314 ( .A(_02899__PTR2), .B(_02897__PTR66), .S(P1_P1_State2_PTR3), .Z(_01921__PTR2) );
  MUX2_X1 U22315 ( .A(_02899__PTR3), .B(_02897__PTR67), .S(P1_P1_State2_PTR3), .Z(_01921__PTR3) );
  MUX2_X1 U22316 ( .A(_02899__PTR4), .B(_02897__PTR68), .S(P1_P1_State2_PTR3), .Z(_01921__PTR4) );
  MUX2_X1 U22317 ( .A(_02899__PTR5), .B(_02897__PTR69), .S(P1_P1_State2_PTR3), .Z(_01921__PTR5) );
  MUX2_X1 U22318 ( .A(_02899__PTR6), .B(_02897__PTR70), .S(P1_P1_State2_PTR3), .Z(_01921__PTR6) );
  MUX2_X1 U22319 ( .A(_02899__PTR7), .B(_02897__PTR71), .S(P1_P1_State2_PTR3), .Z(_01921__PTR7) );
  MUX2_X1 U22320 ( .A(_02898__PTR0), .B(_02898__PTR32), .S(P1_P1_State2_PTR2), .Z(_02899__PTR0) );
  MUX2_X1 U22321 ( .A(_02898__PTR1), .B(_02898__PTR33), .S(P1_P1_State2_PTR2), .Z(_02899__PTR1) );
  MUX2_X1 U22322 ( .A(_02898__PTR2), .B(_02898__PTR34), .S(P1_P1_State2_PTR2), .Z(_02899__PTR2) );
  MUX2_X1 U22323 ( .A(_02898__PTR3), .B(_02898__PTR35), .S(P1_P1_State2_PTR2), .Z(_02899__PTR3) );
  MUX2_X1 U22324 ( .A(_02898__PTR4), .B(_02898__PTR36), .S(P1_P1_State2_PTR2), .Z(_02899__PTR4) );
  MUX2_X1 U22325 ( .A(_02898__PTR5), .B(_02898__PTR37), .S(P1_P1_State2_PTR2), .Z(_02899__PTR5) );
  MUX2_X1 U22326 ( .A(_02898__PTR6), .B(_02898__PTR38), .S(P1_P1_State2_PTR2), .Z(_02899__PTR6) );
  MUX2_X1 U22327 ( .A(_02898__PTR7), .B(_02898__PTR39), .S(P1_P1_State2_PTR2), .Z(_02899__PTR7) );
  MUX2_X1 U22328 ( .A(1'b0), .B(_02897__PTR16), .S(P1_P1_State2_PTR1), .Z(_02898__PTR0) );
  MUX2_X1 U22329 ( .A(1'b0), .B(_02897__PTR17), .S(P1_P1_State2_PTR1), .Z(_02898__PTR1) );
  MUX2_X1 U22330 ( .A(1'b0), .B(_02897__PTR18), .S(P1_P1_State2_PTR1), .Z(_02898__PTR2) );
  MUX2_X1 U22331 ( .A(1'b0), .B(_02897__PTR19), .S(P1_P1_State2_PTR1), .Z(_02898__PTR3) );
  MUX2_X1 U22332 ( .A(1'b0), .B(_02897__PTR20), .S(P1_P1_State2_PTR1), .Z(_02898__PTR4) );
  MUX2_X1 U22333 ( .A(1'b0), .B(_02897__PTR21), .S(P1_P1_State2_PTR1), .Z(_02898__PTR5) );
  MUX2_X1 U22334 ( .A(1'b0), .B(_02897__PTR22), .S(P1_P1_State2_PTR1), .Z(_02898__PTR6) );
  MUX2_X1 U22335 ( .A(1'b0), .B(_02897__PTR23), .S(P1_P1_State2_PTR1), .Z(_02898__PTR7) );
  MUX2_X1 U22336 ( .A(_02897__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02898__PTR32) );
  MUX2_X1 U22337 ( .A(_02897__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02898__PTR33) );
  MUX2_X1 U22338 ( .A(_02897__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02898__PTR34) );
  MUX2_X1 U22339 ( .A(_02897__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02898__PTR35) );
  MUX2_X1 U22340 ( .A(_02897__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02898__PTR36) );
  MUX2_X1 U22341 ( .A(_02897__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02898__PTR37) );
  MUX2_X1 U22342 ( .A(_02897__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02898__PTR38) );
  MUX2_X1 U22343 ( .A(_02897__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02898__PTR39) );
  MUX2_X1 U22344 ( .A(_01920__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR16) );
  MUX2_X1 U22345 ( .A(_01920__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR17) );
  MUX2_X1 U22346 ( .A(_01920__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR18) );
  MUX2_X1 U22347 ( .A(_01920__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR19) );
  MUX2_X1 U22348 ( .A(_01920__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR20) );
  MUX2_X1 U22349 ( .A(_01920__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR21) );
  MUX2_X1 U22350 ( .A(_01920__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR22) );
  MUX2_X1 U22351 ( .A(_01920__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR23) );
  MUX2_X1 U22352 ( .A(_01920__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR32) );
  MUX2_X1 U22353 ( .A(_01920__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR33) );
  MUX2_X1 U22354 ( .A(_01920__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR34) );
  MUX2_X1 U22355 ( .A(_01920__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR35) );
  MUX2_X1 U22356 ( .A(_01920__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR36) );
  MUX2_X1 U22357 ( .A(_01920__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR37) );
  MUX2_X1 U22358 ( .A(_01920__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR38) );
  MUX2_X1 U22359 ( .A(_01920__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR39) );
  MUX2_X1 U22360 ( .A(_01920__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR64) );
  MUX2_X1 U22361 ( .A(_01920__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR65) );
  MUX2_X1 U22362 ( .A(_01920__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR66) );
  MUX2_X1 U22363 ( .A(_01920__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR67) );
  MUX2_X1 U22364 ( .A(_01920__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR68) );
  MUX2_X1 U22365 ( .A(_01920__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR69) );
  MUX2_X1 U22366 ( .A(_01920__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR70) );
  MUX2_X1 U22367 ( .A(_01920__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02897__PTR71) );
  MUX2_X1 U22368 ( .A(_02902__PTR0), .B(_02900__PTR64), .S(P1_P1_State2_PTR3), .Z(_01923__PTR0) );
  MUX2_X1 U22369 ( .A(_02902__PTR1), .B(_02900__PTR65), .S(P1_P1_State2_PTR3), .Z(_01923__PTR1) );
  MUX2_X1 U22370 ( .A(_02902__PTR2), .B(_02900__PTR66), .S(P1_P1_State2_PTR3), .Z(_01923__PTR2) );
  MUX2_X1 U22371 ( .A(_02902__PTR3), .B(_02900__PTR67), .S(P1_P1_State2_PTR3), .Z(_01923__PTR3) );
  MUX2_X1 U22372 ( .A(_02902__PTR4), .B(_02900__PTR68), .S(P1_P1_State2_PTR3), .Z(_01923__PTR4) );
  MUX2_X1 U22373 ( .A(_02902__PTR5), .B(_02900__PTR69), .S(P1_P1_State2_PTR3), .Z(_01923__PTR5) );
  MUX2_X1 U22374 ( .A(_02902__PTR6), .B(_02900__PTR70), .S(P1_P1_State2_PTR3), .Z(_01923__PTR6) );
  MUX2_X1 U22375 ( .A(_02902__PTR7), .B(_02900__PTR71), .S(P1_P1_State2_PTR3), .Z(_01923__PTR7) );
  MUX2_X1 U22376 ( .A(_02901__PTR0), .B(_02901__PTR32), .S(P1_P1_State2_PTR2), .Z(_02902__PTR0) );
  MUX2_X1 U22377 ( .A(_02901__PTR1), .B(_02901__PTR33), .S(P1_P1_State2_PTR2), .Z(_02902__PTR1) );
  MUX2_X1 U22378 ( .A(_02901__PTR2), .B(_02901__PTR34), .S(P1_P1_State2_PTR2), .Z(_02902__PTR2) );
  MUX2_X1 U22379 ( .A(_02901__PTR3), .B(_02901__PTR35), .S(P1_P1_State2_PTR2), .Z(_02902__PTR3) );
  MUX2_X1 U22380 ( .A(_02901__PTR4), .B(_02901__PTR36), .S(P1_P1_State2_PTR2), .Z(_02902__PTR4) );
  MUX2_X1 U22381 ( .A(_02901__PTR5), .B(_02901__PTR37), .S(P1_P1_State2_PTR2), .Z(_02902__PTR5) );
  MUX2_X1 U22382 ( .A(_02901__PTR6), .B(_02901__PTR38), .S(P1_P1_State2_PTR2), .Z(_02902__PTR6) );
  MUX2_X1 U22383 ( .A(_02901__PTR7), .B(_02901__PTR39), .S(P1_P1_State2_PTR2), .Z(_02902__PTR7) );
  MUX2_X1 U22384 ( .A(1'b0), .B(_02900__PTR16), .S(P1_P1_State2_PTR1), .Z(_02901__PTR0) );
  MUX2_X1 U22385 ( .A(1'b0), .B(_02900__PTR17), .S(P1_P1_State2_PTR1), .Z(_02901__PTR1) );
  MUX2_X1 U22386 ( .A(1'b0), .B(_02900__PTR18), .S(P1_P1_State2_PTR1), .Z(_02901__PTR2) );
  MUX2_X1 U22387 ( .A(1'b0), .B(_02900__PTR19), .S(P1_P1_State2_PTR1), .Z(_02901__PTR3) );
  MUX2_X1 U22388 ( .A(1'b0), .B(_02900__PTR20), .S(P1_P1_State2_PTR1), .Z(_02901__PTR4) );
  MUX2_X1 U22389 ( .A(1'b0), .B(_02900__PTR21), .S(P1_P1_State2_PTR1), .Z(_02901__PTR5) );
  MUX2_X1 U22390 ( .A(1'b0), .B(_02900__PTR22), .S(P1_P1_State2_PTR1), .Z(_02901__PTR6) );
  MUX2_X1 U22391 ( .A(1'b0), .B(_02900__PTR23), .S(P1_P1_State2_PTR1), .Z(_02901__PTR7) );
  MUX2_X1 U22392 ( .A(_02900__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02901__PTR32) );
  MUX2_X1 U22393 ( .A(_02900__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02901__PTR33) );
  MUX2_X1 U22394 ( .A(_02900__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02901__PTR34) );
  MUX2_X1 U22395 ( .A(_02900__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02901__PTR35) );
  MUX2_X1 U22396 ( .A(_02900__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02901__PTR36) );
  MUX2_X1 U22397 ( .A(_02900__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02901__PTR37) );
  MUX2_X1 U22398 ( .A(_02900__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02901__PTR38) );
  MUX2_X1 U22399 ( .A(_02900__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02901__PTR39) );
  MUX2_X1 U22400 ( .A(_01922__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR16) );
  MUX2_X1 U22401 ( .A(_01922__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR17) );
  MUX2_X1 U22402 ( .A(_01922__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR18) );
  MUX2_X1 U22403 ( .A(_01922__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR19) );
  MUX2_X1 U22404 ( .A(_01922__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR20) );
  MUX2_X1 U22405 ( .A(_01922__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR21) );
  MUX2_X1 U22406 ( .A(_01922__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR22) );
  MUX2_X1 U22407 ( .A(_01922__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR23) );
  MUX2_X1 U22408 ( .A(_01922__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR32) );
  MUX2_X1 U22409 ( .A(_01922__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR33) );
  MUX2_X1 U22410 ( .A(_01922__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR34) );
  MUX2_X1 U22411 ( .A(_01922__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR35) );
  MUX2_X1 U22412 ( .A(_01922__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR36) );
  MUX2_X1 U22413 ( .A(_01922__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR37) );
  MUX2_X1 U22414 ( .A(_01922__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR38) );
  MUX2_X1 U22415 ( .A(_01922__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR39) );
  MUX2_X1 U22416 ( .A(_01922__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR64) );
  MUX2_X1 U22417 ( .A(_01922__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR65) );
  MUX2_X1 U22418 ( .A(_01922__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR66) );
  MUX2_X1 U22419 ( .A(_01922__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR67) );
  MUX2_X1 U22420 ( .A(_01922__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR68) );
  MUX2_X1 U22421 ( .A(_01922__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR69) );
  MUX2_X1 U22422 ( .A(_01922__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR70) );
  MUX2_X1 U22423 ( .A(_01922__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02900__PTR71) );
  MUX2_X1 U22424 ( .A(_02905__PTR0), .B(_02903__PTR64), .S(P1_P1_State2_PTR3), .Z(_01925__PTR0) );
  MUX2_X1 U22425 ( .A(_02905__PTR1), .B(_02903__PTR65), .S(P1_P1_State2_PTR3), .Z(_01925__PTR1) );
  MUX2_X1 U22426 ( .A(_02905__PTR2), .B(_02903__PTR66), .S(P1_P1_State2_PTR3), .Z(_01925__PTR2) );
  MUX2_X1 U22427 ( .A(_02905__PTR3), .B(_02903__PTR67), .S(P1_P1_State2_PTR3), .Z(_01925__PTR3) );
  MUX2_X1 U22428 ( .A(_02905__PTR4), .B(_02903__PTR68), .S(P1_P1_State2_PTR3), .Z(_01925__PTR4) );
  MUX2_X1 U22429 ( .A(_02905__PTR5), .B(_02903__PTR69), .S(P1_P1_State2_PTR3), .Z(_01925__PTR5) );
  MUX2_X1 U22430 ( .A(_02905__PTR6), .B(_02903__PTR70), .S(P1_P1_State2_PTR3), .Z(_01925__PTR6) );
  MUX2_X1 U22431 ( .A(_02905__PTR7), .B(_02903__PTR71), .S(P1_P1_State2_PTR3), .Z(_01925__PTR7) );
  MUX2_X1 U22432 ( .A(_02904__PTR0), .B(_02904__PTR32), .S(P1_P1_State2_PTR2), .Z(_02905__PTR0) );
  MUX2_X1 U22433 ( .A(_02904__PTR1), .B(_02904__PTR33), .S(P1_P1_State2_PTR2), .Z(_02905__PTR1) );
  MUX2_X1 U22434 ( .A(_02904__PTR2), .B(_02904__PTR34), .S(P1_P1_State2_PTR2), .Z(_02905__PTR2) );
  MUX2_X1 U22435 ( .A(_02904__PTR3), .B(_02904__PTR35), .S(P1_P1_State2_PTR2), .Z(_02905__PTR3) );
  MUX2_X1 U22436 ( .A(_02904__PTR4), .B(_02904__PTR36), .S(P1_P1_State2_PTR2), .Z(_02905__PTR4) );
  MUX2_X1 U22437 ( .A(_02904__PTR5), .B(_02904__PTR37), .S(P1_P1_State2_PTR2), .Z(_02905__PTR5) );
  MUX2_X1 U22438 ( .A(_02904__PTR6), .B(_02904__PTR38), .S(P1_P1_State2_PTR2), .Z(_02905__PTR6) );
  MUX2_X1 U22439 ( .A(_02904__PTR7), .B(_02904__PTR39), .S(P1_P1_State2_PTR2), .Z(_02905__PTR7) );
  MUX2_X1 U22440 ( .A(1'b0), .B(_02903__PTR16), .S(P1_P1_State2_PTR1), .Z(_02904__PTR0) );
  MUX2_X1 U22441 ( .A(1'b0), .B(_02903__PTR17), .S(P1_P1_State2_PTR1), .Z(_02904__PTR1) );
  MUX2_X1 U22442 ( .A(1'b0), .B(_02903__PTR18), .S(P1_P1_State2_PTR1), .Z(_02904__PTR2) );
  MUX2_X1 U22443 ( .A(1'b0), .B(_02903__PTR19), .S(P1_P1_State2_PTR1), .Z(_02904__PTR3) );
  MUX2_X1 U22444 ( .A(1'b0), .B(_02903__PTR20), .S(P1_P1_State2_PTR1), .Z(_02904__PTR4) );
  MUX2_X1 U22445 ( .A(1'b0), .B(_02903__PTR21), .S(P1_P1_State2_PTR1), .Z(_02904__PTR5) );
  MUX2_X1 U22446 ( .A(1'b0), .B(_02903__PTR22), .S(P1_P1_State2_PTR1), .Z(_02904__PTR6) );
  MUX2_X1 U22447 ( .A(1'b0), .B(_02903__PTR23), .S(P1_P1_State2_PTR1), .Z(_02904__PTR7) );
  MUX2_X1 U22448 ( .A(_02903__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02904__PTR32) );
  MUX2_X1 U22449 ( .A(_02903__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02904__PTR33) );
  MUX2_X1 U22450 ( .A(_02903__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02904__PTR34) );
  MUX2_X1 U22451 ( .A(_02903__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02904__PTR35) );
  MUX2_X1 U22452 ( .A(_02903__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02904__PTR36) );
  MUX2_X1 U22453 ( .A(_02903__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02904__PTR37) );
  MUX2_X1 U22454 ( .A(_02903__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02904__PTR38) );
  MUX2_X1 U22455 ( .A(_02903__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02904__PTR39) );
  MUX2_X1 U22456 ( .A(_01924__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR16) );
  MUX2_X1 U22457 ( .A(_01924__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR17) );
  MUX2_X1 U22458 ( .A(_01924__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR18) );
  MUX2_X1 U22459 ( .A(_01924__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR19) );
  MUX2_X1 U22460 ( .A(_01924__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR20) );
  MUX2_X1 U22461 ( .A(_01924__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR21) );
  MUX2_X1 U22462 ( .A(_01924__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR22) );
  MUX2_X1 U22463 ( .A(_01924__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR23) );
  MUX2_X1 U22464 ( .A(_01924__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR32) );
  MUX2_X1 U22465 ( .A(_01924__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR33) );
  MUX2_X1 U22466 ( .A(_01924__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR34) );
  MUX2_X1 U22467 ( .A(_01924__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR35) );
  MUX2_X1 U22468 ( .A(_01924__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR36) );
  MUX2_X1 U22469 ( .A(_01924__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR37) );
  MUX2_X1 U22470 ( .A(_01924__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR38) );
  MUX2_X1 U22471 ( .A(_01924__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR39) );
  MUX2_X1 U22472 ( .A(_01924__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR64) );
  MUX2_X1 U22473 ( .A(_01924__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR65) );
  MUX2_X1 U22474 ( .A(_01924__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR66) );
  MUX2_X1 U22475 ( .A(_01924__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR67) );
  MUX2_X1 U22476 ( .A(_01924__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR68) );
  MUX2_X1 U22477 ( .A(_01924__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR69) );
  MUX2_X1 U22478 ( .A(_01924__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR70) );
  MUX2_X1 U22479 ( .A(_01924__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02903__PTR71) );
  MUX2_X1 U22480 ( .A(_02908__PTR0), .B(_02906__PTR64), .S(P1_P1_State2_PTR3), .Z(_01927__PTR0) );
  MUX2_X1 U22481 ( .A(_02908__PTR1), .B(_02906__PTR65), .S(P1_P1_State2_PTR3), .Z(_01927__PTR1) );
  MUX2_X1 U22482 ( .A(_02908__PTR2), .B(_02906__PTR66), .S(P1_P1_State2_PTR3), .Z(_01927__PTR2) );
  MUX2_X1 U22483 ( .A(_02908__PTR3), .B(_02906__PTR67), .S(P1_P1_State2_PTR3), .Z(_01927__PTR3) );
  MUX2_X1 U22484 ( .A(_02908__PTR4), .B(_02906__PTR68), .S(P1_P1_State2_PTR3), .Z(_01927__PTR4) );
  MUX2_X1 U22485 ( .A(_02908__PTR5), .B(_02906__PTR69), .S(P1_P1_State2_PTR3), .Z(_01927__PTR5) );
  MUX2_X1 U22486 ( .A(_02908__PTR6), .B(_02906__PTR70), .S(P1_P1_State2_PTR3), .Z(_01927__PTR6) );
  MUX2_X1 U22487 ( .A(_02908__PTR7), .B(_02906__PTR71), .S(P1_P1_State2_PTR3), .Z(_01927__PTR7) );
  MUX2_X1 U22488 ( .A(_02907__PTR0), .B(_02907__PTR32), .S(P1_P1_State2_PTR2), .Z(_02908__PTR0) );
  MUX2_X1 U22489 ( .A(_02907__PTR1), .B(_02907__PTR33), .S(P1_P1_State2_PTR2), .Z(_02908__PTR1) );
  MUX2_X1 U22490 ( .A(_02907__PTR2), .B(_02907__PTR34), .S(P1_P1_State2_PTR2), .Z(_02908__PTR2) );
  MUX2_X1 U22491 ( .A(_02907__PTR3), .B(_02907__PTR35), .S(P1_P1_State2_PTR2), .Z(_02908__PTR3) );
  MUX2_X1 U22492 ( .A(_02907__PTR4), .B(_02907__PTR36), .S(P1_P1_State2_PTR2), .Z(_02908__PTR4) );
  MUX2_X1 U22493 ( .A(_02907__PTR5), .B(_02907__PTR37), .S(P1_P1_State2_PTR2), .Z(_02908__PTR5) );
  MUX2_X1 U22494 ( .A(_02907__PTR6), .B(_02907__PTR38), .S(P1_P1_State2_PTR2), .Z(_02908__PTR6) );
  MUX2_X1 U22495 ( .A(_02907__PTR7), .B(_02907__PTR39), .S(P1_P1_State2_PTR2), .Z(_02908__PTR7) );
  MUX2_X1 U22496 ( .A(1'b0), .B(_02906__PTR16), .S(P1_P1_State2_PTR1), .Z(_02907__PTR0) );
  MUX2_X1 U22497 ( .A(1'b0), .B(_02906__PTR17), .S(P1_P1_State2_PTR1), .Z(_02907__PTR1) );
  MUX2_X1 U22498 ( .A(1'b0), .B(_02906__PTR18), .S(P1_P1_State2_PTR1), .Z(_02907__PTR2) );
  MUX2_X1 U22499 ( .A(1'b0), .B(_02906__PTR19), .S(P1_P1_State2_PTR1), .Z(_02907__PTR3) );
  MUX2_X1 U22500 ( .A(1'b0), .B(_02906__PTR20), .S(P1_P1_State2_PTR1), .Z(_02907__PTR4) );
  MUX2_X1 U22501 ( .A(1'b0), .B(_02906__PTR21), .S(P1_P1_State2_PTR1), .Z(_02907__PTR5) );
  MUX2_X1 U22502 ( .A(1'b0), .B(_02906__PTR22), .S(P1_P1_State2_PTR1), .Z(_02907__PTR6) );
  MUX2_X1 U22503 ( .A(1'b0), .B(_02906__PTR23), .S(P1_P1_State2_PTR1), .Z(_02907__PTR7) );
  MUX2_X1 U22504 ( .A(_02906__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02907__PTR32) );
  MUX2_X1 U22505 ( .A(_02906__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02907__PTR33) );
  MUX2_X1 U22506 ( .A(_02906__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02907__PTR34) );
  MUX2_X1 U22507 ( .A(_02906__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02907__PTR35) );
  MUX2_X1 U22508 ( .A(_02906__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02907__PTR36) );
  MUX2_X1 U22509 ( .A(_02906__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02907__PTR37) );
  MUX2_X1 U22510 ( .A(_02906__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02907__PTR38) );
  MUX2_X1 U22511 ( .A(_02906__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02907__PTR39) );
  MUX2_X1 U22512 ( .A(_01926__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR16) );
  MUX2_X1 U22513 ( .A(_01926__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR17) );
  MUX2_X1 U22514 ( .A(_01926__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR18) );
  MUX2_X1 U22515 ( .A(_01926__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR19) );
  MUX2_X1 U22516 ( .A(_01926__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR20) );
  MUX2_X1 U22517 ( .A(_01926__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR21) );
  MUX2_X1 U22518 ( .A(_01926__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR22) );
  MUX2_X1 U22519 ( .A(_01926__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR23) );
  MUX2_X1 U22520 ( .A(_01926__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR32) );
  MUX2_X1 U22521 ( .A(_01926__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR33) );
  MUX2_X1 U22522 ( .A(_01926__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR34) );
  MUX2_X1 U22523 ( .A(_01926__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR35) );
  MUX2_X1 U22524 ( .A(_01926__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR36) );
  MUX2_X1 U22525 ( .A(_01926__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR37) );
  MUX2_X1 U22526 ( .A(_01926__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR38) );
  MUX2_X1 U22527 ( .A(_01926__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR39) );
  MUX2_X1 U22528 ( .A(_01926__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR64) );
  MUX2_X1 U22529 ( .A(_01926__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR65) );
  MUX2_X1 U22530 ( .A(_01926__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR66) );
  MUX2_X1 U22531 ( .A(_01926__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR67) );
  MUX2_X1 U22532 ( .A(_01926__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR68) );
  MUX2_X1 U22533 ( .A(_01926__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR69) );
  MUX2_X1 U22534 ( .A(_01926__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR70) );
  MUX2_X1 U22535 ( .A(_01926__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02906__PTR71) );
  MUX2_X1 U22536 ( .A(_02911__PTR0), .B(_02909__PTR64), .S(P1_P1_State2_PTR3), .Z(_01929__PTR0) );
  MUX2_X1 U22537 ( .A(_02911__PTR1), .B(_02909__PTR65), .S(P1_P1_State2_PTR3), .Z(_01929__PTR1) );
  MUX2_X1 U22538 ( .A(_02911__PTR2), .B(_02909__PTR66), .S(P1_P1_State2_PTR3), .Z(_01929__PTR2) );
  MUX2_X1 U22539 ( .A(_02911__PTR3), .B(_02909__PTR67), .S(P1_P1_State2_PTR3), .Z(_01929__PTR3) );
  MUX2_X1 U22540 ( .A(_02911__PTR4), .B(_02909__PTR68), .S(P1_P1_State2_PTR3), .Z(_01929__PTR4) );
  MUX2_X1 U22541 ( .A(_02911__PTR5), .B(_02909__PTR69), .S(P1_P1_State2_PTR3), .Z(_01929__PTR5) );
  MUX2_X1 U22542 ( .A(_02911__PTR6), .B(_02909__PTR70), .S(P1_P1_State2_PTR3), .Z(_01929__PTR6) );
  MUX2_X1 U22543 ( .A(_02911__PTR7), .B(_02909__PTR71), .S(P1_P1_State2_PTR3), .Z(_01929__PTR7) );
  MUX2_X1 U22544 ( .A(_02910__PTR0), .B(_02910__PTR32), .S(P1_P1_State2_PTR2), .Z(_02911__PTR0) );
  MUX2_X1 U22545 ( .A(_02910__PTR1), .B(_02910__PTR33), .S(P1_P1_State2_PTR2), .Z(_02911__PTR1) );
  MUX2_X1 U22546 ( .A(_02910__PTR2), .B(_02910__PTR34), .S(P1_P1_State2_PTR2), .Z(_02911__PTR2) );
  MUX2_X1 U22547 ( .A(_02910__PTR3), .B(_02910__PTR35), .S(P1_P1_State2_PTR2), .Z(_02911__PTR3) );
  MUX2_X1 U22548 ( .A(_02910__PTR4), .B(_02910__PTR36), .S(P1_P1_State2_PTR2), .Z(_02911__PTR4) );
  MUX2_X1 U22549 ( .A(_02910__PTR5), .B(_02910__PTR37), .S(P1_P1_State2_PTR2), .Z(_02911__PTR5) );
  MUX2_X1 U22550 ( .A(_02910__PTR6), .B(_02910__PTR38), .S(P1_P1_State2_PTR2), .Z(_02911__PTR6) );
  MUX2_X1 U22551 ( .A(_02910__PTR7), .B(_02910__PTR39), .S(P1_P1_State2_PTR2), .Z(_02911__PTR7) );
  MUX2_X1 U22552 ( .A(1'b0), .B(_02909__PTR16), .S(P1_P1_State2_PTR1), .Z(_02910__PTR0) );
  MUX2_X1 U22553 ( .A(1'b0), .B(_02909__PTR17), .S(P1_P1_State2_PTR1), .Z(_02910__PTR1) );
  MUX2_X1 U22554 ( .A(1'b0), .B(_02909__PTR18), .S(P1_P1_State2_PTR1), .Z(_02910__PTR2) );
  MUX2_X1 U22555 ( .A(1'b0), .B(_02909__PTR19), .S(P1_P1_State2_PTR1), .Z(_02910__PTR3) );
  MUX2_X1 U22556 ( .A(1'b0), .B(_02909__PTR20), .S(P1_P1_State2_PTR1), .Z(_02910__PTR4) );
  MUX2_X1 U22557 ( .A(1'b0), .B(_02909__PTR21), .S(P1_P1_State2_PTR1), .Z(_02910__PTR5) );
  MUX2_X1 U22558 ( .A(1'b0), .B(_02909__PTR22), .S(P1_P1_State2_PTR1), .Z(_02910__PTR6) );
  MUX2_X1 U22559 ( .A(1'b0), .B(_02909__PTR23), .S(P1_P1_State2_PTR1), .Z(_02910__PTR7) );
  MUX2_X1 U22560 ( .A(_02909__PTR32), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02910__PTR32) );
  MUX2_X1 U22561 ( .A(_02909__PTR33), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02910__PTR33) );
  MUX2_X1 U22562 ( .A(_02909__PTR34), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02910__PTR34) );
  MUX2_X1 U22563 ( .A(_02909__PTR35), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02910__PTR35) );
  MUX2_X1 U22564 ( .A(_02909__PTR36), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02910__PTR36) );
  MUX2_X1 U22565 ( .A(_02909__PTR37), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02910__PTR37) );
  MUX2_X1 U22566 ( .A(_02909__PTR38), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02910__PTR38) );
  MUX2_X1 U22567 ( .A(_02909__PTR39), .B(1'b0), .S(P1_P1_State2_PTR1), .Z(_02910__PTR39) );
  MUX2_X1 U22568 ( .A(_01928__PTR16), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR16) );
  MUX2_X1 U22569 ( .A(_01928__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR17) );
  MUX2_X1 U22570 ( .A(_01928__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR18) );
  MUX2_X1 U22571 ( .A(_01928__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR19) );
  MUX2_X1 U22572 ( .A(_01928__PTR20), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR20) );
  MUX2_X1 U22573 ( .A(_01928__PTR21), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR21) );
  MUX2_X1 U22574 ( .A(_01928__PTR22), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR22) );
  MUX2_X1 U22575 ( .A(_01928__PTR23), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR23) );
  MUX2_X1 U22576 ( .A(_01928__PTR32), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR32) );
  MUX2_X1 U22577 ( .A(_01928__PTR33), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR33) );
  MUX2_X1 U22578 ( .A(_01928__PTR34), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR34) );
  MUX2_X1 U22579 ( .A(_01928__PTR35), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR35) );
  MUX2_X1 U22580 ( .A(_01928__PTR36), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR36) );
  MUX2_X1 U22581 ( .A(_01928__PTR37), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR37) );
  MUX2_X1 U22582 ( .A(_01928__PTR38), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR38) );
  MUX2_X1 U22583 ( .A(_01928__PTR39), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR39) );
  MUX2_X1 U22584 ( .A(_01928__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR64) );
  MUX2_X1 U22585 ( .A(_01928__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR65) );
  MUX2_X1 U22586 ( .A(_01928__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR66) );
  MUX2_X1 U22587 ( .A(_01928__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR67) );
  MUX2_X1 U22588 ( .A(_01928__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR68) );
  MUX2_X1 U22589 ( .A(_01928__PTR69), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR69) );
  MUX2_X1 U22590 ( .A(_01928__PTR70), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR70) );
  MUX2_X1 U22591 ( .A(_01928__PTR71), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02909__PTR71) );
  MUX2_X1 U22592 ( .A(_02914__PTR0), .B(_02912__PTR64), .S(P1_P1_State2_PTR3), .Z(_01931__PTR0) );
  MUX2_X1 U22593 ( .A(_02914__PTR1), .B(_02912__PTR65), .S(P1_P1_State2_PTR3), .Z(_01931__PTR1) );
  MUX2_X1 U22594 ( .A(_02914__PTR2), .B(_02912__PTR66), .S(P1_P1_State2_PTR3), .Z(_01931__PTR2) );
  MUX2_X1 U22595 ( .A(_02914__PTR3), .B(_02912__PTR67), .S(P1_P1_State2_PTR3), .Z(_01931__PTR3) );
  MUX2_X1 U22596 ( .A(_02914__PTR4), .B(_02912__PTR68), .S(P1_P1_State2_PTR3), .Z(_01931__PTR4) );
  MUX2_X1 U22597 ( .A(1'b0), .B(_02913__PTR32), .S(P1_P1_State2_PTR2), .Z(_02914__PTR0) );
  MUX2_X1 U22598 ( .A(_02913__PTR1), .B(_02913__PTR33), .S(P1_P1_State2_PTR2), .Z(_02914__PTR1) );
  MUX2_X1 U22599 ( .A(_02913__PTR2), .B(_02913__PTR34), .S(P1_P1_State2_PTR2), .Z(_02914__PTR2) );
  MUX2_X1 U22600 ( .A(_02913__PTR3), .B(_02913__PTR35), .S(P1_P1_State2_PTR2), .Z(_02914__PTR3) );
  MUX2_X1 U22601 ( .A(_02913__PTR4), .B(_02913__PTR36), .S(P1_P1_State2_PTR2), .Z(_02914__PTR4) );
  MUX2_X1 U22602 ( .A(1'b0), .B(_02912__PTR17), .S(P1_P1_State2_PTR1), .Z(_02913__PTR1) );
  MUX2_X1 U22603 ( .A(1'b0), .B(_02912__PTR18), .S(P1_P1_State2_PTR1), .Z(_02913__PTR2) );
  MUX2_X1 U22604 ( .A(1'b0), .B(_02912__PTR19), .S(P1_P1_State2_PTR1), .Z(_02913__PTR3) );
  MUX2_X1 U22605 ( .A(1'b0), .B(_02912__PTR36), .S(P1_P1_State2_PTR1), .Z(_02913__PTR4) );
  MUX2_X1 U22606 ( .A(1'b0), .B(_02912__PTR48), .S(P1_P1_State2_PTR1), .Z(_02913__PTR32) );
  MUX2_X1 U22607 ( .A(_02912__PTR33), .B(_02912__PTR52), .S(P1_P1_State2_PTR1), .Z(_02913__PTR33) );
  MUX2_X1 U22608 ( .A(_02912__PTR34), .B(_02912__PTR52), .S(P1_P1_State2_PTR1), .Z(_02913__PTR34) );
  MUX2_X1 U22609 ( .A(_02912__PTR35), .B(_02912__PTR52), .S(P1_P1_State2_PTR1), .Z(_02913__PTR35) );
  MUX2_X1 U22610 ( .A(_02912__PTR36), .B(_02912__PTR52), .S(P1_P1_State2_PTR1), .Z(_02913__PTR36) );
  MUX2_X1 U22611 ( .A(_01930__PTR17), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02912__PTR17) );
  MUX2_X1 U22612 ( .A(_01930__PTR18), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02912__PTR18) );
  MUX2_X1 U22613 ( .A(_01930__PTR19), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02912__PTR19) );
  MUX2_X1 U22614 ( .A(_01838__PTR1), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02912__PTR33) );
  MUX2_X1 U22615 ( .A(_01838__PTR2), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02912__PTR34) );
  MUX2_X1 U22616 ( .A(_01838__PTR3), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02912__PTR35) );
  MUX2_X1 U22617 ( .A(1'b0), .B(P1_P1_InstQueueWr_Addr_PTR4), .S(P1_P1_State2_PTR0), .Z(_02912__PTR36) );
  MUX2_X1 U22618 ( .A(1'b0), .B(_01930__PTR56), .S(P1_P1_State2_PTR0), .Z(_02912__PTR48) );
  MUX2_X1 U22619 ( .A(1'b0), .B(_01930__PTR60), .S(P1_P1_State2_PTR0), .Z(_02912__PTR52) );
  MUX2_X1 U22620 ( .A(_01930__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02912__PTR64) );
  MUX2_X1 U22621 ( .A(_01930__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02912__PTR65) );
  MUX2_X1 U22622 ( .A(_01930__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02912__PTR66) );
  MUX2_X1 U22623 ( .A(_01930__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02912__PTR67) );
  MUX2_X1 U22624 ( .A(_01930__PTR68), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02912__PTR68) );
  MUX2_X1 U22625 ( .A(_02917__PTR0), .B(_02915__PTR64), .S(P1_P1_State2_PTR3), .Z(_01933__PTR0) );
  MUX2_X1 U22626 ( .A(_02917__PTR1), .B(_02915__PTR65), .S(P1_P1_State2_PTR3), .Z(_01933__PTR1) );
  MUX2_X1 U22627 ( .A(_02917__PTR2), .B(_02915__PTR66), .S(P1_P1_State2_PTR3), .Z(_01933__PTR2) );
  MUX2_X1 U22628 ( .A(_02917__PTR3), .B(_02915__PTR67), .S(P1_P1_State2_PTR3), .Z(_01933__PTR3) );
  MUX2_X1 U22629 ( .A(_02917__PTR4), .B(_02861__PTR32), .S(P1_P1_State2_PTR3), .Z(_01933__PTR4) );
  MUX2_X1 U22630 ( .A(1'b0), .B(_02916__PTR32), .S(P1_P1_State2_PTR2), .Z(_02917__PTR0) );
  MUX2_X1 U22631 ( .A(1'b0), .B(_02916__PTR33), .S(P1_P1_State2_PTR2), .Z(_02917__PTR1) );
  MUX2_X1 U22632 ( .A(1'b0), .B(_02916__PTR34), .S(P1_P1_State2_PTR2), .Z(_02917__PTR2) );
  MUX2_X1 U22633 ( .A(1'b0), .B(_02916__PTR35), .S(P1_P1_State2_PTR2), .Z(_02917__PTR3) );
  MUX2_X1 U22634 ( .A(1'b0), .B(_02916__PTR36), .S(P1_P1_State2_PTR2), .Z(_02917__PTR4) );
  MUX2_X1 U22635 ( .A(_02915__PTR32), .B(_02915__PTR48), .S(P1_P1_State2_PTR1), .Z(_02916__PTR32) );
  MUX2_X1 U22636 ( .A(_02915__PTR33), .B(_02915__PTR49), .S(P1_P1_State2_PTR1), .Z(_02916__PTR33) );
  MUX2_X1 U22637 ( .A(_02915__PTR34), .B(_02915__PTR50), .S(P1_P1_State2_PTR1), .Z(_02916__PTR34) );
  MUX2_X1 U22638 ( .A(_02915__PTR35), .B(_02915__PTR51), .S(P1_P1_State2_PTR1), .Z(_02916__PTR35) );
  MUX2_X1 U22639 ( .A(_02915__PTR36), .B(_02915__PTR52), .S(P1_P1_State2_PTR1), .Z(_02916__PTR36) );
  MUX2_X1 U22640 ( .A(1'b0), .B(_01932__PTR40), .S(P1_P1_State2_PTR0), .Z(_02915__PTR32) );
  MUX2_X1 U22641 ( .A(1'b0), .B(_01932__PTR41), .S(P1_P1_State2_PTR0), .Z(_02915__PTR33) );
  MUX2_X1 U22642 ( .A(1'b0), .B(_01932__PTR42), .S(P1_P1_State2_PTR0), .Z(_02915__PTR34) );
  MUX2_X1 U22643 ( .A(1'b0), .B(_01932__PTR43), .S(P1_P1_State2_PTR0), .Z(_02915__PTR35) );
  MUX2_X1 U22644 ( .A(1'b0), .B(_01932__PTR44), .S(P1_P1_State2_PTR0), .Z(_02915__PTR36) );
  MUX2_X1 U22645 ( .A(1'b0), .B(_01932__PTR56), .S(P1_P1_State2_PTR0), .Z(_02915__PTR48) );
  MUX2_X1 U22646 ( .A(1'b0), .B(_01932__PTR57), .S(P1_P1_State2_PTR0), .Z(_02915__PTR49) );
  MUX2_X1 U22647 ( .A(1'b0), .B(_01932__PTR58), .S(P1_P1_State2_PTR0), .Z(_02915__PTR50) );
  MUX2_X1 U22648 ( .A(1'b0), .B(_01932__PTR59), .S(P1_P1_State2_PTR0), .Z(_02915__PTR51) );
  MUX2_X1 U22649 ( .A(1'b0), .B(_01932__PTR60), .S(P1_P1_State2_PTR0), .Z(_02915__PTR52) );
  MUX2_X1 U22650 ( .A(_01932__PTR64), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02915__PTR64) );
  MUX2_X1 U22651 ( .A(_01932__PTR65), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02915__PTR65) );
  MUX2_X1 U22652 ( .A(_01932__PTR66), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02915__PTR66) );
  MUX2_X1 U22653 ( .A(_01932__PTR67), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02915__PTR67) );
  MUX2_X1 U22654 ( .A(_02918__PTR256), .B(_02918__PTR384), .S(P1_P1_State2_PTR1), .Z(_02919__PTR256) );
  MUX2_X1 U22655 ( .A(_02918__PTR257), .B(_02918__PTR385), .S(P1_P1_State2_PTR1), .Z(_02919__PTR257) );
  MUX2_X1 U22656 ( .A(_02918__PTR258), .B(_02918__PTR386), .S(P1_P1_State2_PTR1), .Z(_02919__PTR258) );
  MUX2_X1 U22657 ( .A(_02918__PTR259), .B(_02918__PTR387), .S(P1_P1_State2_PTR1), .Z(_02919__PTR259) );
  MUX2_X1 U22658 ( .A(_02918__PTR260), .B(_02918__PTR388), .S(P1_P1_State2_PTR1), .Z(_02919__PTR260) );
  MUX2_X1 U22659 ( .A(_02918__PTR261), .B(_02918__PTR389), .S(P1_P1_State2_PTR1), .Z(_02919__PTR261) );
  MUX2_X1 U22660 ( .A(_02918__PTR262), .B(_02918__PTR390), .S(P1_P1_State2_PTR1), .Z(_02919__PTR262) );
  MUX2_X1 U22661 ( .A(_02918__PTR263), .B(_02918__PTR391), .S(P1_P1_State2_PTR1), .Z(_02919__PTR263) );
  MUX2_X1 U22662 ( .A(_02918__PTR264), .B(_02918__PTR392), .S(P1_P1_State2_PTR1), .Z(_02919__PTR264) );
  MUX2_X1 U22663 ( .A(_02918__PTR265), .B(_02918__PTR393), .S(P1_P1_State2_PTR1), .Z(_02919__PTR265) );
  MUX2_X1 U22664 ( .A(_02918__PTR266), .B(_02918__PTR394), .S(P1_P1_State2_PTR1), .Z(_02919__PTR266) );
  MUX2_X1 U22665 ( .A(_02918__PTR267), .B(_02918__PTR395), .S(P1_P1_State2_PTR1), .Z(_02919__PTR267) );
  MUX2_X1 U22666 ( .A(_02918__PTR268), .B(_02918__PTR396), .S(P1_P1_State2_PTR1), .Z(_02919__PTR268) );
  MUX2_X1 U22667 ( .A(_02918__PTR269), .B(_02918__PTR397), .S(P1_P1_State2_PTR1), .Z(_02919__PTR269) );
  MUX2_X1 U22668 ( .A(_02918__PTR270), .B(_02918__PTR398), .S(P1_P1_State2_PTR1), .Z(_02919__PTR270) );
  MUX2_X1 U22669 ( .A(_02918__PTR271), .B(_02918__PTR399), .S(P1_P1_State2_PTR1), .Z(_02919__PTR271) );
  MUX2_X1 U22670 ( .A(_02918__PTR272), .B(_02918__PTR400), .S(P1_P1_State2_PTR1), .Z(_02919__PTR272) );
  MUX2_X1 U22671 ( .A(_02918__PTR273), .B(_02918__PTR401), .S(P1_P1_State2_PTR1), .Z(_02919__PTR273) );
  MUX2_X1 U22672 ( .A(_02918__PTR274), .B(_02918__PTR402), .S(P1_P1_State2_PTR1), .Z(_02919__PTR274) );
  MUX2_X1 U22673 ( .A(_02918__PTR275), .B(_02918__PTR403), .S(P1_P1_State2_PTR1), .Z(_02919__PTR275) );
  MUX2_X1 U22674 ( .A(_02918__PTR276), .B(_02918__PTR404), .S(P1_P1_State2_PTR1), .Z(_02919__PTR276) );
  MUX2_X1 U22675 ( .A(_02918__PTR277), .B(_02918__PTR405), .S(P1_P1_State2_PTR1), .Z(_02919__PTR277) );
  MUX2_X1 U22676 ( .A(_02918__PTR278), .B(_02918__PTR406), .S(P1_P1_State2_PTR1), .Z(_02919__PTR278) );
  MUX2_X1 U22677 ( .A(_02918__PTR279), .B(_02918__PTR407), .S(P1_P1_State2_PTR1), .Z(_02919__PTR279) );
  MUX2_X1 U22678 ( .A(_02918__PTR280), .B(_02918__PTR408), .S(P1_P1_State2_PTR1), .Z(_02919__PTR280) );
  MUX2_X1 U22679 ( .A(_02918__PTR281), .B(_02918__PTR409), .S(P1_P1_State2_PTR1), .Z(_02919__PTR281) );
  MUX2_X1 U22680 ( .A(_02918__PTR282), .B(_02918__PTR410), .S(P1_P1_State2_PTR1), .Z(_02919__PTR282) );
  MUX2_X1 U22681 ( .A(_02918__PTR283), .B(_02918__PTR411), .S(P1_P1_State2_PTR1), .Z(_02919__PTR283) );
  MUX2_X1 U22682 ( .A(_02918__PTR284), .B(_02918__PTR412), .S(P1_P1_State2_PTR1), .Z(_02919__PTR284) );
  MUX2_X1 U22683 ( .A(_02918__PTR285), .B(_02918__PTR413), .S(P1_P1_State2_PTR1), .Z(_02919__PTR285) );
  MUX2_X1 U22684 ( .A(_02918__PTR286), .B(_02918__PTR414), .S(P1_P1_State2_PTR1), .Z(_02919__PTR286) );
  MUX2_X1 U22685 ( .A(_02918__PTR288), .B(_02861__PTR32), .S(P1_P1_State2_PTR1), .Z(_02919__PTR288) );
  MUX2_X1 U22686 ( .A(1'b0), .B(_01938__PTR320), .S(P1_P1_State2_PTR0), .Z(_02918__PTR256) );
  MUX2_X1 U22687 ( .A(1'b0), .B(_01938__PTR321), .S(P1_P1_State2_PTR0), .Z(_02918__PTR257) );
  MUX2_X1 U22688 ( .A(1'b0), .B(_01938__PTR322), .S(P1_P1_State2_PTR0), .Z(_02918__PTR258) );
  MUX2_X1 U22689 ( .A(1'b0), .B(_01938__PTR323), .S(P1_P1_State2_PTR0), .Z(_02918__PTR259) );
  MUX2_X1 U22690 ( .A(1'b0), .B(_01938__PTR324), .S(P1_P1_State2_PTR0), .Z(_02918__PTR260) );
  MUX2_X1 U22691 ( .A(1'b0), .B(_01938__PTR325), .S(P1_P1_State2_PTR0), .Z(_02918__PTR261) );
  MUX2_X1 U22692 ( .A(1'b0), .B(_01938__PTR326), .S(P1_P1_State2_PTR0), .Z(_02918__PTR262) );
  MUX2_X1 U22693 ( .A(1'b0), .B(_01938__PTR327), .S(P1_P1_State2_PTR0), .Z(_02918__PTR263) );
  MUX2_X1 U22694 ( .A(1'b0), .B(_01938__PTR328), .S(P1_P1_State2_PTR0), .Z(_02918__PTR264) );
  MUX2_X1 U22695 ( .A(1'b0), .B(_01938__PTR329), .S(P1_P1_State2_PTR0), .Z(_02918__PTR265) );
  MUX2_X1 U22696 ( .A(1'b0), .B(_01938__PTR330), .S(P1_P1_State2_PTR0), .Z(_02918__PTR266) );
  MUX2_X1 U22697 ( .A(1'b0), .B(_01938__PTR331), .S(P1_P1_State2_PTR0), .Z(_02918__PTR267) );
  MUX2_X1 U22698 ( .A(1'b0), .B(_01938__PTR332), .S(P1_P1_State2_PTR0), .Z(_02918__PTR268) );
  MUX2_X1 U22699 ( .A(1'b0), .B(_01938__PTR333), .S(P1_P1_State2_PTR0), .Z(_02918__PTR269) );
  MUX2_X1 U22700 ( .A(1'b0), .B(_01938__PTR334), .S(P1_P1_State2_PTR0), .Z(_02918__PTR270) );
  MUX2_X1 U22701 ( .A(1'b0), .B(_01938__PTR335), .S(P1_P1_State2_PTR0), .Z(_02918__PTR271) );
  MUX2_X1 U22702 ( .A(1'b0), .B(_01938__PTR336), .S(P1_P1_State2_PTR0), .Z(_02918__PTR272) );
  MUX2_X1 U22703 ( .A(1'b0), .B(_01938__PTR337), .S(P1_P1_State2_PTR0), .Z(_02918__PTR273) );
  MUX2_X1 U22704 ( .A(1'b0), .B(_01938__PTR338), .S(P1_P1_State2_PTR0), .Z(_02918__PTR274) );
  MUX2_X1 U22705 ( .A(1'b0), .B(_01938__PTR339), .S(P1_P1_State2_PTR0), .Z(_02918__PTR275) );
  MUX2_X1 U22706 ( .A(1'b0), .B(_01938__PTR340), .S(P1_P1_State2_PTR0), .Z(_02918__PTR276) );
  MUX2_X1 U22707 ( .A(1'b0), .B(_01938__PTR341), .S(P1_P1_State2_PTR0), .Z(_02918__PTR277) );
  MUX2_X1 U22708 ( .A(1'b0), .B(_01938__PTR342), .S(P1_P1_State2_PTR0), .Z(_02918__PTR278) );
  MUX2_X1 U22709 ( .A(1'b0), .B(_01938__PTR343), .S(P1_P1_State2_PTR0), .Z(_02918__PTR279) );
  MUX2_X1 U22710 ( .A(1'b0), .B(_01938__PTR344), .S(P1_P1_State2_PTR0), .Z(_02918__PTR280) );
  MUX2_X1 U22711 ( .A(1'b0), .B(_01938__PTR345), .S(P1_P1_State2_PTR0), .Z(_02918__PTR281) );
  MUX2_X1 U22712 ( .A(1'b0), .B(_01938__PTR346), .S(P1_P1_State2_PTR0), .Z(_02918__PTR282) );
  MUX2_X1 U22713 ( .A(1'b0), .B(_01938__PTR347), .S(P1_P1_State2_PTR0), .Z(_02918__PTR283) );
  MUX2_X1 U22714 ( .A(1'b0), .B(_01938__PTR348), .S(P1_P1_State2_PTR0), .Z(_02918__PTR284) );
  MUX2_X1 U22715 ( .A(1'b0), .B(_01938__PTR349), .S(P1_P1_State2_PTR0), .Z(_02918__PTR285) );
  MUX2_X1 U22716 ( .A(1'b0), .B(_01938__PTR350), .S(P1_P1_State2_PTR0), .Z(_02918__PTR286) );
  MUX2_X1 U22717 ( .A(1'b0), .B(_01938__PTR352), .S(P1_P1_State2_PTR0), .Z(_02918__PTR288) );
  MUX2_X1 U22718 ( .A(P1_P1_lWord_PTR0), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR384) );
  MUX2_X1 U22719 ( .A(P1_P1_lWord_PTR1), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR385) );
  MUX2_X1 U22720 ( .A(P1_P1_lWord_PTR2), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR386) );
  MUX2_X1 U22721 ( .A(P1_P1_lWord_PTR3), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR387) );
  MUX2_X1 U22722 ( .A(P1_P1_lWord_PTR4), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR388) );
  MUX2_X1 U22723 ( .A(P1_P1_lWord_PTR5), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR389) );
  MUX2_X1 U22724 ( .A(P1_P1_lWord_PTR6), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR390) );
  MUX2_X1 U22725 ( .A(P1_P1_lWord_PTR7), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR391) );
  MUX2_X1 U22726 ( .A(P1_P1_lWord_PTR8), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR392) );
  MUX2_X1 U22727 ( .A(P1_P1_lWord_PTR9), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR393) );
  MUX2_X1 U22728 ( .A(P1_P1_lWord_PTR10), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR394) );
  MUX2_X1 U22729 ( .A(P1_P1_lWord_PTR11), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR395) );
  MUX2_X1 U22730 ( .A(P1_P1_lWord_PTR12), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR396) );
  MUX2_X1 U22731 ( .A(P1_P1_lWord_PTR13), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR397) );
  MUX2_X1 U22732 ( .A(P1_P1_lWord_PTR14), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR398) );
  MUX2_X1 U22733 ( .A(P1_P1_lWord_PTR15), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR399) );
  MUX2_X1 U22734 ( .A(P1_P1_uWord_PTR0), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR400) );
  MUX2_X1 U22735 ( .A(P1_P1_uWord_PTR1), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR401) );
  MUX2_X1 U22736 ( .A(P1_P1_uWord_PTR2), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR402) );
  MUX2_X1 U22737 ( .A(P1_P1_uWord_PTR3), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR403) );
  MUX2_X1 U22738 ( .A(P1_P1_uWord_PTR4), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR404) );
  MUX2_X1 U22739 ( .A(P1_P1_uWord_PTR5), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR405) );
  MUX2_X1 U22740 ( .A(P1_P1_uWord_PTR6), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR406) );
  MUX2_X1 U22741 ( .A(P1_P1_uWord_PTR7), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR407) );
  MUX2_X1 U22742 ( .A(P1_P1_uWord_PTR8), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR408) );
  MUX2_X1 U22743 ( .A(P1_P1_uWord_PTR9), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR409) );
  MUX2_X1 U22744 ( .A(P1_P1_uWord_PTR10), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR410) );
  MUX2_X1 U22745 ( .A(P1_P1_uWord_PTR11), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR411) );
  MUX2_X1 U22746 ( .A(P1_P1_uWord_PTR12), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR412) );
  MUX2_X1 U22747 ( .A(P1_P1_uWord_PTR13), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR413) );
  MUX2_X1 U22748 ( .A(P1_P1_uWord_PTR14), .B(1'b0), .S(P1_P1_State2_PTR0), .Z(_02918__PTR414) );
  MUX2_X1 U22749 ( .A(_02951__PTR0), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR0) );
  MUX2_X1 U22750 ( .A(_02951__PTR1), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR1) );
  MUX2_X1 U22751 ( .A(_02951__PTR2), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR2) );
  MUX2_X1 U22752 ( .A(_02951__PTR3), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR3) );
  MUX2_X1 U22753 ( .A(_02951__PTR4), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR4) );
  MUX2_X1 U22754 ( .A(_02951__PTR5), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR5) );
  MUX2_X1 U22755 ( .A(_02951__PTR6), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR6) );
  MUX2_X1 U22756 ( .A(_02951__PTR7), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR7) );
  MUX2_X1 U22757 ( .A(1'b0), .B(_02951__PTR0), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR8) );
  MUX2_X1 U22758 ( .A(1'b0), .B(_02951__PTR1), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR9) );
  MUX2_X1 U22759 ( .A(1'b0), .B(_02951__PTR2), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR10) );
  MUX2_X1 U22760 ( .A(1'b0), .B(_02951__PTR3), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR11) );
  MUX2_X1 U22761 ( .A(1'b0), .B(_02951__PTR4), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR12) );
  MUX2_X1 U22762 ( .A(1'b0), .B(_02951__PTR5), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR13) );
  MUX2_X1 U22763 ( .A(1'b0), .B(_02951__PTR6), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR14) );
  MUX2_X1 U22764 ( .A(1'b0), .B(_02951__PTR7), .S(P2_P1_InstQueueWr_Addr_PTR3), .Z(_02128__PTR15) );
  MUX2_X1 U22765 ( .A(_02950__PTR0), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR2), .Z(_02951__PTR0) );
  MUX2_X1 U22766 ( .A(_02950__PTR1), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR2), .Z(_02951__PTR1) );
  MUX2_X1 U22767 ( .A(_02950__PTR2), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR2), .Z(_02951__PTR2) );
  MUX2_X1 U22768 ( .A(_02950__PTR3), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR2), .Z(_02951__PTR3) );
  MUX2_X1 U22769 ( .A(1'b0), .B(_02950__PTR0), .S(P2_P1_InstQueueWr_Addr_PTR2), .Z(_02951__PTR4) );
  MUX2_X1 U22770 ( .A(1'b0), .B(_02950__PTR1), .S(P2_P1_InstQueueWr_Addr_PTR2), .Z(_02951__PTR5) );
  MUX2_X1 U22771 ( .A(1'b0), .B(_02950__PTR2), .S(P2_P1_InstQueueWr_Addr_PTR2), .Z(_02951__PTR6) );
  MUX2_X1 U22772 ( .A(1'b0), .B(_02950__PTR3), .S(P2_P1_InstQueueWr_Addr_PTR2), .Z(_02951__PTR7) );
  MUX2_X1 U22773 ( .A(_02129__PTR0), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR1), .Z(_02950__PTR0) );
  MUX2_X1 U22774 ( .A(P2_P1_InstQueueWr_Addr_PTR0), .B(1'b0), .S(P2_P1_InstQueueWr_Addr_PTR1), .Z(_02950__PTR1) );
  MUX2_X1 U22775 ( .A(1'b0), .B(_02129__PTR0), .S(P2_P1_InstQueueWr_Addr_PTR1), .Z(_02950__PTR2) );
  MUX2_X1 U22776 ( .A(1'b0), .B(P2_P1_InstQueueWr_Addr_PTR0), .S(P2_P1_InstQueueWr_Addr_PTR1), .Z(_02950__PTR3) );
  MUX2_X1 U22777 ( .A(_02953__PTR0), .B(1'b0), .S(_02129__PTR3), .Z(_02130__PTR0) );
  MUX2_X1 U22778 ( .A(_02953__PTR1), .B(1'b0), .S(_02129__PTR3), .Z(_02130__PTR1) );
  MUX2_X1 U22779 ( .A(_02953__PTR2), .B(1'b0), .S(_02129__PTR3), .Z(_02130__PTR2) );
  MUX2_X1 U22780 ( .A(_02953__PTR3), .B(1'b0), .S(_02129__PTR3), .Z(_02130__PTR3) );
  MUX2_X1 U22781 ( .A(_02953__PTR4), .B(1'b0), .S(_02129__PTR3), .Z(_02130__PTR4) );
  MUX2_X1 U22782 ( .A(_02953__PTR5), .B(1'b0), .S(_02129__PTR3), .Z(_02130__PTR5) );
  MUX2_X1 U22783 ( .A(_02953__PTR6), .B(1'b0), .S(_02129__PTR3), .Z(_02130__PTR6) );
  MUX2_X1 U22784 ( .A(_02953__PTR7), .B(1'b0), .S(_02129__PTR3), .Z(_02130__PTR7) );
  MUX2_X1 U22785 ( .A(1'b0), .B(_02953__PTR0), .S(_02129__PTR3), .Z(_02130__PTR8) );
  MUX2_X1 U22786 ( .A(1'b0), .B(_02953__PTR1), .S(_02129__PTR3), .Z(_02130__PTR9) );
  MUX2_X1 U22787 ( .A(1'b0), .B(_02953__PTR2), .S(_02129__PTR3), .Z(_02130__PTR10) );
  MUX2_X1 U22788 ( .A(1'b0), .B(_02953__PTR3), .S(_02129__PTR3), .Z(_02130__PTR11) );
  MUX2_X1 U22789 ( .A(1'b0), .B(_02953__PTR4), .S(_02129__PTR3), .Z(_02130__PTR12) );
  MUX2_X1 U22790 ( .A(1'b0), .B(_02953__PTR5), .S(_02129__PTR3), .Z(_02130__PTR13) );
  MUX2_X1 U22791 ( .A(1'b0), .B(_02953__PTR6), .S(_02129__PTR3), .Z(_02130__PTR14) );
  MUX2_X1 U22792 ( .A(1'b0), .B(_02953__PTR7), .S(_02129__PTR3), .Z(_02130__PTR15) );
  MUX2_X1 U22793 ( .A(_02952__PTR0), .B(1'b0), .S(_02129__PTR2), .Z(_02953__PTR0) );
  MUX2_X1 U22794 ( .A(_02952__PTR1), .B(1'b0), .S(_02129__PTR2), .Z(_02953__PTR1) );
  MUX2_X1 U22795 ( .A(_02952__PTR2), .B(1'b0), .S(_02129__PTR2), .Z(_02953__PTR2) );
  MUX2_X1 U22796 ( .A(_02952__PTR3), .B(1'b0), .S(_02129__PTR2), .Z(_02953__PTR3) );
  MUX2_X1 U22797 ( .A(1'b0), .B(_02952__PTR0), .S(_02129__PTR2), .Z(_02953__PTR4) );
  MUX2_X1 U22798 ( .A(1'b0), .B(_02952__PTR1), .S(_02129__PTR2), .Z(_02953__PTR5) );
  MUX2_X1 U22799 ( .A(1'b0), .B(_02952__PTR2), .S(_02129__PTR2), .Z(_02953__PTR6) );
  MUX2_X1 U22800 ( .A(1'b0), .B(_02952__PTR3), .S(_02129__PTR2), .Z(_02953__PTR7) );
  MUX2_X1 U22801 ( .A(P2_P1_InstQueueWr_Addr_PTR0), .B(1'b0), .S(_02129__PTR1), .Z(_02952__PTR0) );
  MUX2_X1 U22802 ( .A(_02129__PTR0), .B(1'b0), .S(_02129__PTR1), .Z(_02952__PTR1) );
  MUX2_X1 U22803 ( .A(1'b0), .B(P2_P1_InstQueueWr_Addr_PTR0), .S(_02129__PTR1), .Z(_02952__PTR2) );
  MUX2_X1 U22804 ( .A(1'b0), .B(_02129__PTR0), .S(_02129__PTR1), .Z(_02952__PTR3) );
  MUX2_X1 U22805 ( .A(_02955__PTR0), .B(1'b0), .S(_02131__PTR3), .Z(_02132__PTR0) );
  MUX2_X1 U22806 ( .A(_02955__PTR1), .B(1'b0), .S(_02131__PTR3), .Z(_02132__PTR1) );
  MUX2_X1 U22807 ( .A(_02955__PTR2), .B(1'b0), .S(_02131__PTR3), .Z(_02132__PTR2) );
  MUX2_X1 U22808 ( .A(_02955__PTR3), .B(1'b0), .S(_02131__PTR3), .Z(_02132__PTR3) );
  MUX2_X1 U22809 ( .A(_02955__PTR4), .B(1'b0), .S(_02131__PTR3), .Z(_02132__PTR4) );
  MUX2_X1 U22810 ( .A(_02955__PTR5), .B(1'b0), .S(_02131__PTR3), .Z(_02132__PTR5) );
  MUX2_X1 U22811 ( .A(_02955__PTR6), .B(1'b0), .S(_02131__PTR3), .Z(_02132__PTR6) );
  MUX2_X1 U22812 ( .A(_02955__PTR7), .B(1'b0), .S(_02131__PTR3), .Z(_02132__PTR7) );
  MUX2_X1 U22813 ( .A(1'b0), .B(_02955__PTR0), .S(_02131__PTR3), .Z(_02132__PTR8) );
  MUX2_X1 U22814 ( .A(1'b0), .B(_02955__PTR1), .S(_02131__PTR3), .Z(_02132__PTR9) );
  MUX2_X1 U22815 ( .A(1'b0), .B(_02955__PTR2), .S(_02131__PTR3), .Z(_02132__PTR10) );
  MUX2_X1 U22816 ( .A(1'b0), .B(_02955__PTR3), .S(_02131__PTR3), .Z(_02132__PTR11) );
  MUX2_X1 U22817 ( .A(1'b0), .B(_02955__PTR4), .S(_02131__PTR3), .Z(_02132__PTR12) );
  MUX2_X1 U22818 ( .A(1'b0), .B(_02955__PTR5), .S(_02131__PTR3), .Z(_02132__PTR13) );
  MUX2_X1 U22819 ( .A(1'b0), .B(_02955__PTR6), .S(_02131__PTR3), .Z(_02132__PTR14) );
  MUX2_X1 U22820 ( .A(1'b0), .B(_02955__PTR7), .S(_02131__PTR3), .Z(_02132__PTR15) );
  MUX2_X1 U22821 ( .A(_02954__PTR0), .B(1'b0), .S(_02131__PTR2), .Z(_02955__PTR0) );
  MUX2_X1 U22822 ( .A(_02954__PTR1), .B(1'b0), .S(_02131__PTR2), .Z(_02955__PTR1) );
  MUX2_X1 U22823 ( .A(_02954__PTR2), .B(1'b0), .S(_02131__PTR2), .Z(_02955__PTR2) );
  MUX2_X1 U22824 ( .A(_02954__PTR3), .B(1'b0), .S(_02131__PTR2), .Z(_02955__PTR3) );
  MUX2_X1 U22825 ( .A(1'b0), .B(_02954__PTR0), .S(_02131__PTR2), .Z(_02955__PTR4) );
  MUX2_X1 U22826 ( .A(1'b0), .B(_02954__PTR1), .S(_02131__PTR2), .Z(_02955__PTR5) );
  MUX2_X1 U22827 ( .A(1'b0), .B(_02954__PTR2), .S(_02131__PTR2), .Z(_02955__PTR6) );
  MUX2_X1 U22828 ( .A(1'b0), .B(_02954__PTR3), .S(_02131__PTR2), .Z(_02955__PTR7) );
  MUX2_X1 U22829 ( .A(_02129__PTR0), .B(1'b0), .S(_02131__PTR1), .Z(_02954__PTR0) );
  MUX2_X1 U22830 ( .A(P2_P1_InstQueueWr_Addr_PTR0), .B(1'b0), .S(_02131__PTR1), .Z(_02954__PTR1) );
  MUX2_X1 U22831 ( .A(1'b0), .B(_02129__PTR0), .S(_02131__PTR1), .Z(_02954__PTR2) );
  MUX2_X1 U22832 ( .A(1'b0), .B(P2_P1_InstQueueWr_Addr_PTR0), .S(_02131__PTR1), .Z(_02954__PTR3) );
  MUX2_X1 U22833 ( .A(_02957__PTR0), .B(1'b0), .S(_02133__PTR3), .Z(_02134__PTR0) );
  MUX2_X1 U22834 ( .A(_02957__PTR1), .B(1'b0), .S(_02133__PTR3), .Z(_02134__PTR1) );
  MUX2_X1 U22835 ( .A(_02957__PTR2), .B(1'b0), .S(_02133__PTR3), .Z(_02134__PTR2) );
  MUX2_X1 U22836 ( .A(_02957__PTR3), .B(1'b0), .S(_02133__PTR3), .Z(_02134__PTR3) );
  MUX2_X1 U22837 ( .A(_02957__PTR4), .B(1'b0), .S(_02133__PTR3), .Z(_02134__PTR4) );
  MUX2_X1 U22838 ( .A(_02957__PTR5), .B(1'b0), .S(_02133__PTR3), .Z(_02134__PTR5) );
  MUX2_X1 U22839 ( .A(_02957__PTR6), .B(1'b0), .S(_02133__PTR3), .Z(_02134__PTR6) );
  MUX2_X1 U22840 ( .A(_02957__PTR7), .B(1'b0), .S(_02133__PTR3), .Z(_02134__PTR7) );
  MUX2_X1 U22841 ( .A(1'b0), .B(_02957__PTR0), .S(_02133__PTR3), .Z(_02134__PTR8) );
  MUX2_X1 U22842 ( .A(1'b0), .B(_02957__PTR1), .S(_02133__PTR3), .Z(_02134__PTR9) );
  MUX2_X1 U22843 ( .A(1'b0), .B(_02957__PTR2), .S(_02133__PTR3), .Z(_02134__PTR10) );
  MUX2_X1 U22844 ( .A(1'b0), .B(_02957__PTR3), .S(_02133__PTR3), .Z(_02134__PTR11) );
  MUX2_X1 U22845 ( .A(1'b0), .B(_02957__PTR4), .S(_02133__PTR3), .Z(_02134__PTR12) );
  MUX2_X1 U22846 ( .A(1'b0), .B(_02957__PTR5), .S(_02133__PTR3), .Z(_02134__PTR13) );
  MUX2_X1 U22847 ( .A(1'b0), .B(_02957__PTR6), .S(_02133__PTR3), .Z(_02134__PTR14) );
  MUX2_X1 U22848 ( .A(1'b0), .B(_02957__PTR7), .S(_02133__PTR3), .Z(_02134__PTR15) );
  MUX2_X1 U22849 ( .A(_02956__PTR0), .B(1'b0), .S(_02133__PTR2), .Z(_02957__PTR0) );
  MUX2_X1 U22850 ( .A(_02956__PTR1), .B(1'b0), .S(_02133__PTR2), .Z(_02957__PTR1) );
  MUX2_X1 U22851 ( .A(_02956__PTR2), .B(1'b0), .S(_02133__PTR2), .Z(_02957__PTR2) );
  MUX2_X1 U22852 ( .A(_02956__PTR3), .B(1'b0), .S(_02133__PTR2), .Z(_02957__PTR3) );
  MUX2_X1 U22853 ( .A(1'b0), .B(_02956__PTR0), .S(_02133__PTR2), .Z(_02957__PTR4) );
  MUX2_X1 U22854 ( .A(1'b0), .B(_02956__PTR1), .S(_02133__PTR2), .Z(_02957__PTR5) );
  MUX2_X1 U22855 ( .A(1'b0), .B(_02956__PTR2), .S(_02133__PTR2), .Z(_02957__PTR6) );
  MUX2_X1 U22856 ( .A(1'b0), .B(_02956__PTR3), .S(_02133__PTR2), .Z(_02957__PTR7) );
  MUX2_X1 U22857 ( .A(P2_P1_InstQueueWr_Addr_PTR0), .B(1'b0), .S(_02133__PTR1), .Z(_02956__PTR0) );
  MUX2_X1 U22858 ( .A(_02129__PTR0), .B(1'b0), .S(_02133__PTR1), .Z(_02956__PTR1) );
  MUX2_X1 U22859 ( .A(1'b0), .B(P2_P1_InstQueueWr_Addr_PTR0), .S(_02133__PTR1), .Z(_02956__PTR2) );
  MUX2_X1 U22860 ( .A(1'b0), .B(_02129__PTR0), .S(_02133__PTR1), .Z(_02956__PTR3) );
  MUX2_X1 U22861 ( .A(_03000__PTR0), .B(_03000__PTR4), .S(P2_State_PTR2), .Z(_02136_) );
  MUX2_X1 U22862 ( .A(_02999__PTR0), .B(_02999__PTR6), .S(P2_State_PTR1), .Z(_03000__PTR0) );
  MUX2_X1 U22863 ( .A(1'b0), .B(_02999__PTR6), .S(P2_State_PTR1), .Z(_03000__PTR4) );
  MUX2_X1 U22864 ( .A(1'b1), .B(1'b0), .S(P2_State_PTR0), .Z(_02999__PTR0) );
  MUX2_X1 U22865 ( .A(_02135__PTR6), .B(P2_D_C_n), .S(P2_State_PTR0), .Z(_02999__PTR6) );
  MUX2_X1 U22866 ( .A(_03002__PTR0), .B(_03002__PTR4), .S(P2_State_PTR2), .Z(_02137_) );
  MUX2_X1 U22867 ( .A(_03001__PTR4), .B(P2_State_PTR0), .S(P2_State_PTR1), .Z(_03002__PTR0) );
  MUX2_X1 U22868 ( .A(_03001__PTR4), .B(_03001__PTR6), .S(P2_State_PTR1), .Z(_03002__PTR4) );
  MUX2_X1 U22869 ( .A(1'b1), .B(P2_ADS_n), .S(P2_State_PTR0), .Z(_03001__PTR4) );
  MUX2_X1 U22870 ( .A(1'b0), .B(1'b0), .S(P2_State_PTR0), .Z(_03001__PTR6) );
  MUX2_X1 U22871 ( .A(_03004__PTR0), .B(_03004__PTR4), .S(P2_State_PTR2), .Z(_02138_) );
  MUX2_X1 U22872 ( .A(_02999__PTR0), .B(_03003__PTR2), .S(P2_State_PTR1), .Z(_03004__PTR0) );
  MUX2_X1 U22873 ( .A(_03003__PTR4), .B(1'b0), .S(P2_State_PTR1), .Z(_03004__PTR4) );
  MUX2_X1 U22874 ( .A(1'b0), .B(bs16), .S(P2_State_PTR0), .Z(_03003__PTR2) );
  MUX2_X1 U22875 ( .A(bs16), .B(1'b0), .S(P2_State_PTR0), .Z(_03003__PTR4) );
  MUX2_X1 U22876 ( .A(_03006__PTR0), .B(_03006__PTR4), .S(P2_P1_State2_PTR2), .Z(_03007__PTR0) );
  MUX2_X1 U22877 ( .A(1'b1), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03006__PTR0) );
  MUX2_X1 U22878 ( .A(_03005__PTR4), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03006__PTR4) );
  MUX2_X1 U22879 ( .A(1'b0), .B(_02140__PTR5), .S(P2_P1_State2_PTR0), .Z(_03005__PTR4) );
  MUX2_X1 U22880 ( .A(_03006__PTR0), .B(_03009__PTR4), .S(P2_P1_State2_PTR2), .Z(_03010__PTR0) );
  MUX2_X1 U22881 ( .A(_03008__PTR4), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03009__PTR4) );
  MUX2_X1 U22882 ( .A(1'b0), .B(_02141__PTR5), .S(P2_P1_State2_PTR0), .Z(_03008__PTR4) );
  MUX2_X1 U22883 ( .A(_03012__PTR0), .B(_03012__PTR4), .S(P2_P1_State2_PTR2), .Z(_03013__PTR0) );
  MUX2_X1 U22884 ( .A(1'b1), .B(P2_P1_State2_PTR0), .S(P2_P1_State2_PTR1), .Z(_03012__PTR0) );
  MUX2_X1 U22885 ( .A(_03011__PTR4), .B(_03011__PTR6), .S(P2_P1_State2_PTR1), .Z(_03012__PTR4) );
  MUX2_X1 U22886 ( .A(1'b0), .B(_02142__PTR5), .S(P2_P1_State2_PTR0), .Z(_03011__PTR4) );
  MUX2_X1 U22887 ( .A(_02142__PTR6), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03011__PTR6) );
  MUX2_X1 U22888 ( .A(_03015__PTR0), .B(_03015__PTR4), .S(P2_P1_State2_PTR2), .Z(_03016__PTR0) );
  MUX2_X1 U22889 ( .A(_03014__PTR0), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03015__PTR0) );
  MUX2_X1 U22890 ( .A(_03014__PTR4), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03015__PTR4) );
  MUX2_X1 U22891 ( .A(1'b0), .B(1'b1), .S(P2_P1_State2_PTR0), .Z(_03014__PTR0) );
  MUX2_X1 U22892 ( .A(1'b0), .B(_02143__PTR5), .S(P2_P1_State2_PTR0), .Z(_03014__PTR4) );
  MUX2_X1 U22893 ( .A(_03077__PTR0), .B(_03077__PTR16), .S(P2_State_PTR2), .Z(_02170__PTR0) );
  MUX2_X1 U22894 ( .A(_03077__PTR1), .B(_03077__PTR17), .S(P2_State_PTR2), .Z(_02170__PTR1) );
  MUX2_X1 U22895 ( .A(_03077__PTR2), .B(_03077__PTR18), .S(P2_State_PTR2), .Z(_02170__PTR2) );
  MUX2_X1 U22896 ( .A(_03079__PTR0), .B(_03078__PTR0), .S(P2_State_PTR1), .Z(_03077__PTR0) );
  MUX2_X1 U22897 ( .A(_03079__PTR1), .B(_03078__PTR1), .S(P2_State_PTR1), .Z(_03077__PTR1) );
  MUX2_X1 U22898 ( .A(_03079__PTR2), .B(_03078__PTR2), .S(P2_State_PTR1), .Z(_03077__PTR2) );
  MUX2_X1 U22899 ( .A(_03078__PTR8), .B(_03078__PTR16), .S(P2_State_PTR1), .Z(_03077__PTR16) );
  MUX2_X1 U22900 ( .A(_03078__PTR9), .B(_03078__PTR17), .S(P2_State_PTR1), .Z(_03077__PTR17) );
  MUX2_X1 U22901 ( .A(_03078__PTR10), .B(_03078__PTR18), .S(P2_State_PTR1), .Z(_03077__PTR18) );
  MUX2_X1 U22902 ( .A(1'b1), .B(_02169__PTR4), .S(P2_State_PTR0), .Z(_03079__PTR0) );
  MUX2_X1 U22903 ( .A(1'b0), .B(P2_RequestPending), .S(P2_State_PTR0), .Z(_03079__PTR1) );
  MUX2_X1 U22904 ( .A(1'b0), .B(_02169__PTR6), .S(P2_State_PTR0), .Z(_03079__PTR2) );
  MUX2_X1 U22905 ( .A(1'b1), .B(_02169__PTR12), .S(P2_State_PTR0), .Z(_03078__PTR0) );
  MUX2_X1 U22906 ( .A(1'b1), .B(_02169__PTR13), .S(P2_State_PTR0), .Z(_03078__PTR1) );
  MUX2_X1 U22907 ( .A(1'b0), .B(_02169__PTR14), .S(P2_State_PTR0), .Z(_03078__PTR2) );
  MUX2_X1 U22908 ( .A(_02169__PTR16), .B(_02169__PTR20), .S(P2_State_PTR0), .Z(_03078__PTR8) );
  MUX2_X1 U22909 ( .A(_02169__PTR17), .B(_02169__PTR21), .S(P2_State_PTR0), .Z(_03078__PTR9) );
  MUX2_X1 U22910 ( .A(_02169__PTR18), .B(_02169__PTR22), .S(P2_State_PTR0), .Z(_03078__PTR10) );
  MUX2_X1 U22911 ( .A(1'b0), .B(_02169__PTR28), .S(P2_State_PTR0), .Z(_03078__PTR16) );
  MUX2_X1 U22912 ( .A(P2_READY_n), .B(_02169__PTR29), .S(P2_State_PTR0), .Z(_03078__PTR17) );
  MUX2_X1 U22913 ( .A(1'b1), .B(_02169__PTR30), .S(P2_State_PTR0), .Z(_03078__PTR18) );
  MUX2_X1 U22914 ( .A(_03081__PTR0), .B(_03081__PTR256), .S(P2_State_PTR2), .Z(_02171__PTR0) );
  MUX2_X1 U22915 ( .A(_03081__PTR2), .B(_03081__PTR258), .S(P2_State_PTR2), .Z(_02171__PTR2) );
  MUX2_X1 U22916 ( .A(_03081__PTR3), .B(_03081__PTR259), .S(P2_State_PTR2), .Z(_02171__PTR3) );
  MUX2_X1 U22917 ( .A(_03081__PTR4), .B(_03081__PTR260), .S(P2_State_PTR2), .Z(_02171__PTR4) );
  MUX2_X1 U22918 ( .A(_03081__PTR5), .B(_03081__PTR261), .S(P2_State_PTR2), .Z(_02171__PTR5) );
  MUX2_X1 U22919 ( .A(_03081__PTR6), .B(_03081__PTR262), .S(P2_State_PTR2), .Z(_02171__PTR6) );
  MUX2_X1 U22920 ( .A(_03081__PTR7), .B(_03081__PTR263), .S(P2_State_PTR2), .Z(_02171__PTR7) );
  MUX2_X1 U22921 ( .A(_03081__PTR8), .B(_03081__PTR264), .S(P2_State_PTR2), .Z(_02171__PTR8) );
  MUX2_X1 U22922 ( .A(_03081__PTR9), .B(_03081__PTR265), .S(P2_State_PTR2), .Z(_02171__PTR9) );
  MUX2_X1 U22923 ( .A(_03081__PTR10), .B(_03081__PTR266), .S(P2_State_PTR2), .Z(_02171__PTR10) );
  MUX2_X1 U22924 ( .A(_03081__PTR11), .B(_03081__PTR267), .S(P2_State_PTR2), .Z(_02171__PTR11) );
  MUX2_X1 U22925 ( .A(_03081__PTR12), .B(_03081__PTR268), .S(P2_State_PTR2), .Z(_02171__PTR12) );
  MUX2_X1 U22926 ( .A(_03081__PTR13), .B(_03081__PTR269), .S(P2_State_PTR2), .Z(_02171__PTR13) );
  MUX2_X1 U22927 ( .A(_03081__PTR14), .B(_03081__PTR270), .S(P2_State_PTR2), .Z(_02171__PTR14) );
  MUX2_X1 U22928 ( .A(_03081__PTR15), .B(_03081__PTR271), .S(P2_State_PTR2), .Z(_02171__PTR15) );
  MUX2_X1 U22929 ( .A(_03081__PTR16), .B(_03081__PTR272), .S(P2_State_PTR2), .Z(_02171__PTR16) );
  MUX2_X1 U22930 ( .A(_03081__PTR17), .B(_03081__PTR273), .S(P2_State_PTR2), .Z(_02171__PTR17) );
  MUX2_X1 U22931 ( .A(_03081__PTR18), .B(_03081__PTR274), .S(P2_State_PTR2), .Z(_02171__PTR18) );
  MUX2_X1 U22932 ( .A(_03081__PTR19), .B(_03081__PTR275), .S(P2_State_PTR2), .Z(_02171__PTR19) );
  MUX2_X1 U22933 ( .A(_03081__PTR20), .B(_03081__PTR276), .S(P2_State_PTR2), .Z(_02171__PTR20) );
  MUX2_X1 U22934 ( .A(_03081__PTR21), .B(_03081__PTR277), .S(P2_State_PTR2), .Z(_02171__PTR21) );
  MUX2_X1 U22935 ( .A(_03081__PTR22), .B(_03081__PTR278), .S(P2_State_PTR2), .Z(_02171__PTR22) );
  MUX2_X1 U22936 ( .A(_03081__PTR23), .B(_03081__PTR279), .S(P2_State_PTR2), .Z(_02171__PTR23) );
  MUX2_X1 U22937 ( .A(_03081__PTR24), .B(_03081__PTR280), .S(P2_State_PTR2), .Z(_02171__PTR24) );
  MUX2_X1 U22938 ( .A(_03081__PTR25), .B(_03081__PTR281), .S(P2_State_PTR2), .Z(_02171__PTR25) );
  MUX2_X1 U22939 ( .A(_03081__PTR26), .B(_03081__PTR282), .S(P2_State_PTR2), .Z(_02171__PTR26) );
  MUX2_X1 U22940 ( .A(_03081__PTR27), .B(_03081__PTR283), .S(P2_State_PTR2), .Z(_02171__PTR27) );
  MUX2_X1 U22941 ( .A(_03081__PTR28), .B(_03081__PTR284), .S(P2_State_PTR2), .Z(_02171__PTR28) );
  MUX2_X1 U22942 ( .A(_03081__PTR29), .B(_03081__PTR285), .S(P2_State_PTR2), .Z(_02171__PTR29) );
  MUX2_X1 U22943 ( .A(_03081__PTR30), .B(_03081__PTR286), .S(P2_State_PTR2), .Z(_02171__PTR30) );
  MUX2_X1 U22944 ( .A(_03081__PTR32), .B(_03081__PTR288), .S(P2_State_PTR2), .Z(_02171__PTR32) );
  MUX2_X1 U22945 ( .A(_03001__PTR6), .B(_03080__PTR128), .S(P2_State_PTR1), .Z(_03081__PTR0) );
  MUX2_X1 U22946 ( .A(_03080__PTR258), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR2) );
  MUX2_X1 U22947 ( .A(_03080__PTR259), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR3) );
  MUX2_X1 U22948 ( .A(_03080__PTR260), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR4) );
  MUX2_X1 U22949 ( .A(_03080__PTR261), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR5) );
  MUX2_X1 U22950 ( .A(_03080__PTR262), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR6) );
  MUX2_X1 U22951 ( .A(_03080__PTR263), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR7) );
  MUX2_X1 U22952 ( .A(_03080__PTR264), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR8) );
  MUX2_X1 U22953 ( .A(_03080__PTR265), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR9) );
  MUX2_X1 U22954 ( .A(_03080__PTR266), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR10) );
  MUX2_X1 U22955 ( .A(_03080__PTR267), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR11) );
  MUX2_X1 U22956 ( .A(_03080__PTR268), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR12) );
  MUX2_X1 U22957 ( .A(_03080__PTR269), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR13) );
  MUX2_X1 U22958 ( .A(_03080__PTR270), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR14) );
  MUX2_X1 U22959 ( .A(_03080__PTR271), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR15) );
  MUX2_X1 U22960 ( .A(_03080__PTR272), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR16) );
  MUX2_X1 U22961 ( .A(_03080__PTR273), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR17) );
  MUX2_X1 U22962 ( .A(_03080__PTR274), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR18) );
  MUX2_X1 U22963 ( .A(_03080__PTR275), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR19) );
  MUX2_X1 U22964 ( .A(_03080__PTR276), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR20) );
  MUX2_X1 U22965 ( .A(_03080__PTR277), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR21) );
  MUX2_X1 U22966 ( .A(_03080__PTR278), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR22) );
  MUX2_X1 U22967 ( .A(_03080__PTR279), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR23) );
  MUX2_X1 U22968 ( .A(_03080__PTR280), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR24) );
  MUX2_X1 U22969 ( .A(_03080__PTR281), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR25) );
  MUX2_X1 U22970 ( .A(_03080__PTR282), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR26) );
  MUX2_X1 U22971 ( .A(_03080__PTR283), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR27) );
  MUX2_X1 U22972 ( .A(_03080__PTR284), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR28) );
  MUX2_X1 U22973 ( .A(_03080__PTR285), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR29) );
  MUX2_X1 U22974 ( .A(_03080__PTR286), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR30) );
  MUX2_X1 U22975 ( .A(_03080__PTR288), .B(_03080__PTR160), .S(P2_State_PTR1), .Z(_03081__PTR32) );
  MUX2_X1 U22976 ( .A(_03080__PTR256), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR256) );
  MUX2_X1 U22977 ( .A(_03080__PTR258), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR258) );
  MUX2_X1 U22978 ( .A(_03080__PTR259), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR259) );
  MUX2_X1 U22979 ( .A(_03080__PTR260), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR260) );
  MUX2_X1 U22980 ( .A(_03080__PTR261), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR261) );
  MUX2_X1 U22981 ( .A(_03080__PTR262), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR262) );
  MUX2_X1 U22982 ( .A(_03080__PTR263), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR263) );
  MUX2_X1 U22983 ( .A(_03080__PTR264), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR264) );
  MUX2_X1 U22984 ( .A(_03080__PTR265), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR265) );
  MUX2_X1 U22985 ( .A(_03080__PTR266), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR266) );
  MUX2_X1 U22986 ( .A(_03080__PTR267), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR267) );
  MUX2_X1 U22987 ( .A(_03080__PTR268), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR268) );
  MUX2_X1 U22988 ( .A(_03080__PTR269), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR269) );
  MUX2_X1 U22989 ( .A(_03080__PTR270), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR270) );
  MUX2_X1 U22990 ( .A(_03080__PTR271), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR271) );
  MUX2_X1 U22991 ( .A(_03080__PTR272), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR272) );
  MUX2_X1 U22992 ( .A(_03080__PTR273), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR273) );
  MUX2_X1 U22993 ( .A(_03080__PTR274), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR274) );
  MUX2_X1 U22994 ( .A(_03080__PTR275), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR275) );
  MUX2_X1 U22995 ( .A(_03080__PTR276), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR276) );
  MUX2_X1 U22996 ( .A(_03080__PTR277), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR277) );
  MUX2_X1 U22997 ( .A(_03080__PTR278), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR278) );
  MUX2_X1 U22998 ( .A(_03080__PTR279), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR279) );
  MUX2_X1 U22999 ( .A(_03080__PTR280), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR280) );
  MUX2_X1 U23000 ( .A(_03080__PTR281), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR281) );
  MUX2_X1 U23001 ( .A(_03080__PTR282), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR282) );
  MUX2_X1 U23002 ( .A(_03080__PTR283), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR283) );
  MUX2_X1 U23003 ( .A(_03080__PTR284), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR284) );
  MUX2_X1 U23004 ( .A(_03080__PTR285), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR285) );
  MUX2_X1 U23005 ( .A(_03080__PTR286), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR286) );
  MUX2_X1 U23006 ( .A(_03080__PTR288), .B(1'b0), .S(P2_State_PTR1), .Z(_03081__PTR288) );
  MUX2_X1 U23007 ( .A(1'b0), .B(_01878__PTR256), .S(P2_State_PTR0), .Z(_03080__PTR128) );
  MUX2_X1 U23008 ( .A(1'b0), .B(1'b0), .S(P2_State_PTR0), .Z(_03080__PTR160) );
  MUX2_X1 U23009 ( .A(_01878__PTR256), .B(1'b0), .S(P2_State_PTR0), .Z(_03080__PTR256) );
  MUX2_X1 U23010 ( .A(1'b0), .B(P2_DataWidth_PTR2), .S(P2_State_PTR0), .Z(_03080__PTR258) );
  MUX2_X1 U23011 ( .A(1'b0), .B(P2_DataWidth_PTR3), .S(P2_State_PTR0), .Z(_03080__PTR259) );
  MUX2_X1 U23012 ( .A(1'b0), .B(P2_DataWidth_PTR4), .S(P2_State_PTR0), .Z(_03080__PTR260) );
  MUX2_X1 U23013 ( .A(1'b0), .B(P2_DataWidth_PTR5), .S(P2_State_PTR0), .Z(_03080__PTR261) );
  MUX2_X1 U23014 ( .A(1'b0), .B(P2_DataWidth_PTR6), .S(P2_State_PTR0), .Z(_03080__PTR262) );
  MUX2_X1 U23015 ( .A(1'b0), .B(P2_DataWidth_PTR7), .S(P2_State_PTR0), .Z(_03080__PTR263) );
  MUX2_X1 U23016 ( .A(1'b0), .B(P2_DataWidth_PTR8), .S(P2_State_PTR0), .Z(_03080__PTR264) );
  MUX2_X1 U23017 ( .A(1'b0), .B(P2_DataWidth_PTR9), .S(P2_State_PTR0), .Z(_03080__PTR265) );
  MUX2_X1 U23018 ( .A(1'b0), .B(P2_DataWidth_PTR10), .S(P2_State_PTR0), .Z(_03080__PTR266) );
  MUX2_X1 U23019 ( .A(1'b0), .B(P2_DataWidth_PTR11), .S(P2_State_PTR0), .Z(_03080__PTR267) );
  MUX2_X1 U23020 ( .A(1'b0), .B(P2_DataWidth_PTR12), .S(P2_State_PTR0), .Z(_03080__PTR268) );
  MUX2_X1 U23021 ( .A(1'b0), .B(P2_DataWidth_PTR13), .S(P2_State_PTR0), .Z(_03080__PTR269) );
  MUX2_X1 U23022 ( .A(1'b0), .B(P2_DataWidth_PTR14), .S(P2_State_PTR0), .Z(_03080__PTR270) );
  MUX2_X1 U23023 ( .A(1'b0), .B(P2_DataWidth_PTR15), .S(P2_State_PTR0), .Z(_03080__PTR271) );
  MUX2_X1 U23024 ( .A(1'b0), .B(P2_DataWidth_PTR16), .S(P2_State_PTR0), .Z(_03080__PTR272) );
  MUX2_X1 U23025 ( .A(1'b0), .B(P2_DataWidth_PTR17), .S(P2_State_PTR0), .Z(_03080__PTR273) );
  MUX2_X1 U23026 ( .A(1'b0), .B(P2_DataWidth_PTR18), .S(P2_State_PTR0), .Z(_03080__PTR274) );
  MUX2_X1 U23027 ( .A(1'b0), .B(P2_DataWidth_PTR19), .S(P2_State_PTR0), .Z(_03080__PTR275) );
  MUX2_X1 U23028 ( .A(1'b0), .B(P2_DataWidth_PTR20), .S(P2_State_PTR0), .Z(_03080__PTR276) );
  MUX2_X1 U23029 ( .A(1'b0), .B(P2_DataWidth_PTR21), .S(P2_State_PTR0), .Z(_03080__PTR277) );
  MUX2_X1 U23030 ( .A(1'b0), .B(P2_DataWidth_PTR22), .S(P2_State_PTR0), .Z(_03080__PTR278) );
  MUX2_X1 U23031 ( .A(1'b0), .B(P2_DataWidth_PTR23), .S(P2_State_PTR0), .Z(_03080__PTR279) );
  MUX2_X1 U23032 ( .A(1'b0), .B(P2_DataWidth_PTR24), .S(P2_State_PTR0), .Z(_03080__PTR280) );
  MUX2_X1 U23033 ( .A(1'b0), .B(P2_DataWidth_PTR25), .S(P2_State_PTR0), .Z(_03080__PTR281) );
  MUX2_X1 U23034 ( .A(1'b0), .B(P2_DataWidth_PTR26), .S(P2_State_PTR0), .Z(_03080__PTR282) );
  MUX2_X1 U23035 ( .A(1'b0), .B(P2_DataWidth_PTR27), .S(P2_State_PTR0), .Z(_03080__PTR283) );
  MUX2_X1 U23036 ( .A(1'b0), .B(P2_DataWidth_PTR28), .S(P2_State_PTR0), .Z(_03080__PTR284) );
  MUX2_X1 U23037 ( .A(1'b0), .B(P2_DataWidth_PTR29), .S(P2_State_PTR0), .Z(_03080__PTR285) );
  MUX2_X1 U23038 ( .A(1'b0), .B(P2_DataWidth_PTR30), .S(P2_State_PTR0), .Z(_03080__PTR286) );
  MUX2_X1 U23039 ( .A(1'b0), .B(P2_DataWidth_PTR31), .S(P2_State_PTR0), .Z(_03080__PTR288) );
  MUX2_X1 U23040 ( .A(_03083__PTR0), .B(_03083__PTR128), .S(P2_State_PTR2), .Z(_02173__PTR0) );
  MUX2_X1 U23041 ( .A(_03083__PTR1), .B(_03083__PTR129), .S(P2_State_PTR2), .Z(_02173__PTR1) );
  MUX2_X1 U23042 ( .A(_03083__PTR2), .B(_03083__PTR130), .S(P2_State_PTR2), .Z(_02173__PTR2) );
  MUX2_X1 U23043 ( .A(_03083__PTR3), .B(_03083__PTR131), .S(P2_State_PTR2), .Z(_02173__PTR3) );
  MUX2_X1 U23044 ( .A(_03083__PTR4), .B(_03083__PTR132), .S(P2_State_PTR2), .Z(_02173__PTR4) );
  MUX2_X1 U23045 ( .A(_03083__PTR5), .B(_03083__PTR133), .S(P2_State_PTR2), .Z(_02173__PTR5) );
  MUX2_X1 U23046 ( .A(_03083__PTR6), .B(_03083__PTR134), .S(P2_State_PTR2), .Z(_02173__PTR6) );
  MUX2_X1 U23047 ( .A(_03083__PTR7), .B(_03083__PTR135), .S(P2_State_PTR2), .Z(_02173__PTR7) );
  MUX2_X1 U23048 ( .A(_03083__PTR8), .B(_03083__PTR136), .S(P2_State_PTR2), .Z(_02173__PTR8) );
  MUX2_X1 U23049 ( .A(_03083__PTR9), .B(_03083__PTR137), .S(P2_State_PTR2), .Z(_02173__PTR9) );
  MUX2_X1 U23050 ( .A(_03083__PTR10), .B(_03083__PTR138), .S(P2_State_PTR2), .Z(_02173__PTR10) );
  MUX2_X1 U23051 ( .A(_03083__PTR11), .B(_03083__PTR139), .S(P2_State_PTR2), .Z(_02173__PTR11) );
  MUX2_X1 U23052 ( .A(_03083__PTR12), .B(_03083__PTR140), .S(P2_State_PTR2), .Z(_02173__PTR12) );
  MUX2_X1 U23053 ( .A(_03083__PTR13), .B(_03083__PTR141), .S(P2_State_PTR2), .Z(_02173__PTR13) );
  MUX2_X1 U23054 ( .A(_03083__PTR14), .B(_03083__PTR142), .S(P2_State_PTR2), .Z(_02173__PTR14) );
  MUX2_X1 U23055 ( .A(_03083__PTR15), .B(_03083__PTR143), .S(P2_State_PTR2), .Z(_02173__PTR15) );
  MUX2_X1 U23056 ( .A(_03083__PTR16), .B(_03083__PTR144), .S(P2_State_PTR2), .Z(_02173__PTR16) );
  MUX2_X1 U23057 ( .A(_03083__PTR17), .B(_03083__PTR145), .S(P2_State_PTR2), .Z(_02173__PTR17) );
  MUX2_X1 U23058 ( .A(_03083__PTR18), .B(_03083__PTR146), .S(P2_State_PTR2), .Z(_02173__PTR18) );
  MUX2_X1 U23059 ( .A(_03083__PTR19), .B(_03083__PTR147), .S(P2_State_PTR2), .Z(_02173__PTR19) );
  MUX2_X1 U23060 ( .A(_03083__PTR20), .B(_03083__PTR148), .S(P2_State_PTR2), .Z(_02173__PTR20) );
  MUX2_X1 U23061 ( .A(_03083__PTR21), .B(_03083__PTR149), .S(P2_State_PTR2), .Z(_02173__PTR21) );
  MUX2_X1 U23062 ( .A(_03083__PTR22), .B(_03083__PTR150), .S(P2_State_PTR2), .Z(_02173__PTR22) );
  MUX2_X1 U23063 ( .A(_03083__PTR23), .B(_03083__PTR151), .S(P2_State_PTR2), .Z(_02173__PTR23) );
  MUX2_X1 U23064 ( .A(_03083__PTR24), .B(_03083__PTR152), .S(P2_State_PTR2), .Z(_02173__PTR24) );
  MUX2_X1 U23065 ( .A(_03083__PTR25), .B(_03083__PTR153), .S(P2_State_PTR2), .Z(_02173__PTR25) );
  MUX2_X1 U23066 ( .A(_03083__PTR26), .B(_03083__PTR154), .S(P2_State_PTR2), .Z(_02173__PTR26) );
  MUX2_X1 U23067 ( .A(_03083__PTR27), .B(_03083__PTR155), .S(P2_State_PTR2), .Z(_02173__PTR27) );
  MUX2_X1 U23068 ( .A(_03083__PTR28), .B(_03083__PTR156), .S(P2_State_PTR2), .Z(_02173__PTR28) );
  MUX2_X1 U23069 ( .A(_03083__PTR29), .B(_03083__PTR157), .S(P2_State_PTR2), .Z(_02173__PTR29) );
  MUX2_X1 U23070 ( .A(1'b0), .B(_03082__PTR64), .S(P2_State_PTR1), .Z(_03083__PTR0) );
  MUX2_X1 U23071 ( .A(1'b0), .B(_03082__PTR65), .S(P2_State_PTR1), .Z(_03083__PTR1) );
  MUX2_X1 U23072 ( .A(1'b0), .B(_03082__PTR66), .S(P2_State_PTR1), .Z(_03083__PTR2) );
  MUX2_X1 U23073 ( .A(1'b0), .B(_03082__PTR67), .S(P2_State_PTR1), .Z(_03083__PTR3) );
  MUX2_X1 U23074 ( .A(1'b0), .B(_03082__PTR68), .S(P2_State_PTR1), .Z(_03083__PTR4) );
  MUX2_X1 U23075 ( .A(1'b0), .B(_03082__PTR69), .S(P2_State_PTR1), .Z(_03083__PTR5) );
  MUX2_X1 U23076 ( .A(1'b0), .B(_03082__PTR70), .S(P2_State_PTR1), .Z(_03083__PTR6) );
  MUX2_X1 U23077 ( .A(1'b0), .B(_03082__PTR71), .S(P2_State_PTR1), .Z(_03083__PTR7) );
  MUX2_X1 U23078 ( .A(1'b0), .B(_03082__PTR72), .S(P2_State_PTR1), .Z(_03083__PTR8) );
  MUX2_X1 U23079 ( .A(1'b0), .B(_03082__PTR73), .S(P2_State_PTR1), .Z(_03083__PTR9) );
  MUX2_X1 U23080 ( .A(1'b0), .B(_03082__PTR74), .S(P2_State_PTR1), .Z(_03083__PTR10) );
  MUX2_X1 U23081 ( .A(1'b0), .B(_03082__PTR75), .S(P2_State_PTR1), .Z(_03083__PTR11) );
  MUX2_X1 U23082 ( .A(1'b0), .B(_03082__PTR76), .S(P2_State_PTR1), .Z(_03083__PTR12) );
  MUX2_X1 U23083 ( .A(1'b0), .B(_03082__PTR77), .S(P2_State_PTR1), .Z(_03083__PTR13) );
  MUX2_X1 U23084 ( .A(1'b0), .B(_03082__PTR78), .S(P2_State_PTR1), .Z(_03083__PTR14) );
  MUX2_X1 U23085 ( .A(1'b0), .B(_03082__PTR79), .S(P2_State_PTR1), .Z(_03083__PTR15) );
  MUX2_X1 U23086 ( .A(1'b0), .B(_03082__PTR80), .S(P2_State_PTR1), .Z(_03083__PTR16) );
  MUX2_X1 U23087 ( .A(1'b0), .B(_03082__PTR81), .S(P2_State_PTR1), .Z(_03083__PTR17) );
  MUX2_X1 U23088 ( .A(1'b0), .B(_03082__PTR82), .S(P2_State_PTR1), .Z(_03083__PTR18) );
  MUX2_X1 U23089 ( .A(1'b0), .B(_03082__PTR83), .S(P2_State_PTR1), .Z(_03083__PTR19) );
  MUX2_X1 U23090 ( .A(1'b0), .B(_03082__PTR84), .S(P2_State_PTR1), .Z(_03083__PTR20) );
  MUX2_X1 U23091 ( .A(1'b0), .B(_03082__PTR85), .S(P2_State_PTR1), .Z(_03083__PTR21) );
  MUX2_X1 U23092 ( .A(1'b0), .B(_03082__PTR86), .S(P2_State_PTR1), .Z(_03083__PTR22) );
  MUX2_X1 U23093 ( .A(1'b0), .B(_03082__PTR87), .S(P2_State_PTR1), .Z(_03083__PTR23) );
  MUX2_X1 U23094 ( .A(1'b0), .B(_03082__PTR88), .S(P2_State_PTR1), .Z(_03083__PTR24) );
  MUX2_X1 U23095 ( .A(1'b0), .B(_03082__PTR89), .S(P2_State_PTR1), .Z(_03083__PTR25) );
  MUX2_X1 U23096 ( .A(1'b0), .B(_03082__PTR90), .S(P2_State_PTR1), .Z(_03083__PTR26) );
  MUX2_X1 U23097 ( .A(1'b0), .B(_03082__PTR91), .S(P2_State_PTR1), .Z(_03083__PTR27) );
  MUX2_X1 U23098 ( .A(1'b0), .B(_03082__PTR92), .S(P2_State_PTR1), .Z(_03083__PTR28) );
  MUX2_X1 U23099 ( .A(1'b0), .B(_03082__PTR93), .S(P2_State_PTR1), .Z(_03083__PTR29) );
  MUX2_X1 U23100 ( .A(1'b0), .B(_03082__PTR192), .S(P2_State_PTR1), .Z(_03083__PTR128) );
  MUX2_X1 U23101 ( .A(1'b0), .B(_03082__PTR193), .S(P2_State_PTR1), .Z(_03083__PTR129) );
  MUX2_X1 U23102 ( .A(1'b0), .B(_03082__PTR194), .S(P2_State_PTR1), .Z(_03083__PTR130) );
  MUX2_X1 U23103 ( .A(1'b0), .B(_03082__PTR195), .S(P2_State_PTR1), .Z(_03083__PTR131) );
  MUX2_X1 U23104 ( .A(1'b0), .B(_03082__PTR196), .S(P2_State_PTR1), .Z(_03083__PTR132) );
  MUX2_X1 U23105 ( .A(1'b0), .B(_03082__PTR197), .S(P2_State_PTR1), .Z(_03083__PTR133) );
  MUX2_X1 U23106 ( .A(1'b0), .B(_03082__PTR198), .S(P2_State_PTR1), .Z(_03083__PTR134) );
  MUX2_X1 U23107 ( .A(1'b0), .B(_03082__PTR199), .S(P2_State_PTR1), .Z(_03083__PTR135) );
  MUX2_X1 U23108 ( .A(1'b0), .B(_03082__PTR200), .S(P2_State_PTR1), .Z(_03083__PTR136) );
  MUX2_X1 U23109 ( .A(1'b0), .B(_03082__PTR201), .S(P2_State_PTR1), .Z(_03083__PTR137) );
  MUX2_X1 U23110 ( .A(1'b0), .B(_03082__PTR202), .S(P2_State_PTR1), .Z(_03083__PTR138) );
  MUX2_X1 U23111 ( .A(1'b0), .B(_03082__PTR203), .S(P2_State_PTR1), .Z(_03083__PTR139) );
  MUX2_X1 U23112 ( .A(1'b0), .B(_03082__PTR204), .S(P2_State_PTR1), .Z(_03083__PTR140) );
  MUX2_X1 U23113 ( .A(1'b0), .B(_03082__PTR205), .S(P2_State_PTR1), .Z(_03083__PTR141) );
  MUX2_X1 U23114 ( .A(1'b0), .B(_03082__PTR206), .S(P2_State_PTR1), .Z(_03083__PTR142) );
  MUX2_X1 U23115 ( .A(1'b0), .B(_03082__PTR207), .S(P2_State_PTR1), .Z(_03083__PTR143) );
  MUX2_X1 U23116 ( .A(1'b0), .B(_03082__PTR208), .S(P2_State_PTR1), .Z(_03083__PTR144) );
  MUX2_X1 U23117 ( .A(1'b0), .B(_03082__PTR209), .S(P2_State_PTR1), .Z(_03083__PTR145) );
  MUX2_X1 U23118 ( .A(1'b0), .B(_03082__PTR210), .S(P2_State_PTR1), .Z(_03083__PTR146) );
  MUX2_X1 U23119 ( .A(1'b0), .B(_03082__PTR211), .S(P2_State_PTR1), .Z(_03083__PTR147) );
  MUX2_X1 U23120 ( .A(1'b0), .B(_03082__PTR212), .S(P2_State_PTR1), .Z(_03083__PTR148) );
  MUX2_X1 U23121 ( .A(1'b0), .B(_03082__PTR213), .S(P2_State_PTR1), .Z(_03083__PTR149) );
  MUX2_X1 U23122 ( .A(1'b0), .B(_03082__PTR214), .S(P2_State_PTR1), .Z(_03083__PTR150) );
  MUX2_X1 U23123 ( .A(1'b0), .B(_03082__PTR215), .S(P2_State_PTR1), .Z(_03083__PTR151) );
  MUX2_X1 U23124 ( .A(1'b0), .B(_03082__PTR216), .S(P2_State_PTR1), .Z(_03083__PTR152) );
  MUX2_X1 U23125 ( .A(1'b0), .B(_03082__PTR217), .S(P2_State_PTR1), .Z(_03083__PTR153) );
  MUX2_X1 U23126 ( .A(1'b0), .B(_03082__PTR218), .S(P2_State_PTR1), .Z(_03083__PTR154) );
  MUX2_X1 U23127 ( .A(1'b0), .B(_03082__PTR219), .S(P2_State_PTR1), .Z(_03083__PTR155) );
  MUX2_X1 U23128 ( .A(1'b0), .B(_03082__PTR220), .S(P2_State_PTR1), .Z(_03083__PTR156) );
  MUX2_X1 U23129 ( .A(1'b0), .B(_03082__PTR221), .S(P2_State_PTR1), .Z(_03083__PTR157) );
  MUX2_X1 U23130 ( .A(_02172__PTR64), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR64) );
  MUX2_X1 U23131 ( .A(_02172__PTR65), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR65) );
  MUX2_X1 U23132 ( .A(_02172__PTR66), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR66) );
  MUX2_X1 U23133 ( .A(_02172__PTR67), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR67) );
  MUX2_X1 U23134 ( .A(_02172__PTR68), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR68) );
  MUX2_X1 U23135 ( .A(_02172__PTR69), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR69) );
  MUX2_X1 U23136 ( .A(_02172__PTR70), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR70) );
  MUX2_X1 U23137 ( .A(_02172__PTR71), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR71) );
  MUX2_X1 U23138 ( .A(_02172__PTR72), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR72) );
  MUX2_X1 U23139 ( .A(_02172__PTR73), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR73) );
  MUX2_X1 U23140 ( .A(_02172__PTR74), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR74) );
  MUX2_X1 U23141 ( .A(_02172__PTR75), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR75) );
  MUX2_X1 U23142 ( .A(_02172__PTR76), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR76) );
  MUX2_X1 U23143 ( .A(_02172__PTR77), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR77) );
  MUX2_X1 U23144 ( .A(_02172__PTR78), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR78) );
  MUX2_X1 U23145 ( .A(_02172__PTR79), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR79) );
  MUX2_X1 U23146 ( .A(_02172__PTR80), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR80) );
  MUX2_X1 U23147 ( .A(_02172__PTR81), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR81) );
  MUX2_X1 U23148 ( .A(_02172__PTR82), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR82) );
  MUX2_X1 U23149 ( .A(_02172__PTR83), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR83) );
  MUX2_X1 U23150 ( .A(_02172__PTR84), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR84) );
  MUX2_X1 U23151 ( .A(_02172__PTR85), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR85) );
  MUX2_X1 U23152 ( .A(_02172__PTR86), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR86) );
  MUX2_X1 U23153 ( .A(_02172__PTR87), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR87) );
  MUX2_X1 U23154 ( .A(_02172__PTR88), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR88) );
  MUX2_X1 U23155 ( .A(_02172__PTR89), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR89) );
  MUX2_X1 U23156 ( .A(_02172__PTR90), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR90) );
  MUX2_X1 U23157 ( .A(_02172__PTR91), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR91) );
  MUX2_X1 U23158 ( .A(_02172__PTR92), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR92) );
  MUX2_X1 U23159 ( .A(_02172__PTR93), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR93) );
  MUX2_X1 U23160 ( .A(_02172__PTR192), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR192) );
  MUX2_X1 U23161 ( .A(_02172__PTR193), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR193) );
  MUX2_X1 U23162 ( .A(_02172__PTR194), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR194) );
  MUX2_X1 U23163 ( .A(_02172__PTR195), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR195) );
  MUX2_X1 U23164 ( .A(_02172__PTR196), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR196) );
  MUX2_X1 U23165 ( .A(_02172__PTR197), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR197) );
  MUX2_X1 U23166 ( .A(_02172__PTR198), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR198) );
  MUX2_X1 U23167 ( .A(_02172__PTR199), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR199) );
  MUX2_X1 U23168 ( .A(_02172__PTR200), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR200) );
  MUX2_X1 U23169 ( .A(_02172__PTR201), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR201) );
  MUX2_X1 U23170 ( .A(_02172__PTR202), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR202) );
  MUX2_X1 U23171 ( .A(_02172__PTR203), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR203) );
  MUX2_X1 U23172 ( .A(_02172__PTR204), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR204) );
  MUX2_X1 U23173 ( .A(_02172__PTR205), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR205) );
  MUX2_X1 U23174 ( .A(_02172__PTR206), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR206) );
  MUX2_X1 U23175 ( .A(_02172__PTR207), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR207) );
  MUX2_X1 U23176 ( .A(_02172__PTR208), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR208) );
  MUX2_X1 U23177 ( .A(_02172__PTR209), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR209) );
  MUX2_X1 U23178 ( .A(_02172__PTR210), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR210) );
  MUX2_X1 U23179 ( .A(_02172__PTR211), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR211) );
  MUX2_X1 U23180 ( .A(_02172__PTR212), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR212) );
  MUX2_X1 U23181 ( .A(_02172__PTR213), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR213) );
  MUX2_X1 U23182 ( .A(_02172__PTR214), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR214) );
  MUX2_X1 U23183 ( .A(_02172__PTR215), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR215) );
  MUX2_X1 U23184 ( .A(_02172__PTR216), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR216) );
  MUX2_X1 U23185 ( .A(_02172__PTR217), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR217) );
  MUX2_X1 U23186 ( .A(_02172__PTR218), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR218) );
  MUX2_X1 U23187 ( .A(_02172__PTR219), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR219) );
  MUX2_X1 U23188 ( .A(_02172__PTR220), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR220) );
  MUX2_X1 U23189 ( .A(_02172__PTR221), .B(1'b0), .S(P2_State_PTR0), .Z(_03082__PTR221) );
  INV_X1 U23190 ( .A(P2_rEIP_PTR0), .ZN(_03084__PTR43) );
  MUX2_X1 U23191 ( .A(1'b0), .B(P2_rEIP_PTR0), .S(P2_rEIP_PTR1), .Z(_02174__PTR2) );
  MUX2_X1 U23192 ( .A(_03084__PTR43), .B(P2_rEIP_PTR0), .S(P2_rEIP_PTR1), .Z(_02174__PTR6) );
  MUX2_X1 U23193 ( .A(P2_rEIP_PTR0), .B(1'b1), .S(P2_rEIP_PTR1), .Z(_02174__PTR8) );
  MUX2_X1 U23194 ( .A(_03084__PTR43), .B(1'b1), .S(P2_rEIP_PTR1), .Z(_02174__PTR9) );
  MUX2_X1 U23195 ( .A(1'b1), .B(P2_rEIP_PTR0), .S(P2_rEIP_PTR1), .Z(_02174__PTR10) );
  MUX2_X1 U23196 ( .A(1'b1), .B(_03084__PTR43), .S(P2_rEIP_PTR1), .Z(_02174__PTR11) );
  MUX2_X1 U23197 ( .A(_03087__PTR0), .B(_03087__PTR64), .S(P2_P1_InstQueueRd_Addr_PTR3), .Z(_02175__PTR0) );
  MUX2_X1 U23198 ( .A(_03087__PTR1), .B(_03087__PTR65), .S(P2_P1_InstQueueRd_Addr_PTR3), .Z(_02175__PTR1) );
  MUX2_X1 U23199 ( .A(_03087__PTR2), .B(_03087__PTR66), .S(P2_P1_InstQueueRd_Addr_PTR3), .Z(_02175__PTR2) );
  MUX2_X1 U23200 ( .A(_03087__PTR3), .B(_03087__PTR67), .S(P2_P1_InstQueueRd_Addr_PTR3), .Z(_02175__PTR3) );
  MUX2_X1 U23201 ( .A(_03087__PTR4), .B(_03087__PTR68), .S(P2_P1_InstQueueRd_Addr_PTR3), .Z(_02175__PTR4) );
  MUX2_X1 U23202 ( .A(_03087__PTR5), .B(_03087__PTR69), .S(P2_P1_InstQueueRd_Addr_PTR3), .Z(_02175__PTR5) );
  MUX2_X1 U23203 ( .A(_03087__PTR6), .B(_03087__PTR70), .S(P2_P1_InstQueueRd_Addr_PTR3), .Z(_02175__PTR6) );
  MUX2_X1 U23204 ( .A(_03087__PTR7), .B(_03087__PTR71), .S(P2_P1_InstQueueRd_Addr_PTR3), .Z(_02175__PTR7) );
  MUX2_X1 U23205 ( .A(_03086__PTR0), .B(_03086__PTR32), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR0) );
  MUX2_X1 U23206 ( .A(_03086__PTR1), .B(_03086__PTR33), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR1) );
  MUX2_X1 U23207 ( .A(_03086__PTR2), .B(_03086__PTR34), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR2) );
  MUX2_X1 U23208 ( .A(_03086__PTR3), .B(_03086__PTR35), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR3) );
  MUX2_X1 U23209 ( .A(_03086__PTR4), .B(_03086__PTR36), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR4) );
  MUX2_X1 U23210 ( .A(_03086__PTR5), .B(_03086__PTR37), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR5) );
  MUX2_X1 U23211 ( .A(_03086__PTR6), .B(_03086__PTR38), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR6) );
  MUX2_X1 U23212 ( .A(_03086__PTR7), .B(_03086__PTR39), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR7) );
  MUX2_X1 U23213 ( .A(_03086__PTR64), .B(_03086__PTR96), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR64) );
  MUX2_X1 U23214 ( .A(_03086__PTR65), .B(_03086__PTR97), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR65) );
  MUX2_X1 U23215 ( .A(_03086__PTR66), .B(_03086__PTR98), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR66) );
  MUX2_X1 U23216 ( .A(_03086__PTR67), .B(_03086__PTR99), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR67) );
  MUX2_X1 U23217 ( .A(_03086__PTR68), .B(_03086__PTR100), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR68) );
  MUX2_X1 U23218 ( .A(_03086__PTR69), .B(_03086__PTR101), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR69) );
  MUX2_X1 U23219 ( .A(_03086__PTR70), .B(_03086__PTR102), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR70) );
  MUX2_X1 U23220 ( .A(_03086__PTR71), .B(_03086__PTR103), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03087__PTR71) );
  MUX2_X1 U23221 ( .A(_03085__PTR0), .B(_03085__PTR16), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR0) );
  MUX2_X1 U23222 ( .A(_03085__PTR1), .B(_03085__PTR17), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR1) );
  MUX2_X1 U23223 ( .A(_03085__PTR2), .B(_03085__PTR18), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR2) );
  MUX2_X1 U23224 ( .A(_03085__PTR3), .B(_03085__PTR19), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR3) );
  MUX2_X1 U23225 ( .A(_03085__PTR4), .B(_03085__PTR20), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR4) );
  MUX2_X1 U23226 ( .A(_03085__PTR5), .B(_03085__PTR21), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR5) );
  MUX2_X1 U23227 ( .A(_03085__PTR6), .B(_03085__PTR22), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR6) );
  MUX2_X1 U23228 ( .A(_03085__PTR7), .B(_03085__PTR23), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR7) );
  MUX2_X1 U23229 ( .A(_03085__PTR32), .B(_03085__PTR48), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR32) );
  MUX2_X1 U23230 ( .A(_03085__PTR33), .B(_03085__PTR49), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR33) );
  MUX2_X1 U23231 ( .A(_03085__PTR34), .B(_03085__PTR50), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR34) );
  MUX2_X1 U23232 ( .A(_03085__PTR35), .B(_03085__PTR51), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR35) );
  MUX2_X1 U23233 ( .A(_03085__PTR36), .B(_03085__PTR52), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR36) );
  MUX2_X1 U23234 ( .A(_03085__PTR37), .B(_03085__PTR53), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR37) );
  MUX2_X1 U23235 ( .A(_03085__PTR38), .B(_03085__PTR54), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR38) );
  MUX2_X1 U23236 ( .A(_03085__PTR39), .B(_03085__PTR55), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR39) );
  MUX2_X1 U23237 ( .A(_03085__PTR64), .B(_03085__PTR80), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR64) );
  MUX2_X1 U23238 ( .A(_03085__PTR65), .B(_03085__PTR81), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR65) );
  MUX2_X1 U23239 ( .A(_03085__PTR66), .B(_03085__PTR82), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR66) );
  MUX2_X1 U23240 ( .A(_03085__PTR67), .B(_03085__PTR83), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR67) );
  MUX2_X1 U23241 ( .A(_03085__PTR68), .B(_03085__PTR84), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR68) );
  MUX2_X1 U23242 ( .A(_03085__PTR69), .B(_03085__PTR85), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR69) );
  MUX2_X1 U23243 ( .A(_03085__PTR70), .B(_03085__PTR86), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR70) );
  MUX2_X1 U23244 ( .A(_03085__PTR71), .B(_03085__PTR87), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR71) );
  MUX2_X1 U23245 ( .A(_03085__PTR96), .B(_03085__PTR112), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR96) );
  MUX2_X1 U23246 ( .A(_03085__PTR97), .B(_03085__PTR113), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR97) );
  MUX2_X1 U23247 ( .A(_03085__PTR98), .B(_03085__PTR114), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR98) );
  MUX2_X1 U23248 ( .A(_03085__PTR99), .B(_03085__PTR115), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR99) );
  MUX2_X1 U23249 ( .A(_03085__PTR100), .B(_03085__PTR116), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR100) );
  MUX2_X1 U23250 ( .A(_03085__PTR101), .B(_03085__PTR117), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR101) );
  MUX2_X1 U23251 ( .A(_03085__PTR102), .B(_03085__PTR118), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR102) );
  MUX2_X1 U23252 ( .A(_03085__PTR103), .B(_03085__PTR119), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03086__PTR103) );
  MUX2_X1 U23253 ( .A(P2_P1_InstQueue_PTR0_PTR0), .B(P2_P1_InstQueue_PTR1_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR0) );
  MUX2_X1 U23254 ( .A(P2_P1_InstQueue_PTR0_PTR1), .B(P2_P1_InstQueue_PTR1_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR1) );
  MUX2_X1 U23255 ( .A(P2_P1_InstQueue_PTR0_PTR2), .B(P2_P1_InstQueue_PTR1_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR2) );
  MUX2_X1 U23256 ( .A(P2_P1_InstQueue_PTR0_PTR3), .B(P2_P1_InstQueue_PTR1_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR3) );
  MUX2_X1 U23257 ( .A(P2_P1_InstQueue_PTR0_PTR4), .B(P2_P1_InstQueue_PTR1_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR4) );
  MUX2_X1 U23258 ( .A(P2_P1_InstQueue_PTR0_PTR5), .B(P2_P1_InstQueue_PTR1_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR5) );
  MUX2_X1 U23259 ( .A(P2_P1_InstQueue_PTR0_PTR6), .B(P2_P1_InstQueue_PTR1_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR6) );
  MUX2_X1 U23260 ( .A(P2_P1_InstQueue_PTR0_PTR7), .B(P2_P1_InstQueue_PTR1_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR7) );
  MUX2_X1 U23261 ( .A(P2_P1_InstQueue_PTR2_PTR0), .B(P2_P1_InstQueue_PTR3_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR16) );
  MUX2_X1 U23262 ( .A(P2_P1_InstQueue_PTR2_PTR1), .B(P2_P1_InstQueue_PTR3_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR17) );
  MUX2_X1 U23263 ( .A(P2_P1_InstQueue_PTR2_PTR2), .B(P2_P1_InstQueue_PTR3_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR18) );
  MUX2_X1 U23264 ( .A(P2_P1_InstQueue_PTR2_PTR3), .B(P2_P1_InstQueue_PTR3_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR19) );
  MUX2_X1 U23265 ( .A(P2_P1_InstQueue_PTR2_PTR4), .B(P2_P1_InstQueue_PTR3_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR20) );
  MUX2_X1 U23266 ( .A(P2_P1_InstQueue_PTR2_PTR5), .B(P2_P1_InstQueue_PTR3_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR21) );
  MUX2_X1 U23267 ( .A(P2_P1_InstQueue_PTR2_PTR6), .B(P2_P1_InstQueue_PTR3_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR22) );
  MUX2_X1 U23268 ( .A(P2_P1_InstQueue_PTR2_PTR7), .B(P2_P1_InstQueue_PTR3_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR23) );
  MUX2_X1 U23269 ( .A(P2_P1_InstQueue_PTR4_PTR0), .B(P2_P1_InstQueue_PTR5_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR32) );
  MUX2_X1 U23270 ( .A(P2_P1_InstQueue_PTR4_PTR1), .B(P2_P1_InstQueue_PTR5_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR33) );
  MUX2_X1 U23271 ( .A(P2_P1_InstQueue_PTR4_PTR2), .B(P2_P1_InstQueue_PTR5_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR34) );
  MUX2_X1 U23272 ( .A(P2_P1_InstQueue_PTR4_PTR3), .B(P2_P1_InstQueue_PTR5_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR35) );
  MUX2_X1 U23273 ( .A(P2_P1_InstQueue_PTR4_PTR4), .B(P2_P1_InstQueue_PTR5_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR36) );
  MUX2_X1 U23274 ( .A(P2_P1_InstQueue_PTR4_PTR5), .B(P2_P1_InstQueue_PTR5_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR37) );
  MUX2_X1 U23275 ( .A(P2_P1_InstQueue_PTR4_PTR6), .B(P2_P1_InstQueue_PTR5_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR38) );
  MUX2_X1 U23276 ( .A(P2_P1_InstQueue_PTR4_PTR7), .B(P2_P1_InstQueue_PTR5_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR39) );
  MUX2_X1 U23277 ( .A(P2_P1_InstQueue_PTR6_PTR0), .B(P2_P1_InstQueue_PTR7_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR48) );
  MUX2_X1 U23278 ( .A(P2_P1_InstQueue_PTR6_PTR1), .B(P2_P1_InstQueue_PTR7_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR49) );
  MUX2_X1 U23279 ( .A(P2_P1_InstQueue_PTR6_PTR2), .B(P2_P1_InstQueue_PTR7_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR50) );
  MUX2_X1 U23280 ( .A(P2_P1_InstQueue_PTR6_PTR3), .B(P2_P1_InstQueue_PTR7_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR51) );
  MUX2_X1 U23281 ( .A(P2_P1_InstQueue_PTR6_PTR4), .B(P2_P1_InstQueue_PTR7_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR52) );
  MUX2_X1 U23282 ( .A(P2_P1_InstQueue_PTR6_PTR5), .B(P2_P1_InstQueue_PTR7_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR53) );
  MUX2_X1 U23283 ( .A(P2_P1_InstQueue_PTR6_PTR6), .B(P2_P1_InstQueue_PTR7_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR54) );
  MUX2_X1 U23284 ( .A(P2_P1_InstQueue_PTR6_PTR7), .B(P2_P1_InstQueue_PTR7_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR55) );
  MUX2_X1 U23285 ( .A(P2_P1_InstQueue_PTR8_PTR0), .B(P2_P1_InstQueue_PTR9_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR64) );
  MUX2_X1 U23286 ( .A(P2_P1_InstQueue_PTR8_PTR1), .B(P2_P1_InstQueue_PTR9_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR65) );
  MUX2_X1 U23287 ( .A(P2_P1_InstQueue_PTR8_PTR2), .B(P2_P1_InstQueue_PTR9_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR66) );
  MUX2_X1 U23288 ( .A(P2_P1_InstQueue_PTR8_PTR3), .B(P2_P1_InstQueue_PTR9_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR67) );
  MUX2_X1 U23289 ( .A(P2_P1_InstQueue_PTR8_PTR4), .B(P2_P1_InstQueue_PTR9_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR68) );
  MUX2_X1 U23290 ( .A(P2_P1_InstQueue_PTR8_PTR5), .B(P2_P1_InstQueue_PTR9_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR69) );
  MUX2_X1 U23291 ( .A(P2_P1_InstQueue_PTR8_PTR6), .B(P2_P1_InstQueue_PTR9_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR70) );
  MUX2_X1 U23292 ( .A(P2_P1_InstQueue_PTR8_PTR7), .B(P2_P1_InstQueue_PTR9_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR71) );
  MUX2_X1 U23293 ( .A(P2_P1_InstQueue_PTR10_PTR0), .B(P2_P1_InstQueue_PTR11_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR80) );
  MUX2_X1 U23294 ( .A(P2_P1_InstQueue_PTR10_PTR1), .B(P2_P1_InstQueue_PTR11_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR81) );
  MUX2_X1 U23295 ( .A(P2_P1_InstQueue_PTR10_PTR2), .B(P2_P1_InstQueue_PTR11_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR82) );
  MUX2_X1 U23296 ( .A(P2_P1_InstQueue_PTR10_PTR3), .B(P2_P1_InstQueue_PTR11_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR83) );
  MUX2_X1 U23297 ( .A(P2_P1_InstQueue_PTR10_PTR4), .B(P2_P1_InstQueue_PTR11_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR84) );
  MUX2_X1 U23298 ( .A(P2_P1_InstQueue_PTR10_PTR5), .B(P2_P1_InstQueue_PTR11_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR85) );
  MUX2_X1 U23299 ( .A(P2_P1_InstQueue_PTR10_PTR6), .B(P2_P1_InstQueue_PTR11_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR86) );
  MUX2_X1 U23300 ( .A(P2_P1_InstQueue_PTR10_PTR7), .B(P2_P1_InstQueue_PTR11_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR87) );
  MUX2_X1 U23301 ( .A(P2_P1_InstQueue_PTR12_PTR0), .B(P2_P1_InstQueue_PTR13_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR96) );
  MUX2_X1 U23302 ( .A(P2_P1_InstQueue_PTR12_PTR1), .B(P2_P1_InstQueue_PTR13_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR97) );
  MUX2_X1 U23303 ( .A(P2_P1_InstQueue_PTR12_PTR2), .B(P2_P1_InstQueue_PTR13_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR98) );
  MUX2_X1 U23304 ( .A(P2_P1_InstQueue_PTR12_PTR3), .B(P2_P1_InstQueue_PTR13_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR99) );
  MUX2_X1 U23305 ( .A(P2_P1_InstQueue_PTR12_PTR4), .B(P2_P1_InstQueue_PTR13_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR100) );
  MUX2_X1 U23306 ( .A(P2_P1_InstQueue_PTR12_PTR5), .B(P2_P1_InstQueue_PTR13_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR101) );
  MUX2_X1 U23307 ( .A(P2_P1_InstQueue_PTR12_PTR6), .B(P2_P1_InstQueue_PTR13_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR102) );
  MUX2_X1 U23308 ( .A(P2_P1_InstQueue_PTR12_PTR7), .B(P2_P1_InstQueue_PTR13_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR103) );
  MUX2_X1 U23309 ( .A(P2_P1_InstQueue_PTR14_PTR0), .B(P2_P1_InstQueue_PTR15_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR112) );
  MUX2_X1 U23310 ( .A(P2_P1_InstQueue_PTR14_PTR1), .B(P2_P1_InstQueue_PTR15_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR113) );
  MUX2_X1 U23311 ( .A(P2_P1_InstQueue_PTR14_PTR2), .B(P2_P1_InstQueue_PTR15_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR114) );
  MUX2_X1 U23312 ( .A(P2_P1_InstQueue_PTR14_PTR3), .B(P2_P1_InstQueue_PTR15_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR115) );
  MUX2_X1 U23313 ( .A(P2_P1_InstQueue_PTR14_PTR4), .B(P2_P1_InstQueue_PTR15_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR116) );
  MUX2_X1 U23314 ( .A(P2_P1_InstQueue_PTR14_PTR5), .B(P2_P1_InstQueue_PTR15_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR117) );
  MUX2_X1 U23315 ( .A(P2_P1_InstQueue_PTR14_PTR6), .B(P2_P1_InstQueue_PTR15_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR118) );
  MUX2_X1 U23316 ( .A(P2_P1_InstQueue_PTR14_PTR7), .B(P2_P1_InstQueue_PTR15_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03085__PTR119) );
  MUX2_X1 U23317 ( .A(_03090__PTR0), .B(_03090__PTR64), .S(_02176__PTR6), .Z(_02177__PTR0) );
  MUX2_X1 U23318 ( .A(_03090__PTR1), .B(_03090__PTR65), .S(_02176__PTR6), .Z(_02177__PTR1) );
  MUX2_X1 U23319 ( .A(_03090__PTR2), .B(_03090__PTR66), .S(_02176__PTR6), .Z(_02177__PTR2) );
  MUX2_X1 U23320 ( .A(_03090__PTR3), .B(_03090__PTR67), .S(_02176__PTR6), .Z(_02177__PTR3) );
  MUX2_X1 U23321 ( .A(_03090__PTR4), .B(_03090__PTR68), .S(_02176__PTR6), .Z(_02177__PTR4) );
  MUX2_X1 U23322 ( .A(_03090__PTR5), .B(_03090__PTR69), .S(_02176__PTR6), .Z(_02177__PTR5) );
  MUX2_X1 U23323 ( .A(_03090__PTR6), .B(_03090__PTR70), .S(_02176__PTR6), .Z(_02177__PTR6) );
  MUX2_X1 U23324 ( .A(_03090__PTR7), .B(_03090__PTR71), .S(_02176__PTR6), .Z(_02177__PTR7) );
  MUX2_X1 U23325 ( .A(_03089__PTR0), .B(_03089__PTR32), .S(_02176__PTR5), .Z(_03090__PTR0) );
  MUX2_X1 U23326 ( .A(_03089__PTR1), .B(_03089__PTR33), .S(_02176__PTR5), .Z(_03090__PTR1) );
  MUX2_X1 U23327 ( .A(_03089__PTR2), .B(_03089__PTR34), .S(_02176__PTR5), .Z(_03090__PTR2) );
  MUX2_X1 U23328 ( .A(_03089__PTR3), .B(_03089__PTR35), .S(_02176__PTR5), .Z(_03090__PTR3) );
  MUX2_X1 U23329 ( .A(_03089__PTR4), .B(_03089__PTR36), .S(_02176__PTR5), .Z(_03090__PTR4) );
  MUX2_X1 U23330 ( .A(_03089__PTR5), .B(_03089__PTR37), .S(_02176__PTR5), .Z(_03090__PTR5) );
  MUX2_X1 U23331 ( .A(_03089__PTR6), .B(_03089__PTR38), .S(_02176__PTR5), .Z(_03090__PTR6) );
  MUX2_X1 U23332 ( .A(_03089__PTR7), .B(_03089__PTR39), .S(_02176__PTR5), .Z(_03090__PTR7) );
  MUX2_X1 U23333 ( .A(_03089__PTR64), .B(_03089__PTR96), .S(_02176__PTR5), .Z(_03090__PTR64) );
  MUX2_X1 U23334 ( .A(_03089__PTR65), .B(_03089__PTR97), .S(_02176__PTR5), .Z(_03090__PTR65) );
  MUX2_X1 U23335 ( .A(_03089__PTR66), .B(_03089__PTR98), .S(_02176__PTR5), .Z(_03090__PTR66) );
  MUX2_X1 U23336 ( .A(_03089__PTR67), .B(_03089__PTR99), .S(_02176__PTR5), .Z(_03090__PTR67) );
  MUX2_X1 U23337 ( .A(_03089__PTR68), .B(_03089__PTR100), .S(_02176__PTR5), .Z(_03090__PTR68) );
  MUX2_X1 U23338 ( .A(_03089__PTR69), .B(_03089__PTR101), .S(_02176__PTR5), .Z(_03090__PTR69) );
  MUX2_X1 U23339 ( .A(_03089__PTR70), .B(_03089__PTR102), .S(_02176__PTR5), .Z(_03090__PTR70) );
  MUX2_X1 U23340 ( .A(_03089__PTR71), .B(_03089__PTR103), .S(_02176__PTR5), .Z(_03090__PTR71) );
  MUX2_X1 U23341 ( .A(_03088__PTR0), .B(_03088__PTR16), .S(_02176__PTR4), .Z(_03089__PTR0) );
  MUX2_X1 U23342 ( .A(_03088__PTR1), .B(_03088__PTR17), .S(_02176__PTR4), .Z(_03089__PTR1) );
  MUX2_X1 U23343 ( .A(_03088__PTR2), .B(_03088__PTR18), .S(_02176__PTR4), .Z(_03089__PTR2) );
  MUX2_X1 U23344 ( .A(_03088__PTR3), .B(_03088__PTR19), .S(_02176__PTR4), .Z(_03089__PTR3) );
  MUX2_X1 U23345 ( .A(_03088__PTR4), .B(_03088__PTR20), .S(_02176__PTR4), .Z(_03089__PTR4) );
  MUX2_X1 U23346 ( .A(_03088__PTR5), .B(_03088__PTR21), .S(_02176__PTR4), .Z(_03089__PTR5) );
  MUX2_X1 U23347 ( .A(_03088__PTR6), .B(_03088__PTR22), .S(_02176__PTR4), .Z(_03089__PTR6) );
  MUX2_X1 U23348 ( .A(_03088__PTR7), .B(_03088__PTR23), .S(_02176__PTR4), .Z(_03089__PTR7) );
  MUX2_X1 U23349 ( .A(_03088__PTR32), .B(_03088__PTR48), .S(_02176__PTR4), .Z(_03089__PTR32) );
  MUX2_X1 U23350 ( .A(_03088__PTR33), .B(_03088__PTR49), .S(_02176__PTR4), .Z(_03089__PTR33) );
  MUX2_X1 U23351 ( .A(_03088__PTR34), .B(_03088__PTR50), .S(_02176__PTR4), .Z(_03089__PTR34) );
  MUX2_X1 U23352 ( .A(_03088__PTR35), .B(_03088__PTR51), .S(_02176__PTR4), .Z(_03089__PTR35) );
  MUX2_X1 U23353 ( .A(_03088__PTR36), .B(_03088__PTR52), .S(_02176__PTR4), .Z(_03089__PTR36) );
  MUX2_X1 U23354 ( .A(_03088__PTR37), .B(_03088__PTR53), .S(_02176__PTR4), .Z(_03089__PTR37) );
  MUX2_X1 U23355 ( .A(_03088__PTR38), .B(_03088__PTR54), .S(_02176__PTR4), .Z(_03089__PTR38) );
  MUX2_X1 U23356 ( .A(_03088__PTR39), .B(_03088__PTR55), .S(_02176__PTR4), .Z(_03089__PTR39) );
  MUX2_X1 U23357 ( .A(_03088__PTR64), .B(_03088__PTR80), .S(_02176__PTR4), .Z(_03089__PTR64) );
  MUX2_X1 U23358 ( .A(_03088__PTR65), .B(_03088__PTR81), .S(_02176__PTR4), .Z(_03089__PTR65) );
  MUX2_X1 U23359 ( .A(_03088__PTR66), .B(_03088__PTR82), .S(_02176__PTR4), .Z(_03089__PTR66) );
  MUX2_X1 U23360 ( .A(_03088__PTR67), .B(_03088__PTR83), .S(_02176__PTR4), .Z(_03089__PTR67) );
  MUX2_X1 U23361 ( .A(_03088__PTR68), .B(_03088__PTR84), .S(_02176__PTR4), .Z(_03089__PTR68) );
  MUX2_X1 U23362 ( .A(_03088__PTR69), .B(_03088__PTR85), .S(_02176__PTR4), .Z(_03089__PTR69) );
  MUX2_X1 U23363 ( .A(_03088__PTR70), .B(_03088__PTR86), .S(_02176__PTR4), .Z(_03089__PTR70) );
  MUX2_X1 U23364 ( .A(_03088__PTR71), .B(_03088__PTR87), .S(_02176__PTR4), .Z(_03089__PTR71) );
  MUX2_X1 U23365 ( .A(_03088__PTR96), .B(_03088__PTR112), .S(_02176__PTR4), .Z(_03089__PTR96) );
  MUX2_X1 U23366 ( .A(_03088__PTR97), .B(_03088__PTR113), .S(_02176__PTR4), .Z(_03089__PTR97) );
  MUX2_X1 U23367 ( .A(_03088__PTR98), .B(_03088__PTR114), .S(_02176__PTR4), .Z(_03089__PTR98) );
  MUX2_X1 U23368 ( .A(_03088__PTR99), .B(_03088__PTR115), .S(_02176__PTR4), .Z(_03089__PTR99) );
  MUX2_X1 U23369 ( .A(_03088__PTR100), .B(_03088__PTR116), .S(_02176__PTR4), .Z(_03089__PTR100) );
  MUX2_X1 U23370 ( .A(_03088__PTR101), .B(_03088__PTR117), .S(_02176__PTR4), .Z(_03089__PTR101) );
  MUX2_X1 U23371 ( .A(_03088__PTR102), .B(_03088__PTR118), .S(_02176__PTR4), .Z(_03089__PTR102) );
  MUX2_X1 U23372 ( .A(_03088__PTR103), .B(_03088__PTR119), .S(_02176__PTR4), .Z(_03089__PTR103) );
  MUX2_X1 U23373 ( .A(P2_P1_InstQueue_PTR1_PTR0), .B(P2_P1_InstQueue_PTR0_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR0) );
  MUX2_X1 U23374 ( .A(P2_P1_InstQueue_PTR1_PTR1), .B(P2_P1_InstQueue_PTR0_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR1) );
  MUX2_X1 U23375 ( .A(P2_P1_InstQueue_PTR1_PTR2), .B(P2_P1_InstQueue_PTR0_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR2) );
  MUX2_X1 U23376 ( .A(P2_P1_InstQueue_PTR1_PTR3), .B(P2_P1_InstQueue_PTR0_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR3) );
  MUX2_X1 U23377 ( .A(P2_P1_InstQueue_PTR1_PTR4), .B(P2_P1_InstQueue_PTR0_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR4) );
  MUX2_X1 U23378 ( .A(P2_P1_InstQueue_PTR1_PTR5), .B(P2_P1_InstQueue_PTR0_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR5) );
  MUX2_X1 U23379 ( .A(P2_P1_InstQueue_PTR1_PTR6), .B(P2_P1_InstQueue_PTR0_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR6) );
  MUX2_X1 U23380 ( .A(P2_P1_InstQueue_PTR1_PTR7), .B(P2_P1_InstQueue_PTR0_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR7) );
  MUX2_X1 U23381 ( .A(P2_P1_InstQueue_PTR3_PTR0), .B(P2_P1_InstQueue_PTR2_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR16) );
  MUX2_X1 U23382 ( .A(P2_P1_InstQueue_PTR3_PTR1), .B(P2_P1_InstQueue_PTR2_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR17) );
  MUX2_X1 U23383 ( .A(P2_P1_InstQueue_PTR3_PTR2), .B(P2_P1_InstQueue_PTR2_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR18) );
  MUX2_X1 U23384 ( .A(P2_P1_InstQueue_PTR3_PTR3), .B(P2_P1_InstQueue_PTR2_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR19) );
  MUX2_X1 U23385 ( .A(P2_P1_InstQueue_PTR3_PTR4), .B(P2_P1_InstQueue_PTR2_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR20) );
  MUX2_X1 U23386 ( .A(P2_P1_InstQueue_PTR3_PTR5), .B(P2_P1_InstQueue_PTR2_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR21) );
  MUX2_X1 U23387 ( .A(P2_P1_InstQueue_PTR3_PTR6), .B(P2_P1_InstQueue_PTR2_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR22) );
  MUX2_X1 U23388 ( .A(P2_P1_InstQueue_PTR3_PTR7), .B(P2_P1_InstQueue_PTR2_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR23) );
  MUX2_X1 U23389 ( .A(P2_P1_InstQueue_PTR5_PTR0), .B(P2_P1_InstQueue_PTR4_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR32) );
  MUX2_X1 U23390 ( .A(P2_P1_InstQueue_PTR5_PTR1), .B(P2_P1_InstQueue_PTR4_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR33) );
  MUX2_X1 U23391 ( .A(P2_P1_InstQueue_PTR5_PTR2), .B(P2_P1_InstQueue_PTR4_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR34) );
  MUX2_X1 U23392 ( .A(P2_P1_InstQueue_PTR5_PTR3), .B(P2_P1_InstQueue_PTR4_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR35) );
  MUX2_X1 U23393 ( .A(P2_P1_InstQueue_PTR5_PTR4), .B(P2_P1_InstQueue_PTR4_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR36) );
  MUX2_X1 U23394 ( .A(P2_P1_InstQueue_PTR5_PTR5), .B(P2_P1_InstQueue_PTR4_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR37) );
  MUX2_X1 U23395 ( .A(P2_P1_InstQueue_PTR5_PTR6), .B(P2_P1_InstQueue_PTR4_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR38) );
  MUX2_X1 U23396 ( .A(P2_P1_InstQueue_PTR5_PTR7), .B(P2_P1_InstQueue_PTR4_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR39) );
  MUX2_X1 U23397 ( .A(P2_P1_InstQueue_PTR7_PTR0), .B(P2_P1_InstQueue_PTR6_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR48) );
  MUX2_X1 U23398 ( .A(P2_P1_InstQueue_PTR7_PTR1), .B(P2_P1_InstQueue_PTR6_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR49) );
  MUX2_X1 U23399 ( .A(P2_P1_InstQueue_PTR7_PTR2), .B(P2_P1_InstQueue_PTR6_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR50) );
  MUX2_X1 U23400 ( .A(P2_P1_InstQueue_PTR7_PTR3), .B(P2_P1_InstQueue_PTR6_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR51) );
  MUX2_X1 U23401 ( .A(P2_P1_InstQueue_PTR7_PTR4), .B(P2_P1_InstQueue_PTR6_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR52) );
  MUX2_X1 U23402 ( .A(P2_P1_InstQueue_PTR7_PTR5), .B(P2_P1_InstQueue_PTR6_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR53) );
  MUX2_X1 U23403 ( .A(P2_P1_InstQueue_PTR7_PTR6), .B(P2_P1_InstQueue_PTR6_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR54) );
  MUX2_X1 U23404 ( .A(P2_P1_InstQueue_PTR7_PTR7), .B(P2_P1_InstQueue_PTR6_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR55) );
  MUX2_X1 U23405 ( .A(P2_P1_InstQueue_PTR9_PTR0), .B(P2_P1_InstQueue_PTR8_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR64) );
  MUX2_X1 U23406 ( .A(P2_P1_InstQueue_PTR9_PTR1), .B(P2_P1_InstQueue_PTR8_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR65) );
  MUX2_X1 U23407 ( .A(P2_P1_InstQueue_PTR9_PTR2), .B(P2_P1_InstQueue_PTR8_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR66) );
  MUX2_X1 U23408 ( .A(P2_P1_InstQueue_PTR9_PTR3), .B(P2_P1_InstQueue_PTR8_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR67) );
  MUX2_X1 U23409 ( .A(P2_P1_InstQueue_PTR9_PTR4), .B(P2_P1_InstQueue_PTR8_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR68) );
  MUX2_X1 U23410 ( .A(P2_P1_InstQueue_PTR9_PTR5), .B(P2_P1_InstQueue_PTR8_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR69) );
  MUX2_X1 U23411 ( .A(P2_P1_InstQueue_PTR9_PTR6), .B(P2_P1_InstQueue_PTR8_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR70) );
  MUX2_X1 U23412 ( .A(P2_P1_InstQueue_PTR9_PTR7), .B(P2_P1_InstQueue_PTR8_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR71) );
  MUX2_X1 U23413 ( .A(P2_P1_InstQueue_PTR11_PTR0), .B(P2_P1_InstQueue_PTR10_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR80) );
  MUX2_X1 U23414 ( .A(P2_P1_InstQueue_PTR11_PTR1), .B(P2_P1_InstQueue_PTR10_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR81) );
  MUX2_X1 U23415 ( .A(P2_P1_InstQueue_PTR11_PTR2), .B(P2_P1_InstQueue_PTR10_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR82) );
  MUX2_X1 U23416 ( .A(P2_P1_InstQueue_PTR11_PTR3), .B(P2_P1_InstQueue_PTR10_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR83) );
  MUX2_X1 U23417 ( .A(P2_P1_InstQueue_PTR11_PTR4), .B(P2_P1_InstQueue_PTR10_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR84) );
  MUX2_X1 U23418 ( .A(P2_P1_InstQueue_PTR11_PTR5), .B(P2_P1_InstQueue_PTR10_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR85) );
  MUX2_X1 U23419 ( .A(P2_P1_InstQueue_PTR11_PTR6), .B(P2_P1_InstQueue_PTR10_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR86) );
  MUX2_X1 U23420 ( .A(P2_P1_InstQueue_PTR11_PTR7), .B(P2_P1_InstQueue_PTR10_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR87) );
  MUX2_X1 U23421 ( .A(P2_P1_InstQueue_PTR13_PTR0), .B(P2_P1_InstQueue_PTR12_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR96) );
  MUX2_X1 U23422 ( .A(P2_P1_InstQueue_PTR13_PTR1), .B(P2_P1_InstQueue_PTR12_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR97) );
  MUX2_X1 U23423 ( .A(P2_P1_InstQueue_PTR13_PTR2), .B(P2_P1_InstQueue_PTR12_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR98) );
  MUX2_X1 U23424 ( .A(P2_P1_InstQueue_PTR13_PTR3), .B(P2_P1_InstQueue_PTR12_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR99) );
  MUX2_X1 U23425 ( .A(P2_P1_InstQueue_PTR13_PTR4), .B(P2_P1_InstQueue_PTR12_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR100) );
  MUX2_X1 U23426 ( .A(P2_P1_InstQueue_PTR13_PTR5), .B(P2_P1_InstQueue_PTR12_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR101) );
  MUX2_X1 U23427 ( .A(P2_P1_InstQueue_PTR13_PTR6), .B(P2_P1_InstQueue_PTR12_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR102) );
  MUX2_X1 U23428 ( .A(P2_P1_InstQueue_PTR13_PTR7), .B(P2_P1_InstQueue_PTR12_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR103) );
  MUX2_X1 U23429 ( .A(P2_P1_InstQueue_PTR15_PTR0), .B(P2_P1_InstQueue_PTR14_PTR0), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR112) );
  MUX2_X1 U23430 ( .A(P2_P1_InstQueue_PTR15_PTR1), .B(P2_P1_InstQueue_PTR14_PTR1), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR113) );
  MUX2_X1 U23431 ( .A(P2_P1_InstQueue_PTR15_PTR2), .B(P2_P1_InstQueue_PTR14_PTR2), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR114) );
  MUX2_X1 U23432 ( .A(P2_P1_InstQueue_PTR15_PTR3), .B(P2_P1_InstQueue_PTR14_PTR3), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR115) );
  MUX2_X1 U23433 ( .A(P2_P1_InstQueue_PTR15_PTR4), .B(P2_P1_InstQueue_PTR14_PTR4), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR116) );
  MUX2_X1 U23434 ( .A(P2_P1_InstQueue_PTR15_PTR5), .B(P2_P1_InstQueue_PTR14_PTR5), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR117) );
  MUX2_X1 U23435 ( .A(P2_P1_InstQueue_PTR15_PTR6), .B(P2_P1_InstQueue_PTR14_PTR6), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR118) );
  MUX2_X1 U23436 ( .A(P2_P1_InstQueue_PTR15_PTR7), .B(P2_P1_InstQueue_PTR14_PTR7), .S(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03088__PTR119) );
  MUX2_X1 U23437 ( .A(_03091__PTR0), .B(_03091__PTR64), .S(_02178__PTR6), .Z(_02179__PTR0) );
  MUX2_X1 U23438 ( .A(_03091__PTR1), .B(_03091__PTR65), .S(_02178__PTR6), .Z(_02179__PTR1) );
  MUX2_X1 U23439 ( .A(_03091__PTR2), .B(_03091__PTR66), .S(_02178__PTR6), .Z(_02179__PTR2) );
  MUX2_X1 U23440 ( .A(_03091__PTR3), .B(_03091__PTR67), .S(_02178__PTR6), .Z(_02179__PTR3) );
  MUX2_X1 U23441 ( .A(_03091__PTR4), .B(_03091__PTR68), .S(_02178__PTR6), .Z(_02179__PTR4) );
  MUX2_X1 U23442 ( .A(_03091__PTR5), .B(_03091__PTR69), .S(_02178__PTR6), .Z(_02179__PTR5) );
  MUX2_X1 U23443 ( .A(_03091__PTR6), .B(_03091__PTR70), .S(_02178__PTR6), .Z(_02179__PTR6) );
  MUX2_X1 U23444 ( .A(_03091__PTR7), .B(_03091__PTR71), .S(_02178__PTR6), .Z(_02179__PTR7) );
  MUX2_X1 U23445 ( .A(_03086__PTR32), .B(_03086__PTR0), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR0) );
  MUX2_X1 U23446 ( .A(_03086__PTR33), .B(_03086__PTR1), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR1) );
  MUX2_X1 U23447 ( .A(_03086__PTR34), .B(_03086__PTR2), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR2) );
  MUX2_X1 U23448 ( .A(_03086__PTR35), .B(_03086__PTR3), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR3) );
  MUX2_X1 U23449 ( .A(_03086__PTR36), .B(_03086__PTR4), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR4) );
  MUX2_X1 U23450 ( .A(_03086__PTR37), .B(_03086__PTR5), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR5) );
  MUX2_X1 U23451 ( .A(_03086__PTR38), .B(_03086__PTR6), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR6) );
  MUX2_X1 U23452 ( .A(_03086__PTR39), .B(_03086__PTR7), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR7) );
  MUX2_X1 U23453 ( .A(_03086__PTR96), .B(_03086__PTR64), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR64) );
  MUX2_X1 U23454 ( .A(_03086__PTR97), .B(_03086__PTR65), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR65) );
  MUX2_X1 U23455 ( .A(_03086__PTR98), .B(_03086__PTR66), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR66) );
  MUX2_X1 U23456 ( .A(_03086__PTR99), .B(_03086__PTR67), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR67) );
  MUX2_X1 U23457 ( .A(_03086__PTR100), .B(_03086__PTR68), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR68) );
  MUX2_X1 U23458 ( .A(_03086__PTR101), .B(_03086__PTR69), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR69) );
  MUX2_X1 U23459 ( .A(_03086__PTR102), .B(_03086__PTR70), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR70) );
  MUX2_X1 U23460 ( .A(_03086__PTR103), .B(_03086__PTR71), .S(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03091__PTR71) );
  MUX2_X1 U23461 ( .A(_03093__PTR0), .B(_03093__PTR64), .S(_02180__PTR6), .Z(_02181__PTR0) );
  MUX2_X1 U23462 ( .A(_03093__PTR1), .B(_03093__PTR65), .S(_02180__PTR6), .Z(_02181__PTR1) );
  MUX2_X1 U23463 ( .A(_03093__PTR2), .B(_03093__PTR66), .S(_02180__PTR6), .Z(_02181__PTR2) );
  MUX2_X1 U23464 ( .A(_03093__PTR3), .B(_03093__PTR67), .S(_02180__PTR6), .Z(_02181__PTR3) );
  MUX2_X1 U23465 ( .A(_03093__PTR4), .B(_03093__PTR68), .S(_02180__PTR6), .Z(_02181__PTR4) );
  MUX2_X1 U23466 ( .A(_03093__PTR5), .B(_03093__PTR69), .S(_02180__PTR6), .Z(_02181__PTR5) );
  MUX2_X1 U23467 ( .A(_03093__PTR6), .B(_03093__PTR70), .S(_02180__PTR6), .Z(_02181__PTR6) );
  MUX2_X1 U23468 ( .A(_03093__PTR7), .B(_03093__PTR71), .S(_02180__PTR6), .Z(_02181__PTR7) );
  MUX2_X1 U23469 ( .A(_03092__PTR0), .B(_03092__PTR32), .S(_02180__PTR5), .Z(_03093__PTR0) );
  MUX2_X1 U23470 ( .A(_03092__PTR1), .B(_03092__PTR33), .S(_02180__PTR5), .Z(_03093__PTR1) );
  MUX2_X1 U23471 ( .A(_03092__PTR2), .B(_03092__PTR34), .S(_02180__PTR5), .Z(_03093__PTR2) );
  MUX2_X1 U23472 ( .A(_03092__PTR3), .B(_03092__PTR35), .S(_02180__PTR5), .Z(_03093__PTR3) );
  MUX2_X1 U23473 ( .A(_03092__PTR4), .B(_03092__PTR36), .S(_02180__PTR5), .Z(_03093__PTR4) );
  MUX2_X1 U23474 ( .A(_03092__PTR5), .B(_03092__PTR37), .S(_02180__PTR5), .Z(_03093__PTR5) );
  MUX2_X1 U23475 ( .A(_03092__PTR6), .B(_03092__PTR38), .S(_02180__PTR5), .Z(_03093__PTR6) );
  MUX2_X1 U23476 ( .A(_03092__PTR7), .B(_03092__PTR39), .S(_02180__PTR5), .Z(_03093__PTR7) );
  MUX2_X1 U23477 ( .A(_03092__PTR64), .B(_03092__PTR96), .S(_02180__PTR5), .Z(_03093__PTR64) );
  MUX2_X1 U23478 ( .A(_03092__PTR65), .B(_03092__PTR97), .S(_02180__PTR5), .Z(_03093__PTR65) );
  MUX2_X1 U23479 ( .A(_03092__PTR66), .B(_03092__PTR98), .S(_02180__PTR5), .Z(_03093__PTR66) );
  MUX2_X1 U23480 ( .A(_03092__PTR67), .B(_03092__PTR99), .S(_02180__PTR5), .Z(_03093__PTR67) );
  MUX2_X1 U23481 ( .A(_03092__PTR68), .B(_03092__PTR100), .S(_02180__PTR5), .Z(_03093__PTR68) );
  MUX2_X1 U23482 ( .A(_03092__PTR69), .B(_03092__PTR101), .S(_02180__PTR5), .Z(_03093__PTR69) );
  MUX2_X1 U23483 ( .A(_03092__PTR70), .B(_03092__PTR102), .S(_02180__PTR5), .Z(_03093__PTR70) );
  MUX2_X1 U23484 ( .A(_03092__PTR71), .B(_03092__PTR103), .S(_02180__PTR5), .Z(_03093__PTR71) );
  MUX2_X1 U23485 ( .A(_03088__PTR0), .B(_03088__PTR16), .S(_02180__PTR4), .Z(_03092__PTR0) );
  MUX2_X1 U23486 ( .A(_03088__PTR1), .B(_03088__PTR17), .S(_02180__PTR4), .Z(_03092__PTR1) );
  MUX2_X1 U23487 ( .A(_03088__PTR2), .B(_03088__PTR18), .S(_02180__PTR4), .Z(_03092__PTR2) );
  MUX2_X1 U23488 ( .A(_03088__PTR3), .B(_03088__PTR19), .S(_02180__PTR4), .Z(_03092__PTR3) );
  MUX2_X1 U23489 ( .A(_03088__PTR4), .B(_03088__PTR20), .S(_02180__PTR4), .Z(_03092__PTR4) );
  MUX2_X1 U23490 ( .A(_03088__PTR5), .B(_03088__PTR21), .S(_02180__PTR4), .Z(_03092__PTR5) );
  MUX2_X1 U23491 ( .A(_03088__PTR6), .B(_03088__PTR22), .S(_02180__PTR4), .Z(_03092__PTR6) );
  MUX2_X1 U23492 ( .A(_03088__PTR7), .B(_03088__PTR23), .S(_02180__PTR4), .Z(_03092__PTR7) );
  MUX2_X1 U23493 ( .A(_03088__PTR32), .B(_03088__PTR48), .S(_02180__PTR4), .Z(_03092__PTR32) );
  MUX2_X1 U23494 ( .A(_03088__PTR33), .B(_03088__PTR49), .S(_02180__PTR4), .Z(_03092__PTR33) );
  MUX2_X1 U23495 ( .A(_03088__PTR34), .B(_03088__PTR50), .S(_02180__PTR4), .Z(_03092__PTR34) );
  MUX2_X1 U23496 ( .A(_03088__PTR35), .B(_03088__PTR51), .S(_02180__PTR4), .Z(_03092__PTR35) );
  MUX2_X1 U23497 ( .A(_03088__PTR36), .B(_03088__PTR52), .S(_02180__PTR4), .Z(_03092__PTR36) );
  MUX2_X1 U23498 ( .A(_03088__PTR37), .B(_03088__PTR53), .S(_02180__PTR4), .Z(_03092__PTR37) );
  MUX2_X1 U23499 ( .A(_03088__PTR38), .B(_03088__PTR54), .S(_02180__PTR4), .Z(_03092__PTR38) );
  MUX2_X1 U23500 ( .A(_03088__PTR39), .B(_03088__PTR55), .S(_02180__PTR4), .Z(_03092__PTR39) );
  MUX2_X1 U23501 ( .A(_03088__PTR64), .B(_03088__PTR80), .S(_02180__PTR4), .Z(_03092__PTR64) );
  MUX2_X1 U23502 ( .A(_03088__PTR65), .B(_03088__PTR81), .S(_02180__PTR4), .Z(_03092__PTR65) );
  MUX2_X1 U23503 ( .A(_03088__PTR66), .B(_03088__PTR82), .S(_02180__PTR4), .Z(_03092__PTR66) );
  MUX2_X1 U23504 ( .A(_03088__PTR67), .B(_03088__PTR83), .S(_02180__PTR4), .Z(_03092__PTR67) );
  MUX2_X1 U23505 ( .A(_03088__PTR68), .B(_03088__PTR84), .S(_02180__PTR4), .Z(_03092__PTR68) );
  MUX2_X1 U23506 ( .A(_03088__PTR69), .B(_03088__PTR85), .S(_02180__PTR4), .Z(_03092__PTR69) );
  MUX2_X1 U23507 ( .A(_03088__PTR70), .B(_03088__PTR86), .S(_02180__PTR4), .Z(_03092__PTR70) );
  MUX2_X1 U23508 ( .A(_03088__PTR71), .B(_03088__PTR87), .S(_02180__PTR4), .Z(_03092__PTR71) );
  MUX2_X1 U23509 ( .A(_03088__PTR96), .B(_03088__PTR112), .S(_02180__PTR4), .Z(_03092__PTR96) );
  MUX2_X1 U23510 ( .A(_03088__PTR97), .B(_03088__PTR113), .S(_02180__PTR4), .Z(_03092__PTR97) );
  MUX2_X1 U23511 ( .A(_03088__PTR98), .B(_03088__PTR114), .S(_02180__PTR4), .Z(_03092__PTR98) );
  MUX2_X1 U23512 ( .A(_03088__PTR99), .B(_03088__PTR115), .S(_02180__PTR4), .Z(_03092__PTR99) );
  MUX2_X1 U23513 ( .A(_03088__PTR100), .B(_03088__PTR116), .S(_02180__PTR4), .Z(_03092__PTR100) );
  MUX2_X1 U23514 ( .A(_03088__PTR101), .B(_03088__PTR117), .S(_02180__PTR4), .Z(_03092__PTR101) );
  MUX2_X1 U23515 ( .A(_03088__PTR102), .B(_03088__PTR118), .S(_02180__PTR4), .Z(_03092__PTR102) );
  MUX2_X1 U23516 ( .A(_03088__PTR103), .B(_03088__PTR119), .S(_02180__PTR4), .Z(_03092__PTR103) );
  MUX2_X1 U23517 ( .A(_03095__PTR0), .B(_03095__PTR64), .S(_02182__PTR6), .Z(_02183__PTR0) );
  MUX2_X1 U23518 ( .A(_03095__PTR1), .B(_03095__PTR65), .S(_02182__PTR6), .Z(_02183__PTR1) );
  MUX2_X1 U23519 ( .A(_03095__PTR2), .B(_03095__PTR66), .S(_02182__PTR6), .Z(_02183__PTR2) );
  MUX2_X1 U23520 ( .A(_03095__PTR3), .B(_03095__PTR67), .S(_02182__PTR6), .Z(_02183__PTR3) );
  MUX2_X1 U23521 ( .A(_03095__PTR4), .B(_03095__PTR68), .S(_02182__PTR6), .Z(_02183__PTR4) );
  MUX2_X1 U23522 ( .A(_03095__PTR5), .B(_03095__PTR69), .S(_02182__PTR6), .Z(_02183__PTR5) );
  MUX2_X1 U23523 ( .A(_03095__PTR6), .B(_03095__PTR70), .S(_02182__PTR6), .Z(_02183__PTR6) );
  MUX2_X1 U23524 ( .A(_03095__PTR7), .B(_03095__PTR71), .S(_02182__PTR6), .Z(_02183__PTR7) );
  MUX2_X1 U23525 ( .A(_03094__PTR0), .B(_03094__PTR32), .S(_02182__PTR5), .Z(_03095__PTR0) );
  MUX2_X1 U23526 ( .A(_03094__PTR1), .B(_03094__PTR33), .S(_02182__PTR5), .Z(_03095__PTR1) );
  MUX2_X1 U23527 ( .A(_03094__PTR2), .B(_03094__PTR34), .S(_02182__PTR5), .Z(_03095__PTR2) );
  MUX2_X1 U23528 ( .A(_03094__PTR3), .B(_03094__PTR35), .S(_02182__PTR5), .Z(_03095__PTR3) );
  MUX2_X1 U23529 ( .A(_03094__PTR4), .B(_03094__PTR36), .S(_02182__PTR5), .Z(_03095__PTR4) );
  MUX2_X1 U23530 ( .A(_03094__PTR5), .B(_03094__PTR37), .S(_02182__PTR5), .Z(_03095__PTR5) );
  MUX2_X1 U23531 ( .A(_03094__PTR6), .B(_03094__PTR38), .S(_02182__PTR5), .Z(_03095__PTR6) );
  MUX2_X1 U23532 ( .A(_03094__PTR7), .B(_03094__PTR39), .S(_02182__PTR5), .Z(_03095__PTR7) );
  MUX2_X1 U23533 ( .A(_03094__PTR64), .B(_03094__PTR96), .S(_02182__PTR5), .Z(_03095__PTR64) );
  MUX2_X1 U23534 ( .A(_03094__PTR65), .B(_03094__PTR97), .S(_02182__PTR5), .Z(_03095__PTR65) );
  MUX2_X1 U23535 ( .A(_03094__PTR66), .B(_03094__PTR98), .S(_02182__PTR5), .Z(_03095__PTR66) );
  MUX2_X1 U23536 ( .A(_03094__PTR67), .B(_03094__PTR99), .S(_02182__PTR5), .Z(_03095__PTR67) );
  MUX2_X1 U23537 ( .A(_03094__PTR68), .B(_03094__PTR100), .S(_02182__PTR5), .Z(_03095__PTR68) );
  MUX2_X1 U23538 ( .A(_03094__PTR69), .B(_03094__PTR101), .S(_02182__PTR5), .Z(_03095__PTR69) );
  MUX2_X1 U23539 ( .A(_03094__PTR70), .B(_03094__PTR102), .S(_02182__PTR5), .Z(_03095__PTR70) );
  MUX2_X1 U23540 ( .A(_03094__PTR71), .B(_03094__PTR103), .S(_02182__PTR5), .Z(_03095__PTR71) );
  MUX2_X1 U23541 ( .A(_03085__PTR16), .B(_03085__PTR0), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR0) );
  MUX2_X1 U23542 ( .A(_03085__PTR17), .B(_03085__PTR1), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR1) );
  MUX2_X1 U23543 ( .A(_03085__PTR18), .B(_03085__PTR2), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR2) );
  MUX2_X1 U23544 ( .A(_03085__PTR19), .B(_03085__PTR3), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR3) );
  MUX2_X1 U23545 ( .A(_03085__PTR20), .B(_03085__PTR4), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR4) );
  MUX2_X1 U23546 ( .A(_03085__PTR21), .B(_03085__PTR5), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR5) );
  MUX2_X1 U23547 ( .A(_03085__PTR22), .B(_03085__PTR6), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR6) );
  MUX2_X1 U23548 ( .A(_03085__PTR23), .B(_03085__PTR7), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR7) );
  MUX2_X1 U23549 ( .A(_03085__PTR48), .B(_03085__PTR32), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR32) );
  MUX2_X1 U23550 ( .A(_03085__PTR49), .B(_03085__PTR33), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR33) );
  MUX2_X1 U23551 ( .A(_03085__PTR50), .B(_03085__PTR34), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR34) );
  MUX2_X1 U23552 ( .A(_03085__PTR51), .B(_03085__PTR35), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR35) );
  MUX2_X1 U23553 ( .A(_03085__PTR52), .B(_03085__PTR36), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR36) );
  MUX2_X1 U23554 ( .A(_03085__PTR53), .B(_03085__PTR37), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR37) );
  MUX2_X1 U23555 ( .A(_03085__PTR54), .B(_03085__PTR38), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR38) );
  MUX2_X1 U23556 ( .A(_03085__PTR55), .B(_03085__PTR39), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR39) );
  MUX2_X1 U23557 ( .A(_03085__PTR80), .B(_03085__PTR64), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR64) );
  MUX2_X1 U23558 ( .A(_03085__PTR81), .B(_03085__PTR65), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR65) );
  MUX2_X1 U23559 ( .A(_03085__PTR82), .B(_03085__PTR66), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR66) );
  MUX2_X1 U23560 ( .A(_03085__PTR83), .B(_03085__PTR67), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR67) );
  MUX2_X1 U23561 ( .A(_03085__PTR84), .B(_03085__PTR68), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR68) );
  MUX2_X1 U23562 ( .A(_03085__PTR85), .B(_03085__PTR69), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR69) );
  MUX2_X1 U23563 ( .A(_03085__PTR86), .B(_03085__PTR70), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR70) );
  MUX2_X1 U23564 ( .A(_03085__PTR87), .B(_03085__PTR71), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR71) );
  MUX2_X1 U23565 ( .A(_03085__PTR112), .B(_03085__PTR96), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR96) );
  MUX2_X1 U23566 ( .A(_03085__PTR113), .B(_03085__PTR97), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR97) );
  MUX2_X1 U23567 ( .A(_03085__PTR114), .B(_03085__PTR98), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR98) );
  MUX2_X1 U23568 ( .A(_03085__PTR115), .B(_03085__PTR99), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR99) );
  MUX2_X1 U23569 ( .A(_03085__PTR116), .B(_03085__PTR100), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR100) );
  MUX2_X1 U23570 ( .A(_03085__PTR117), .B(_03085__PTR101), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR101) );
  MUX2_X1 U23571 ( .A(_03085__PTR118), .B(_03085__PTR102), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR102) );
  MUX2_X1 U23572 ( .A(_03085__PTR119), .B(_03085__PTR103), .S(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03094__PTR103) );
  MUX2_X1 U23573 ( .A(_03097__PTR0), .B(_03097__PTR128), .S(P2_P1_State2_PTR2), .Z(_03098__PTR0) );
  MUX2_X1 U23574 ( .A(_03097__PTR1), .B(_03097__PTR129), .S(P2_P1_State2_PTR2), .Z(_03098__PTR1) );
  MUX2_X1 U23575 ( .A(_03097__PTR2), .B(_03097__PTR130), .S(P2_P1_State2_PTR2), .Z(_03098__PTR2) );
  MUX2_X1 U23576 ( .A(_03097__PTR3), .B(_03097__PTR131), .S(P2_P1_State2_PTR2), .Z(_03098__PTR3) );
  MUX2_X1 U23577 ( .A(_03097__PTR4), .B(_03097__PTR132), .S(P2_P1_State2_PTR2), .Z(_03098__PTR4) );
  MUX2_X1 U23578 ( .A(_03097__PTR5), .B(_03097__PTR133), .S(P2_P1_State2_PTR2), .Z(_03098__PTR5) );
  MUX2_X1 U23579 ( .A(_03097__PTR6), .B(_03097__PTR134), .S(P2_P1_State2_PTR2), .Z(_03098__PTR6) );
  MUX2_X1 U23580 ( .A(_03097__PTR7), .B(_03097__PTR135), .S(P2_P1_State2_PTR2), .Z(_03098__PTR7) );
  MUX2_X1 U23581 ( .A(_03097__PTR8), .B(_03097__PTR136), .S(P2_P1_State2_PTR2), .Z(_03098__PTR8) );
  MUX2_X1 U23582 ( .A(_03097__PTR9), .B(_03097__PTR137), .S(P2_P1_State2_PTR2), .Z(_03098__PTR9) );
  MUX2_X1 U23583 ( .A(_03097__PTR10), .B(_03097__PTR138), .S(P2_P1_State2_PTR2), .Z(_03098__PTR10) );
  MUX2_X1 U23584 ( .A(_03097__PTR11), .B(_03097__PTR139), .S(P2_P1_State2_PTR2), .Z(_03098__PTR11) );
  MUX2_X1 U23585 ( .A(_03097__PTR12), .B(_03097__PTR140), .S(P2_P1_State2_PTR2), .Z(_03098__PTR12) );
  MUX2_X1 U23586 ( .A(_03097__PTR13), .B(_03097__PTR141), .S(P2_P1_State2_PTR2), .Z(_03098__PTR13) );
  MUX2_X1 U23587 ( .A(_03097__PTR14), .B(_03097__PTR142), .S(P2_P1_State2_PTR2), .Z(_03098__PTR14) );
  MUX2_X1 U23588 ( .A(_03097__PTR15), .B(_03097__PTR143), .S(P2_P1_State2_PTR2), .Z(_03098__PTR15) );
  MUX2_X1 U23589 ( .A(_03097__PTR16), .B(_03097__PTR144), .S(P2_P1_State2_PTR2), .Z(_03098__PTR16) );
  MUX2_X1 U23590 ( .A(_03097__PTR17), .B(_03097__PTR145), .S(P2_P1_State2_PTR2), .Z(_03098__PTR17) );
  MUX2_X1 U23591 ( .A(_03097__PTR18), .B(_03097__PTR146), .S(P2_P1_State2_PTR2), .Z(_03098__PTR18) );
  MUX2_X1 U23592 ( .A(_03097__PTR19), .B(_03097__PTR147), .S(P2_P1_State2_PTR2), .Z(_03098__PTR19) );
  MUX2_X1 U23593 ( .A(_03097__PTR20), .B(_03097__PTR148), .S(P2_P1_State2_PTR2), .Z(_03098__PTR20) );
  MUX2_X1 U23594 ( .A(_03097__PTR21), .B(_03097__PTR149), .S(P2_P1_State2_PTR2), .Z(_03098__PTR21) );
  MUX2_X1 U23595 ( .A(_03097__PTR22), .B(_03097__PTR150), .S(P2_P1_State2_PTR2), .Z(_03098__PTR22) );
  MUX2_X1 U23596 ( .A(_03097__PTR23), .B(_03097__PTR151), .S(P2_P1_State2_PTR2), .Z(_03098__PTR23) );
  MUX2_X1 U23597 ( .A(_03097__PTR24), .B(_03097__PTR152), .S(P2_P1_State2_PTR2), .Z(_03098__PTR24) );
  MUX2_X1 U23598 ( .A(_03097__PTR25), .B(_03097__PTR153), .S(P2_P1_State2_PTR2), .Z(_03098__PTR25) );
  MUX2_X1 U23599 ( .A(_03097__PTR26), .B(_03097__PTR154), .S(P2_P1_State2_PTR2), .Z(_03098__PTR26) );
  MUX2_X1 U23600 ( .A(_03097__PTR27), .B(_03097__PTR155), .S(P2_P1_State2_PTR2), .Z(_03098__PTR27) );
  MUX2_X1 U23601 ( .A(_03097__PTR28), .B(_03097__PTR156), .S(P2_P1_State2_PTR2), .Z(_03098__PTR28) );
  MUX2_X1 U23602 ( .A(_03097__PTR29), .B(_03097__PTR157), .S(P2_P1_State2_PTR2), .Z(_03098__PTR29) );
  MUX2_X1 U23603 ( .A(_03097__PTR30), .B(_03097__PTR158), .S(P2_P1_State2_PTR2), .Z(_03098__PTR30) );
  MUX2_X1 U23604 ( .A(_03097__PTR31), .B(_03097__PTR159), .S(P2_P1_State2_PTR2), .Z(_03098__PTR31) );
  MUX2_X1 U23605 ( .A(_03096__PTR0), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR0) );
  MUX2_X1 U23606 ( .A(_03096__PTR1), .B(_03096__PTR65), .S(P2_P1_State2_PTR1), .Z(_03097__PTR1) );
  MUX2_X1 U23607 ( .A(_03096__PTR2), .B(_03096__PTR66), .S(P2_P1_State2_PTR1), .Z(_03097__PTR2) );
  MUX2_X1 U23608 ( .A(_03096__PTR3), .B(_03096__PTR67), .S(P2_P1_State2_PTR1), .Z(_03097__PTR3) );
  MUX2_X1 U23609 ( .A(_03096__PTR4), .B(_03096__PTR68), .S(P2_P1_State2_PTR1), .Z(_03097__PTR4) );
  MUX2_X1 U23610 ( .A(_03096__PTR5), .B(_03096__PTR69), .S(P2_P1_State2_PTR1), .Z(_03097__PTR5) );
  MUX2_X1 U23611 ( .A(_03096__PTR6), .B(_03096__PTR70), .S(P2_P1_State2_PTR1), .Z(_03097__PTR6) );
  MUX2_X1 U23612 ( .A(_03096__PTR7), .B(_03096__PTR71), .S(P2_P1_State2_PTR1), .Z(_03097__PTR7) );
  MUX2_X1 U23613 ( .A(_03096__PTR8), .B(_03096__PTR72), .S(P2_P1_State2_PTR1), .Z(_03097__PTR8) );
  MUX2_X1 U23614 ( .A(_03096__PTR9), .B(_03096__PTR73), .S(P2_P1_State2_PTR1), .Z(_03097__PTR9) );
  MUX2_X1 U23615 ( .A(_03096__PTR10), .B(_03096__PTR74), .S(P2_P1_State2_PTR1), .Z(_03097__PTR10) );
  MUX2_X1 U23616 ( .A(_03096__PTR11), .B(_03096__PTR75), .S(P2_P1_State2_PTR1), .Z(_03097__PTR11) );
  MUX2_X1 U23617 ( .A(_03096__PTR12), .B(_03096__PTR76), .S(P2_P1_State2_PTR1), .Z(_03097__PTR12) );
  MUX2_X1 U23618 ( .A(_03096__PTR13), .B(_03096__PTR77), .S(P2_P1_State2_PTR1), .Z(_03097__PTR13) );
  MUX2_X1 U23619 ( .A(_03096__PTR14), .B(_03096__PTR78), .S(P2_P1_State2_PTR1), .Z(_03097__PTR14) );
  MUX2_X1 U23620 ( .A(_03096__PTR15), .B(_03096__PTR79), .S(P2_P1_State2_PTR1), .Z(_03097__PTR15) );
  MUX2_X1 U23621 ( .A(_03096__PTR16), .B(_03096__PTR80), .S(P2_P1_State2_PTR1), .Z(_03097__PTR16) );
  MUX2_X1 U23622 ( .A(_03096__PTR17), .B(_03096__PTR81), .S(P2_P1_State2_PTR1), .Z(_03097__PTR17) );
  MUX2_X1 U23623 ( .A(_03096__PTR18), .B(_03096__PTR82), .S(P2_P1_State2_PTR1), .Z(_03097__PTR18) );
  MUX2_X1 U23624 ( .A(_03096__PTR19), .B(_03096__PTR83), .S(P2_P1_State2_PTR1), .Z(_03097__PTR19) );
  MUX2_X1 U23625 ( .A(_03096__PTR20), .B(_03096__PTR84), .S(P2_P1_State2_PTR1), .Z(_03097__PTR20) );
  MUX2_X1 U23626 ( .A(_03096__PTR21), .B(_03096__PTR85), .S(P2_P1_State2_PTR1), .Z(_03097__PTR21) );
  MUX2_X1 U23627 ( .A(_03096__PTR22), .B(_03096__PTR86), .S(P2_P1_State2_PTR1), .Z(_03097__PTR22) );
  MUX2_X1 U23628 ( .A(_03096__PTR23), .B(_03096__PTR87), .S(P2_P1_State2_PTR1), .Z(_03097__PTR23) );
  MUX2_X1 U23629 ( .A(_03096__PTR24), .B(_03096__PTR88), .S(P2_P1_State2_PTR1), .Z(_03097__PTR24) );
  MUX2_X1 U23630 ( .A(_03096__PTR25), .B(_03096__PTR89), .S(P2_P1_State2_PTR1), .Z(_03097__PTR25) );
  MUX2_X1 U23631 ( .A(_03096__PTR26), .B(_03096__PTR90), .S(P2_P1_State2_PTR1), .Z(_03097__PTR26) );
  MUX2_X1 U23632 ( .A(_03096__PTR27), .B(_03096__PTR91), .S(P2_P1_State2_PTR1), .Z(_03097__PTR27) );
  MUX2_X1 U23633 ( .A(_03096__PTR28), .B(_03096__PTR92), .S(P2_P1_State2_PTR1), .Z(_03097__PTR28) );
  MUX2_X1 U23634 ( .A(_03096__PTR29), .B(_03096__PTR93), .S(P2_P1_State2_PTR1), .Z(_03097__PTR29) );
  MUX2_X1 U23635 ( .A(_03096__PTR30), .B(_03096__PTR94), .S(P2_P1_State2_PTR1), .Z(_03097__PTR30) );
  MUX2_X1 U23636 ( .A(_03096__PTR31), .B(_03096__PTR95), .S(P2_P1_State2_PTR1), .Z(_03097__PTR31) );
  MUX2_X1 U23637 ( .A(_03096__PTR128), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR128) );
  MUX2_X1 U23638 ( .A(_03096__PTR129), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR129) );
  MUX2_X1 U23639 ( .A(_03096__PTR130), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR130) );
  MUX2_X1 U23640 ( .A(_03096__PTR131), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR131) );
  MUX2_X1 U23641 ( .A(_03096__PTR132), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR132) );
  MUX2_X1 U23642 ( .A(_03096__PTR133), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR133) );
  MUX2_X1 U23643 ( .A(_03096__PTR134), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR134) );
  MUX2_X1 U23644 ( .A(_03096__PTR135), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR135) );
  MUX2_X1 U23645 ( .A(_03096__PTR136), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR136) );
  MUX2_X1 U23646 ( .A(_03096__PTR137), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR137) );
  MUX2_X1 U23647 ( .A(_03096__PTR138), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR138) );
  MUX2_X1 U23648 ( .A(_03096__PTR139), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR139) );
  MUX2_X1 U23649 ( .A(_03096__PTR140), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR140) );
  MUX2_X1 U23650 ( .A(_03096__PTR141), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR141) );
  MUX2_X1 U23651 ( .A(_03096__PTR142), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR142) );
  MUX2_X1 U23652 ( .A(_03096__PTR143), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR143) );
  MUX2_X1 U23653 ( .A(_03096__PTR144), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR144) );
  MUX2_X1 U23654 ( .A(_03096__PTR145), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR145) );
  MUX2_X1 U23655 ( .A(_03096__PTR146), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR146) );
  MUX2_X1 U23656 ( .A(_03096__PTR147), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR147) );
  MUX2_X1 U23657 ( .A(_03096__PTR148), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR148) );
  MUX2_X1 U23658 ( .A(_03096__PTR149), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR149) );
  MUX2_X1 U23659 ( .A(_03096__PTR150), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR150) );
  MUX2_X1 U23660 ( .A(_03096__PTR151), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR151) );
  MUX2_X1 U23661 ( .A(_03096__PTR152), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR152) );
  MUX2_X1 U23662 ( .A(_03096__PTR153), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR153) );
  MUX2_X1 U23663 ( .A(_03096__PTR154), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR154) );
  MUX2_X1 U23664 ( .A(_03096__PTR155), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR155) );
  MUX2_X1 U23665 ( .A(_03096__PTR156), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR156) );
  MUX2_X1 U23666 ( .A(_03096__PTR157), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR157) );
  MUX2_X1 U23667 ( .A(_03096__PTR158), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR158) );
  MUX2_X1 U23668 ( .A(_03096__PTR159), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03097__PTR159) );
  MUX2_X1 U23669 ( .A(P2_rEIP_PTR0), .B(P2_P1_PhyAddrPointer_PTR0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR0) );
  MUX2_X1 U23670 ( .A(P2_rEIP_PTR1), .B(P2_P1_PhyAddrPointer_PTR1), .S(P2_P1_State2_PTR0), .Z(_03096__PTR1) );
  MUX2_X1 U23671 ( .A(P2_rEIP_PTR2), .B(P2_P1_PhyAddrPointer_PTR2), .S(P2_P1_State2_PTR0), .Z(_03096__PTR2) );
  MUX2_X1 U23672 ( .A(P2_rEIP_PTR3), .B(P2_P1_PhyAddrPointer_PTR3), .S(P2_P1_State2_PTR0), .Z(_03096__PTR3) );
  MUX2_X1 U23673 ( .A(P2_rEIP_PTR4), .B(P2_P1_PhyAddrPointer_PTR4), .S(P2_P1_State2_PTR0), .Z(_03096__PTR4) );
  MUX2_X1 U23674 ( .A(P2_rEIP_PTR5), .B(P2_P1_PhyAddrPointer_PTR5), .S(P2_P1_State2_PTR0), .Z(_03096__PTR5) );
  MUX2_X1 U23675 ( .A(P2_rEIP_PTR6), .B(P2_P1_PhyAddrPointer_PTR6), .S(P2_P1_State2_PTR0), .Z(_03096__PTR6) );
  MUX2_X1 U23676 ( .A(P2_rEIP_PTR7), .B(P2_P1_PhyAddrPointer_PTR7), .S(P2_P1_State2_PTR0), .Z(_03096__PTR7) );
  MUX2_X1 U23677 ( .A(P2_rEIP_PTR8), .B(P2_P1_PhyAddrPointer_PTR8), .S(P2_P1_State2_PTR0), .Z(_03096__PTR8) );
  MUX2_X1 U23678 ( .A(P2_rEIP_PTR9), .B(P2_P1_PhyAddrPointer_PTR9), .S(P2_P1_State2_PTR0), .Z(_03096__PTR9) );
  MUX2_X1 U23679 ( .A(P2_rEIP_PTR10), .B(P2_P1_PhyAddrPointer_PTR10), .S(P2_P1_State2_PTR0), .Z(_03096__PTR10) );
  MUX2_X1 U23680 ( .A(P2_rEIP_PTR11), .B(P2_P1_PhyAddrPointer_PTR11), .S(P2_P1_State2_PTR0), .Z(_03096__PTR11) );
  MUX2_X1 U23681 ( .A(P2_rEIP_PTR12), .B(P2_P1_PhyAddrPointer_PTR12), .S(P2_P1_State2_PTR0), .Z(_03096__PTR12) );
  MUX2_X1 U23682 ( .A(P2_rEIP_PTR13), .B(P2_P1_PhyAddrPointer_PTR13), .S(P2_P1_State2_PTR0), .Z(_03096__PTR13) );
  MUX2_X1 U23683 ( .A(P2_rEIP_PTR14), .B(P2_P1_PhyAddrPointer_PTR14), .S(P2_P1_State2_PTR0), .Z(_03096__PTR14) );
  MUX2_X1 U23684 ( .A(P2_rEIP_PTR15), .B(P2_P1_PhyAddrPointer_PTR15), .S(P2_P1_State2_PTR0), .Z(_03096__PTR15) );
  MUX2_X1 U23685 ( .A(P2_rEIP_PTR16), .B(P2_P1_PhyAddrPointer_PTR16), .S(P2_P1_State2_PTR0), .Z(_03096__PTR16) );
  MUX2_X1 U23686 ( .A(P2_rEIP_PTR17), .B(P2_P1_PhyAddrPointer_PTR17), .S(P2_P1_State2_PTR0), .Z(_03096__PTR17) );
  MUX2_X1 U23687 ( .A(P2_rEIP_PTR18), .B(P2_P1_PhyAddrPointer_PTR18), .S(P2_P1_State2_PTR0), .Z(_03096__PTR18) );
  MUX2_X1 U23688 ( .A(P2_rEIP_PTR19), .B(P2_P1_PhyAddrPointer_PTR19), .S(P2_P1_State2_PTR0), .Z(_03096__PTR19) );
  MUX2_X1 U23689 ( .A(P2_rEIP_PTR20), .B(P2_P1_PhyAddrPointer_PTR20), .S(P2_P1_State2_PTR0), .Z(_03096__PTR20) );
  MUX2_X1 U23690 ( .A(P2_rEIP_PTR21), .B(P2_P1_PhyAddrPointer_PTR21), .S(P2_P1_State2_PTR0), .Z(_03096__PTR21) );
  MUX2_X1 U23691 ( .A(P2_rEIP_PTR22), .B(P2_P1_PhyAddrPointer_PTR22), .S(P2_P1_State2_PTR0), .Z(_03096__PTR22) );
  MUX2_X1 U23692 ( .A(P2_rEIP_PTR23), .B(P2_P1_PhyAddrPointer_PTR23), .S(P2_P1_State2_PTR0), .Z(_03096__PTR23) );
  MUX2_X1 U23693 ( .A(P2_rEIP_PTR24), .B(P2_P1_PhyAddrPointer_PTR24), .S(P2_P1_State2_PTR0), .Z(_03096__PTR24) );
  MUX2_X1 U23694 ( .A(P2_rEIP_PTR25), .B(P2_P1_PhyAddrPointer_PTR25), .S(P2_P1_State2_PTR0), .Z(_03096__PTR25) );
  MUX2_X1 U23695 ( .A(P2_rEIP_PTR26), .B(P2_P1_PhyAddrPointer_PTR26), .S(P2_P1_State2_PTR0), .Z(_03096__PTR26) );
  MUX2_X1 U23696 ( .A(P2_rEIP_PTR27), .B(P2_P1_PhyAddrPointer_PTR27), .S(P2_P1_State2_PTR0), .Z(_03096__PTR27) );
  MUX2_X1 U23697 ( .A(P2_rEIP_PTR28), .B(P2_P1_PhyAddrPointer_PTR28), .S(P2_P1_State2_PTR0), .Z(_03096__PTR28) );
  MUX2_X1 U23698 ( .A(P2_rEIP_PTR29), .B(P2_P1_PhyAddrPointer_PTR29), .S(P2_P1_State2_PTR0), .Z(_03096__PTR29) );
  MUX2_X1 U23699 ( .A(P2_rEIP_PTR30), .B(P2_P1_PhyAddrPointer_PTR30), .S(P2_P1_State2_PTR0), .Z(_03096__PTR30) );
  MUX2_X1 U23700 ( .A(P2_rEIP_PTR31), .B(P2_P1_PhyAddrPointer_PTR31), .S(P2_P1_State2_PTR0), .Z(_03096__PTR31) );
  MUX2_X1 U23701 ( .A(_02184__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR65) );
  MUX2_X1 U23702 ( .A(_02184__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR66) );
  MUX2_X1 U23703 ( .A(_02184__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR67) );
  MUX2_X1 U23704 ( .A(_02184__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR68) );
  MUX2_X1 U23705 ( .A(_02184__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR69) );
  MUX2_X1 U23706 ( .A(_02184__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR70) );
  MUX2_X1 U23707 ( .A(_02184__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR71) );
  MUX2_X1 U23708 ( .A(_02184__PTR72), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR72) );
  MUX2_X1 U23709 ( .A(_02184__PTR73), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR73) );
  MUX2_X1 U23710 ( .A(_02184__PTR74), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR74) );
  MUX2_X1 U23711 ( .A(_02184__PTR75), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR75) );
  MUX2_X1 U23712 ( .A(_02184__PTR76), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR76) );
  MUX2_X1 U23713 ( .A(_02184__PTR77), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR77) );
  MUX2_X1 U23714 ( .A(_02184__PTR78), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR78) );
  MUX2_X1 U23715 ( .A(_02184__PTR79), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR79) );
  MUX2_X1 U23716 ( .A(_02184__PTR80), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR80) );
  MUX2_X1 U23717 ( .A(_02184__PTR81), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR81) );
  MUX2_X1 U23718 ( .A(_02184__PTR82), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR82) );
  MUX2_X1 U23719 ( .A(_02184__PTR83), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR83) );
  MUX2_X1 U23720 ( .A(_02184__PTR84), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR84) );
  MUX2_X1 U23721 ( .A(_02184__PTR85), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR85) );
  MUX2_X1 U23722 ( .A(_02184__PTR86), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR86) );
  MUX2_X1 U23723 ( .A(_02184__PTR87), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR87) );
  MUX2_X1 U23724 ( .A(_02184__PTR88), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR88) );
  MUX2_X1 U23725 ( .A(_02184__PTR89), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR89) );
  MUX2_X1 U23726 ( .A(_02184__PTR90), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR90) );
  MUX2_X1 U23727 ( .A(_02184__PTR91), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR91) );
  MUX2_X1 U23728 ( .A(_02184__PTR92), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR92) );
  MUX2_X1 U23729 ( .A(_02184__PTR93), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR93) );
  MUX2_X1 U23730 ( .A(_02184__PTR94), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR94) );
  MUX2_X1 U23731 ( .A(_02184__PTR95), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03096__PTR95) );
  MUX2_X1 U23732 ( .A(1'b0), .B(_02184__PTR160), .S(P2_P1_State2_PTR0), .Z(_03096__PTR128) );
  MUX2_X1 U23733 ( .A(_02184__PTR129), .B(_02184__PTR161), .S(P2_P1_State2_PTR0), .Z(_03096__PTR129) );
  MUX2_X1 U23734 ( .A(_02184__PTR130), .B(_02184__PTR162), .S(P2_P1_State2_PTR0), .Z(_03096__PTR130) );
  MUX2_X1 U23735 ( .A(_02184__PTR131), .B(_02184__PTR163), .S(P2_P1_State2_PTR0), .Z(_03096__PTR131) );
  MUX2_X1 U23736 ( .A(_02184__PTR132), .B(_02184__PTR164), .S(P2_P1_State2_PTR0), .Z(_03096__PTR132) );
  MUX2_X1 U23737 ( .A(_02184__PTR133), .B(_02184__PTR165), .S(P2_P1_State2_PTR0), .Z(_03096__PTR133) );
  MUX2_X1 U23738 ( .A(_02184__PTR134), .B(_02184__PTR166), .S(P2_P1_State2_PTR0), .Z(_03096__PTR134) );
  MUX2_X1 U23739 ( .A(_02184__PTR135), .B(_02184__PTR167), .S(P2_P1_State2_PTR0), .Z(_03096__PTR135) );
  MUX2_X1 U23740 ( .A(_02184__PTR136), .B(_02184__PTR168), .S(P2_P1_State2_PTR0), .Z(_03096__PTR136) );
  MUX2_X1 U23741 ( .A(_02184__PTR137), .B(_02184__PTR169), .S(P2_P1_State2_PTR0), .Z(_03096__PTR137) );
  MUX2_X1 U23742 ( .A(_02184__PTR138), .B(_02184__PTR170), .S(P2_P1_State2_PTR0), .Z(_03096__PTR138) );
  MUX2_X1 U23743 ( .A(_02184__PTR139), .B(_02184__PTR171), .S(P2_P1_State2_PTR0), .Z(_03096__PTR139) );
  MUX2_X1 U23744 ( .A(_02184__PTR140), .B(_02184__PTR172), .S(P2_P1_State2_PTR0), .Z(_03096__PTR140) );
  MUX2_X1 U23745 ( .A(_02184__PTR141), .B(_02184__PTR173), .S(P2_P1_State2_PTR0), .Z(_03096__PTR141) );
  MUX2_X1 U23746 ( .A(_02184__PTR142), .B(_02184__PTR174), .S(P2_P1_State2_PTR0), .Z(_03096__PTR142) );
  MUX2_X1 U23747 ( .A(_02184__PTR143), .B(_02184__PTR175), .S(P2_P1_State2_PTR0), .Z(_03096__PTR143) );
  MUX2_X1 U23748 ( .A(_02184__PTR144), .B(_02184__PTR176), .S(P2_P1_State2_PTR0), .Z(_03096__PTR144) );
  MUX2_X1 U23749 ( .A(_02184__PTR145), .B(_02184__PTR177), .S(P2_P1_State2_PTR0), .Z(_03096__PTR145) );
  MUX2_X1 U23750 ( .A(_02184__PTR146), .B(_02184__PTR178), .S(P2_P1_State2_PTR0), .Z(_03096__PTR146) );
  MUX2_X1 U23751 ( .A(_02184__PTR147), .B(_02184__PTR179), .S(P2_P1_State2_PTR0), .Z(_03096__PTR147) );
  MUX2_X1 U23752 ( .A(_02184__PTR148), .B(_02184__PTR180), .S(P2_P1_State2_PTR0), .Z(_03096__PTR148) );
  MUX2_X1 U23753 ( .A(_02184__PTR149), .B(_02184__PTR181), .S(P2_P1_State2_PTR0), .Z(_03096__PTR149) );
  MUX2_X1 U23754 ( .A(_02184__PTR150), .B(_02184__PTR182), .S(P2_P1_State2_PTR0), .Z(_03096__PTR150) );
  MUX2_X1 U23755 ( .A(_02184__PTR151), .B(_02184__PTR183), .S(P2_P1_State2_PTR0), .Z(_03096__PTR151) );
  MUX2_X1 U23756 ( .A(_02184__PTR152), .B(_02184__PTR184), .S(P2_P1_State2_PTR0), .Z(_03096__PTR152) );
  MUX2_X1 U23757 ( .A(_02184__PTR153), .B(_02184__PTR185), .S(P2_P1_State2_PTR0), .Z(_03096__PTR153) );
  MUX2_X1 U23758 ( .A(_02184__PTR154), .B(_02184__PTR186), .S(P2_P1_State2_PTR0), .Z(_03096__PTR154) );
  MUX2_X1 U23759 ( .A(_02184__PTR155), .B(_02184__PTR187), .S(P2_P1_State2_PTR0), .Z(_03096__PTR155) );
  MUX2_X1 U23760 ( .A(_02184__PTR156), .B(_02184__PTR188), .S(P2_P1_State2_PTR0), .Z(_03096__PTR156) );
  MUX2_X1 U23761 ( .A(_02184__PTR157), .B(_02184__PTR189), .S(P2_P1_State2_PTR0), .Z(_03096__PTR157) );
  MUX2_X1 U23762 ( .A(_02184__PTR158), .B(_02184__PTR190), .S(P2_P1_State2_PTR0), .Z(_03096__PTR158) );
  MUX2_X1 U23763 ( .A(_02184__PTR159), .B(_02184__PTR191), .S(P2_P1_State2_PTR0), .Z(_03096__PTR159) );
  MUX2_X1 U23764 ( .A(_03100__PTR0), .B(_03100__PTR128), .S(P2_P1_State2_PTR2), .Z(_03101__PTR0) );
  MUX2_X1 U23765 ( .A(_03100__PTR1), .B(_03100__PTR129), .S(P2_P1_State2_PTR2), .Z(_03101__PTR1) );
  MUX2_X1 U23766 ( .A(_03100__PTR2), .B(_03100__PTR130), .S(P2_P1_State2_PTR2), .Z(_03101__PTR2) );
  MUX2_X1 U23767 ( .A(_03100__PTR3), .B(_03100__PTR131), .S(P2_P1_State2_PTR2), .Z(_03101__PTR3) );
  MUX2_X1 U23768 ( .A(_03100__PTR4), .B(_03100__PTR132), .S(P2_P1_State2_PTR2), .Z(_03101__PTR4) );
  MUX2_X1 U23769 ( .A(_03100__PTR5), .B(_03100__PTR133), .S(P2_P1_State2_PTR2), .Z(_03101__PTR5) );
  MUX2_X1 U23770 ( .A(_03100__PTR6), .B(_03100__PTR134), .S(P2_P1_State2_PTR2), .Z(_03101__PTR6) );
  MUX2_X1 U23771 ( .A(_03100__PTR7), .B(_03100__PTR135), .S(P2_P1_State2_PTR2), .Z(_03101__PTR7) );
  MUX2_X1 U23772 ( .A(_03100__PTR8), .B(_03100__PTR136), .S(P2_P1_State2_PTR2), .Z(_03101__PTR8) );
  MUX2_X1 U23773 ( .A(_03100__PTR9), .B(_03100__PTR137), .S(P2_P1_State2_PTR2), .Z(_03101__PTR9) );
  MUX2_X1 U23774 ( .A(_03100__PTR10), .B(_03100__PTR138), .S(P2_P1_State2_PTR2), .Z(_03101__PTR10) );
  MUX2_X1 U23775 ( .A(_03100__PTR11), .B(_03100__PTR139), .S(P2_P1_State2_PTR2), .Z(_03101__PTR11) );
  MUX2_X1 U23776 ( .A(_03100__PTR12), .B(_03100__PTR140), .S(P2_P1_State2_PTR2), .Z(_03101__PTR12) );
  MUX2_X1 U23777 ( .A(_03100__PTR13), .B(_03100__PTR141), .S(P2_P1_State2_PTR2), .Z(_03101__PTR13) );
  MUX2_X1 U23778 ( .A(_03100__PTR14), .B(_03100__PTR142), .S(P2_P1_State2_PTR2), .Z(_03101__PTR14) );
  MUX2_X1 U23779 ( .A(_03100__PTR15), .B(_03100__PTR143), .S(P2_P1_State2_PTR2), .Z(_03101__PTR15) );
  MUX2_X1 U23780 ( .A(_03100__PTR16), .B(_03100__PTR144), .S(P2_P1_State2_PTR2), .Z(_03101__PTR16) );
  MUX2_X1 U23781 ( .A(_03100__PTR17), .B(_03100__PTR145), .S(P2_P1_State2_PTR2), .Z(_03101__PTR17) );
  MUX2_X1 U23782 ( .A(_03100__PTR18), .B(_03100__PTR146), .S(P2_P1_State2_PTR2), .Z(_03101__PTR18) );
  MUX2_X1 U23783 ( .A(_03100__PTR19), .B(_03100__PTR147), .S(P2_P1_State2_PTR2), .Z(_03101__PTR19) );
  MUX2_X1 U23784 ( .A(_03100__PTR20), .B(_03100__PTR148), .S(P2_P1_State2_PTR2), .Z(_03101__PTR20) );
  MUX2_X1 U23785 ( .A(_03100__PTR21), .B(_03100__PTR149), .S(P2_P1_State2_PTR2), .Z(_03101__PTR21) );
  MUX2_X1 U23786 ( .A(_03100__PTR22), .B(_03100__PTR150), .S(P2_P1_State2_PTR2), .Z(_03101__PTR22) );
  MUX2_X1 U23787 ( .A(_03100__PTR23), .B(_03100__PTR151), .S(P2_P1_State2_PTR2), .Z(_03101__PTR23) );
  MUX2_X1 U23788 ( .A(_03100__PTR24), .B(_03100__PTR152), .S(P2_P1_State2_PTR2), .Z(_03101__PTR24) );
  MUX2_X1 U23789 ( .A(_03100__PTR25), .B(_03100__PTR153), .S(P2_P1_State2_PTR2), .Z(_03101__PTR25) );
  MUX2_X1 U23790 ( .A(_03100__PTR26), .B(_03100__PTR154), .S(P2_P1_State2_PTR2), .Z(_03101__PTR26) );
  MUX2_X1 U23791 ( .A(_03100__PTR27), .B(_03100__PTR155), .S(P2_P1_State2_PTR2), .Z(_03101__PTR27) );
  MUX2_X1 U23792 ( .A(_03100__PTR28), .B(_03100__PTR156), .S(P2_P1_State2_PTR2), .Z(_03101__PTR28) );
  MUX2_X1 U23793 ( .A(_03100__PTR29), .B(_03100__PTR157), .S(P2_P1_State2_PTR2), .Z(_03101__PTR29) );
  MUX2_X1 U23794 ( .A(_03100__PTR30), .B(_03100__PTR158), .S(P2_P1_State2_PTR2), .Z(_03101__PTR30) );
  MUX2_X1 U23795 ( .A(_03100__PTR31), .B(_03100__PTR159), .S(P2_P1_State2_PTR2), .Z(_03101__PTR31) );
  MUX2_X1 U23796 ( .A(_03099__PTR0), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR0) );
  MUX2_X1 U23797 ( .A(_03099__PTR1), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR1) );
  MUX2_X1 U23798 ( .A(_03099__PTR2), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR2) );
  MUX2_X1 U23799 ( .A(_03099__PTR3), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR3) );
  MUX2_X1 U23800 ( .A(_03099__PTR4), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR4) );
  MUX2_X1 U23801 ( .A(_03099__PTR5), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR5) );
  MUX2_X1 U23802 ( .A(_03099__PTR6), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR6) );
  MUX2_X1 U23803 ( .A(_03099__PTR7), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR7) );
  MUX2_X1 U23804 ( .A(_03099__PTR8), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR8) );
  MUX2_X1 U23805 ( .A(_03099__PTR9), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR9) );
  MUX2_X1 U23806 ( .A(_03099__PTR10), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR10) );
  MUX2_X1 U23807 ( .A(_03099__PTR11), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR11) );
  MUX2_X1 U23808 ( .A(_03099__PTR12), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR12) );
  MUX2_X1 U23809 ( .A(_03099__PTR13), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR13) );
  MUX2_X1 U23810 ( .A(_03099__PTR14), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR14) );
  MUX2_X1 U23811 ( .A(_03099__PTR15), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR15) );
  MUX2_X1 U23812 ( .A(_03099__PTR16), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR16) );
  MUX2_X1 U23813 ( .A(_03099__PTR17), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR17) );
  MUX2_X1 U23814 ( .A(_03099__PTR18), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR18) );
  MUX2_X1 U23815 ( .A(_03099__PTR19), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR19) );
  MUX2_X1 U23816 ( .A(_03099__PTR20), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR20) );
  MUX2_X1 U23817 ( .A(_03099__PTR21), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR21) );
  MUX2_X1 U23818 ( .A(_03099__PTR22), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR22) );
  MUX2_X1 U23819 ( .A(_03099__PTR23), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR23) );
  MUX2_X1 U23820 ( .A(_03099__PTR24), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR24) );
  MUX2_X1 U23821 ( .A(_03099__PTR25), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR25) );
  MUX2_X1 U23822 ( .A(_03099__PTR26), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR26) );
  MUX2_X1 U23823 ( .A(_03099__PTR27), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR27) );
  MUX2_X1 U23824 ( .A(_03099__PTR28), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR28) );
  MUX2_X1 U23825 ( .A(_03099__PTR29), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR29) );
  MUX2_X1 U23826 ( .A(_03099__PTR30), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR30) );
  MUX2_X1 U23827 ( .A(_03099__PTR31), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR31) );
  MUX2_X1 U23828 ( .A(_03099__PTR128), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR128) );
  MUX2_X1 U23829 ( .A(_03099__PTR129), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR129) );
  MUX2_X1 U23830 ( .A(_03099__PTR130), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR130) );
  MUX2_X1 U23831 ( .A(_03099__PTR131), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR131) );
  MUX2_X1 U23832 ( .A(_03099__PTR132), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR132) );
  MUX2_X1 U23833 ( .A(_03099__PTR133), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR133) );
  MUX2_X1 U23834 ( .A(_03099__PTR134), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR134) );
  MUX2_X1 U23835 ( .A(_03099__PTR135), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR135) );
  MUX2_X1 U23836 ( .A(_03099__PTR136), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR136) );
  MUX2_X1 U23837 ( .A(_03099__PTR137), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR137) );
  MUX2_X1 U23838 ( .A(_03099__PTR138), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR138) );
  MUX2_X1 U23839 ( .A(_03099__PTR139), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR139) );
  MUX2_X1 U23840 ( .A(_03099__PTR140), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR140) );
  MUX2_X1 U23841 ( .A(_03099__PTR141), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR141) );
  MUX2_X1 U23842 ( .A(_03099__PTR142), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR142) );
  MUX2_X1 U23843 ( .A(_03099__PTR143), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR143) );
  MUX2_X1 U23844 ( .A(_03099__PTR144), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR144) );
  MUX2_X1 U23845 ( .A(_03099__PTR145), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR145) );
  MUX2_X1 U23846 ( .A(_03099__PTR146), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR146) );
  MUX2_X1 U23847 ( .A(_03099__PTR147), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR147) );
  MUX2_X1 U23848 ( .A(_03099__PTR148), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR148) );
  MUX2_X1 U23849 ( .A(_03099__PTR149), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR149) );
  MUX2_X1 U23850 ( .A(_03099__PTR150), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR150) );
  MUX2_X1 U23851 ( .A(_03099__PTR151), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR151) );
  MUX2_X1 U23852 ( .A(_03099__PTR152), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR152) );
  MUX2_X1 U23853 ( .A(_03099__PTR153), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR153) );
  MUX2_X1 U23854 ( .A(_03099__PTR154), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR154) );
  MUX2_X1 U23855 ( .A(_03099__PTR155), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR155) );
  MUX2_X1 U23856 ( .A(_03099__PTR156), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR156) );
  MUX2_X1 U23857 ( .A(_03099__PTR157), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR157) );
  MUX2_X1 U23858 ( .A(_03099__PTR158), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR158) );
  MUX2_X1 U23859 ( .A(_03099__PTR159), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03100__PTR159) );
  MUX2_X1 U23860 ( .A(P2_rEIP_PTR0), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR0) );
  MUX2_X1 U23861 ( .A(P2_rEIP_PTR1), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR1) );
  MUX2_X1 U23862 ( .A(P2_rEIP_PTR2), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR2) );
  MUX2_X1 U23863 ( .A(P2_rEIP_PTR3), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR3) );
  MUX2_X1 U23864 ( .A(P2_rEIP_PTR4), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR4) );
  MUX2_X1 U23865 ( .A(P2_rEIP_PTR5), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR5) );
  MUX2_X1 U23866 ( .A(P2_rEIP_PTR6), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR6) );
  MUX2_X1 U23867 ( .A(P2_rEIP_PTR7), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR7) );
  MUX2_X1 U23868 ( .A(P2_rEIP_PTR8), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR8) );
  MUX2_X1 U23869 ( .A(P2_rEIP_PTR9), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR9) );
  MUX2_X1 U23870 ( .A(P2_rEIP_PTR10), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR10) );
  MUX2_X1 U23871 ( .A(P2_rEIP_PTR11), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR11) );
  MUX2_X1 U23872 ( .A(P2_rEIP_PTR12), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR12) );
  MUX2_X1 U23873 ( .A(P2_rEIP_PTR13), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR13) );
  MUX2_X1 U23874 ( .A(P2_rEIP_PTR14), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR14) );
  MUX2_X1 U23875 ( .A(P2_rEIP_PTR15), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR15) );
  MUX2_X1 U23876 ( .A(P2_rEIP_PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR16) );
  MUX2_X1 U23877 ( .A(P2_rEIP_PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR17) );
  MUX2_X1 U23878 ( .A(P2_rEIP_PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR18) );
  MUX2_X1 U23879 ( .A(P2_rEIP_PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR19) );
  MUX2_X1 U23880 ( .A(P2_rEIP_PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR20) );
  MUX2_X1 U23881 ( .A(P2_rEIP_PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR21) );
  MUX2_X1 U23882 ( .A(P2_rEIP_PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR22) );
  MUX2_X1 U23883 ( .A(P2_rEIP_PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR23) );
  MUX2_X1 U23884 ( .A(P2_rEIP_PTR24), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR24) );
  MUX2_X1 U23885 ( .A(P2_rEIP_PTR25), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR25) );
  MUX2_X1 U23886 ( .A(P2_rEIP_PTR26), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR26) );
  MUX2_X1 U23887 ( .A(P2_rEIP_PTR27), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR27) );
  MUX2_X1 U23888 ( .A(P2_rEIP_PTR28), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR28) );
  MUX2_X1 U23889 ( .A(P2_rEIP_PTR29), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR29) );
  MUX2_X1 U23890 ( .A(P2_rEIP_PTR30), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR30) );
  MUX2_X1 U23891 ( .A(P2_rEIP_PTR31), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03099__PTR31) );
  MUX2_X1 U23892 ( .A(1'b0), .B(_02185__PTR160), .S(P2_P1_State2_PTR0), .Z(_03099__PTR128) );
  MUX2_X1 U23893 ( .A(1'b0), .B(_02185__PTR161), .S(P2_P1_State2_PTR0), .Z(_03099__PTR129) );
  MUX2_X1 U23894 ( .A(1'b0), .B(_02185__PTR162), .S(P2_P1_State2_PTR0), .Z(_03099__PTR130) );
  MUX2_X1 U23895 ( .A(1'b0), .B(_02185__PTR163), .S(P2_P1_State2_PTR0), .Z(_03099__PTR131) );
  MUX2_X1 U23896 ( .A(1'b0), .B(_02185__PTR164), .S(P2_P1_State2_PTR0), .Z(_03099__PTR132) );
  MUX2_X1 U23897 ( .A(1'b0), .B(_02185__PTR165), .S(P2_P1_State2_PTR0), .Z(_03099__PTR133) );
  MUX2_X1 U23898 ( .A(1'b0), .B(_02185__PTR166), .S(P2_P1_State2_PTR0), .Z(_03099__PTR134) );
  MUX2_X1 U23899 ( .A(1'b0), .B(_02185__PTR167), .S(P2_P1_State2_PTR0), .Z(_03099__PTR135) );
  MUX2_X1 U23900 ( .A(1'b0), .B(_02185__PTR168), .S(P2_P1_State2_PTR0), .Z(_03099__PTR136) );
  MUX2_X1 U23901 ( .A(1'b0), .B(_02185__PTR169), .S(P2_P1_State2_PTR0), .Z(_03099__PTR137) );
  MUX2_X1 U23902 ( .A(1'b0), .B(_02185__PTR170), .S(P2_P1_State2_PTR0), .Z(_03099__PTR138) );
  MUX2_X1 U23903 ( .A(1'b0), .B(_02185__PTR171), .S(P2_P1_State2_PTR0), .Z(_03099__PTR139) );
  MUX2_X1 U23904 ( .A(1'b0), .B(_02185__PTR172), .S(P2_P1_State2_PTR0), .Z(_03099__PTR140) );
  MUX2_X1 U23905 ( .A(1'b0), .B(_02185__PTR173), .S(P2_P1_State2_PTR0), .Z(_03099__PTR141) );
  MUX2_X1 U23906 ( .A(1'b0), .B(_02185__PTR174), .S(P2_P1_State2_PTR0), .Z(_03099__PTR142) );
  MUX2_X1 U23907 ( .A(1'b0), .B(_02185__PTR175), .S(P2_P1_State2_PTR0), .Z(_03099__PTR143) );
  MUX2_X1 U23908 ( .A(1'b0), .B(_02185__PTR176), .S(P2_P1_State2_PTR0), .Z(_03099__PTR144) );
  MUX2_X1 U23909 ( .A(1'b0), .B(_02185__PTR177), .S(P2_P1_State2_PTR0), .Z(_03099__PTR145) );
  MUX2_X1 U23910 ( .A(1'b0), .B(_02185__PTR178), .S(P2_P1_State2_PTR0), .Z(_03099__PTR146) );
  MUX2_X1 U23911 ( .A(1'b0), .B(_02185__PTR179), .S(P2_P1_State2_PTR0), .Z(_03099__PTR147) );
  MUX2_X1 U23912 ( .A(1'b0), .B(_02185__PTR180), .S(P2_P1_State2_PTR0), .Z(_03099__PTR148) );
  MUX2_X1 U23913 ( .A(1'b0), .B(_02185__PTR181), .S(P2_P1_State2_PTR0), .Z(_03099__PTR149) );
  MUX2_X1 U23914 ( .A(1'b0), .B(_02185__PTR182), .S(P2_P1_State2_PTR0), .Z(_03099__PTR150) );
  MUX2_X1 U23915 ( .A(1'b0), .B(_02185__PTR183), .S(P2_P1_State2_PTR0), .Z(_03099__PTR151) );
  MUX2_X1 U23916 ( .A(1'b0), .B(_02185__PTR184), .S(P2_P1_State2_PTR0), .Z(_03099__PTR152) );
  MUX2_X1 U23917 ( .A(1'b0), .B(_02185__PTR185), .S(P2_P1_State2_PTR0), .Z(_03099__PTR153) );
  MUX2_X1 U23918 ( .A(1'b0), .B(_02185__PTR186), .S(P2_P1_State2_PTR0), .Z(_03099__PTR154) );
  MUX2_X1 U23919 ( .A(1'b0), .B(_02185__PTR187), .S(P2_P1_State2_PTR0), .Z(_03099__PTR155) );
  MUX2_X1 U23920 ( .A(1'b0), .B(_02185__PTR188), .S(P2_P1_State2_PTR0), .Z(_03099__PTR156) );
  MUX2_X1 U23921 ( .A(1'b0), .B(_02185__PTR189), .S(P2_P1_State2_PTR0), .Z(_03099__PTR157) );
  MUX2_X1 U23922 ( .A(1'b0), .B(_02185__PTR190), .S(P2_P1_State2_PTR0), .Z(_03099__PTR158) );
  MUX2_X1 U23923 ( .A(1'b0), .B(_02185__PTR191), .S(P2_P1_State2_PTR0), .Z(_03099__PTR159) );
  MUX2_X1 U23924 ( .A(_03104__PTR0), .B(_03102__PTR32), .S(P2_P1_State2_PTR3), .Z(_02187__PTR0) );
  MUX2_X1 U23925 ( .A(_03104__PTR1), .B(1'b0), .S(P2_P1_State2_PTR3), .Z(_02187__PTR1) );
  MUX2_X1 U23926 ( .A(_03104__PTR2), .B(1'b0), .S(P2_P1_State2_PTR3), .Z(_02187__PTR2) );
  MUX2_X1 U23927 ( .A(_03104__PTR3), .B(_00300_), .S(P2_P1_State2_PTR3), .Z(_02187__PTR3) );
  MUX2_X1 U23928 ( .A(_03102__PTR0), .B(_03102__PTR16), .S(P2_P1_State2_PTR2), .Z(_03104__PTR0) );
  MUX2_X1 U23929 ( .A(_03102__PTR1), .B(_03102__PTR17), .S(P2_P1_State2_PTR2), .Z(_03104__PTR1) );
  MUX2_X1 U23930 ( .A(_03102__PTR2), .B(_03102__PTR18), .S(P2_P1_State2_PTR2), .Z(_03104__PTR2) );
  MUX2_X1 U23931 ( .A(1'b0), .B(_03102__PTR19), .S(P2_P1_State2_PTR2), .Z(_03104__PTR3) );
  MUX2_X1 U23932 ( .A(_03105__PTR1), .B(_03103__PTR1), .S(P2_P1_State2_PTR1), .Z(_03102__PTR1) );
  MUX2_X1 U23933 ( .A(1'b0), .B(_03103__PTR2), .S(P2_P1_State2_PTR1), .Z(_03102__PTR2) );
  MUX2_X1 U23934 ( .A(_03103__PTR8), .B(_03103__PTR16), .S(P2_P1_State2_PTR1), .Z(_03102__PTR16) );
  MUX2_X1 U23935 ( .A(_03103__PTR9), .B(_03103__PTR17), .S(P2_P1_State2_PTR1), .Z(_03102__PTR17) );
  MUX2_X1 U23936 ( .A(_03103__PTR10), .B(_03103__PTR18), .S(P2_P1_State2_PTR1), .Z(_03102__PTR18) );
  MUX2_X1 U23937 ( .A(_03103__PTR11), .B(_03103__PTR19), .S(P2_P1_State2_PTR1), .Z(_03102__PTR19) );
  MUX2_X1 U23938 ( .A(1'b0), .B(_02186__PTR14), .S(P2_P1_State2_PTR0), .Z(_03105__PTR1) );
  MUX2_X1 U23939 ( .A(1'b1), .B(P2_READY_n), .S(P2_P1_State2_PTR0), .Z(_03102__PTR0) );
  MUX2_X1 U23940 ( .A(_02186__PTR9), .B(P2_READY_n), .S(P2_P1_State2_PTR0), .Z(_03103__PTR1) );
  MUX2_X1 U23941 ( .A(P2_StateBS16), .B(_02186__PTR14), .S(P2_P1_State2_PTR0), .Z(_03103__PTR2) );
  MUX2_X1 U23942 ( .A(1'b1), .B(_02186__PTR20), .S(P2_P1_State2_PTR0), .Z(_03103__PTR8) );
  MUX2_X1 U23943 ( .A(1'b0), .B(_02186__PTR21), .S(P2_P1_State2_PTR0), .Z(_03103__PTR9) );
  MUX2_X1 U23944 ( .A(1'b1), .B(_02186__PTR22), .S(P2_P1_State2_PTR0), .Z(_03103__PTR10) );
  MUX2_X1 U23945 ( .A(1'b0), .B(_02186__PTR23), .S(P2_P1_State2_PTR0), .Z(_03103__PTR11) );
  MUX2_X1 U23946 ( .A(_02186__PTR26), .B(_02186__PTR28), .S(P2_P1_State2_PTR0), .Z(_03103__PTR16) );
  MUX2_X1 U23947 ( .A(_02142__PTR6), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03103__PTR17) );
  MUX2_X1 U23948 ( .A(_02186__PTR26), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03103__PTR18) );
  MUX2_X1 U23949 ( .A(_02142__PTR6), .B(1'b1), .S(P2_P1_State2_PTR0), .Z(_03103__PTR19) );
  MUX2_X1 U23950 ( .A(_02186__PTR32), .B(1'b1), .S(P2_P1_State2_PTR0), .Z(_03102__PTR32) );
  MUX2_X1 U23951 ( .A(_03106__PTR32), .B(_03106__PTR128), .S(P2_P1_State2_PTR1), .Z(_03107__PTR0) );
  MUX2_X1 U23952 ( .A(_03106__PTR32), .B(_03106__PTR129), .S(P2_P1_State2_PTR1), .Z(_03107__PTR1) );
  MUX2_X1 U23953 ( .A(_03106__PTR32), .B(_03106__PTR130), .S(P2_P1_State2_PTR1), .Z(_03107__PTR2) );
  MUX2_X1 U23954 ( .A(_03106__PTR32), .B(_03106__PTR131), .S(P2_P1_State2_PTR1), .Z(_03107__PTR3) );
  MUX2_X1 U23955 ( .A(_03106__PTR19), .B(_03106__PTR132), .S(P2_P1_State2_PTR1), .Z(_03107__PTR4) );
  MUX2_X1 U23956 ( .A(_03106__PTR19), .B(_03106__PTR133), .S(P2_P1_State2_PTR1), .Z(_03107__PTR5) );
  MUX2_X1 U23957 ( .A(_03106__PTR19), .B(_03106__PTR134), .S(P2_P1_State2_PTR1), .Z(_03107__PTR6) );
  MUX2_X1 U23958 ( .A(_03106__PTR19), .B(_03106__PTR135), .S(P2_P1_State2_PTR1), .Z(_03107__PTR7) );
  MUX2_X1 U23959 ( .A(_03106__PTR19), .B(_03106__PTR136), .S(P2_P1_State2_PTR1), .Z(_03107__PTR8) );
  MUX2_X1 U23960 ( .A(_03106__PTR19), .B(_03106__PTR137), .S(P2_P1_State2_PTR1), .Z(_03107__PTR9) );
  MUX2_X1 U23961 ( .A(_03106__PTR19), .B(_03106__PTR138), .S(P2_P1_State2_PTR1), .Z(_03107__PTR10) );
  MUX2_X1 U23962 ( .A(_03106__PTR19), .B(_03106__PTR139), .S(P2_P1_State2_PTR1), .Z(_03107__PTR11) );
  MUX2_X1 U23963 ( .A(_03106__PTR19), .B(_03106__PTR140), .S(P2_P1_State2_PTR1), .Z(_03107__PTR12) );
  MUX2_X1 U23964 ( .A(_03106__PTR19), .B(_03106__PTR141), .S(P2_P1_State2_PTR1), .Z(_03107__PTR13) );
  MUX2_X1 U23965 ( .A(_03106__PTR19), .B(_03106__PTR142), .S(P2_P1_State2_PTR1), .Z(_03107__PTR14) );
  MUX2_X1 U23966 ( .A(_03106__PTR19), .B(_03106__PTR143), .S(P2_P1_State2_PTR1), .Z(_03107__PTR15) );
  MUX2_X1 U23967 ( .A(_03106__PTR19), .B(_03106__PTR144), .S(P2_P1_State2_PTR1), .Z(_03107__PTR16) );
  MUX2_X1 U23968 ( .A(_03106__PTR19), .B(_03106__PTR145), .S(P2_P1_State2_PTR1), .Z(_03107__PTR17) );
  MUX2_X1 U23969 ( .A(_03106__PTR19), .B(_03106__PTR146), .S(P2_P1_State2_PTR1), .Z(_03107__PTR18) );
  MUX2_X1 U23970 ( .A(_03106__PTR19), .B(_03106__PTR147), .S(P2_P1_State2_PTR1), .Z(_03107__PTR19) );
  MUX2_X1 U23971 ( .A(_03106__PTR32), .B(_03106__PTR148), .S(P2_P1_State2_PTR1), .Z(_03107__PTR20) );
  MUX2_X1 U23972 ( .A(_03106__PTR32), .B(_03106__PTR149), .S(P2_P1_State2_PTR1), .Z(_03107__PTR21) );
  MUX2_X1 U23973 ( .A(_03106__PTR32), .B(_03106__PTR150), .S(P2_P1_State2_PTR1), .Z(_03107__PTR22) );
  MUX2_X1 U23974 ( .A(_03106__PTR32), .B(_03106__PTR151), .S(P2_P1_State2_PTR1), .Z(_03107__PTR23) );
  MUX2_X1 U23975 ( .A(_03106__PTR32), .B(_03106__PTR152), .S(P2_P1_State2_PTR1), .Z(_03107__PTR24) );
  MUX2_X1 U23976 ( .A(_03106__PTR32), .B(_03106__PTR153), .S(P2_P1_State2_PTR1), .Z(_03107__PTR25) );
  MUX2_X1 U23977 ( .A(_03106__PTR32), .B(_03106__PTR154), .S(P2_P1_State2_PTR1), .Z(_03107__PTR26) );
  MUX2_X1 U23978 ( .A(_03106__PTR32), .B(_03106__PTR155), .S(P2_P1_State2_PTR1), .Z(_03107__PTR27) );
  MUX2_X1 U23979 ( .A(_03106__PTR32), .B(_03106__PTR156), .S(P2_P1_State2_PTR1), .Z(_03107__PTR28) );
  MUX2_X1 U23980 ( .A(_03106__PTR32), .B(_03106__PTR157), .S(P2_P1_State2_PTR1), .Z(_03107__PTR29) );
  MUX2_X1 U23981 ( .A(_03106__PTR32), .B(_03106__PTR158), .S(P2_P1_State2_PTR1), .Z(_03107__PTR30) );
  MUX2_X1 U23982 ( .A(_03106__PTR32), .B(_03106__PTR160), .S(P2_P1_State2_PTR1), .Z(_03107__PTR32) );
  MUX2_X1 U23983 ( .A(_03106__PTR256), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR256) );
  MUX2_X1 U23984 ( .A(_03106__PTR257), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR257) );
  MUX2_X1 U23985 ( .A(_03106__PTR258), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR258) );
  MUX2_X1 U23986 ( .A(_03106__PTR259), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR259) );
  MUX2_X1 U23987 ( .A(_03106__PTR260), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR260) );
  MUX2_X1 U23988 ( .A(_03106__PTR261), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR261) );
  MUX2_X1 U23989 ( .A(_03106__PTR262), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR262) );
  MUX2_X1 U23990 ( .A(_03106__PTR263), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR263) );
  MUX2_X1 U23991 ( .A(_03106__PTR264), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR264) );
  MUX2_X1 U23992 ( .A(_03106__PTR265), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR265) );
  MUX2_X1 U23993 ( .A(_03106__PTR266), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR266) );
  MUX2_X1 U23994 ( .A(_03106__PTR267), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR267) );
  MUX2_X1 U23995 ( .A(_03106__PTR268), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR268) );
  MUX2_X1 U23996 ( .A(_03106__PTR269), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR269) );
  MUX2_X1 U23997 ( .A(_03106__PTR270), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR270) );
  MUX2_X1 U23998 ( .A(_03106__PTR271), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR271) );
  MUX2_X1 U23999 ( .A(_03106__PTR272), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR272) );
  MUX2_X1 U24000 ( .A(_03106__PTR273), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR273) );
  MUX2_X1 U24001 ( .A(_03106__PTR274), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR274) );
  MUX2_X1 U24002 ( .A(_03106__PTR275), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR275) );
  MUX2_X1 U24003 ( .A(_03106__PTR276), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR276) );
  MUX2_X1 U24004 ( .A(_03106__PTR277), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR277) );
  MUX2_X1 U24005 ( .A(_03106__PTR278), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR278) );
  MUX2_X1 U24006 ( .A(_03106__PTR279), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR279) );
  MUX2_X1 U24007 ( .A(_03106__PTR280), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR280) );
  MUX2_X1 U24008 ( .A(_03106__PTR281), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR281) );
  MUX2_X1 U24009 ( .A(_03106__PTR282), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR282) );
  MUX2_X1 U24010 ( .A(_03106__PTR283), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR283) );
  MUX2_X1 U24011 ( .A(_03106__PTR284), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR284) );
  MUX2_X1 U24012 ( .A(_03106__PTR285), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR285) );
  MUX2_X1 U24013 ( .A(_03106__PTR286), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR286) );
  MUX2_X1 U24014 ( .A(_03106__PTR288), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03107__PTR288) );
  MUX2_X1 U24015 ( .A(1'b0), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR32) );
  MUX2_X1 U24016 ( .A(1'b1), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR19) );
  MUX2_X1 U24017 ( .A(_02188__PTR128), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR128) );
  MUX2_X1 U24018 ( .A(_02188__PTR129), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR129) );
  MUX2_X1 U24019 ( .A(_02188__PTR130), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR130) );
  MUX2_X1 U24020 ( .A(_02188__PTR131), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR131) );
  MUX2_X1 U24021 ( .A(_02188__PTR132), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR132) );
  MUX2_X1 U24022 ( .A(_02188__PTR133), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR133) );
  MUX2_X1 U24023 ( .A(_02188__PTR134), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR134) );
  MUX2_X1 U24024 ( .A(_02188__PTR135), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR135) );
  MUX2_X1 U24025 ( .A(_02188__PTR136), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR136) );
  MUX2_X1 U24026 ( .A(_02188__PTR137), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR137) );
  MUX2_X1 U24027 ( .A(_02188__PTR138), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR138) );
  MUX2_X1 U24028 ( .A(_02188__PTR139), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR139) );
  MUX2_X1 U24029 ( .A(_02188__PTR140), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR140) );
  MUX2_X1 U24030 ( .A(_02188__PTR141), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR141) );
  MUX2_X1 U24031 ( .A(_02188__PTR142), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR142) );
  MUX2_X1 U24032 ( .A(_02188__PTR143), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR143) );
  MUX2_X1 U24033 ( .A(_02188__PTR144), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR144) );
  MUX2_X1 U24034 ( .A(_02188__PTR145), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR145) );
  MUX2_X1 U24035 ( .A(_02188__PTR146), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR146) );
  MUX2_X1 U24036 ( .A(_02188__PTR147), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR147) );
  MUX2_X1 U24037 ( .A(_02188__PTR148), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR148) );
  MUX2_X1 U24038 ( .A(_02188__PTR149), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR149) );
  MUX2_X1 U24039 ( .A(_02188__PTR150), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR150) );
  MUX2_X1 U24040 ( .A(_02188__PTR151), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR151) );
  MUX2_X1 U24041 ( .A(_02188__PTR152), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR152) );
  MUX2_X1 U24042 ( .A(_02188__PTR153), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR153) );
  MUX2_X1 U24043 ( .A(_02188__PTR154), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR154) );
  MUX2_X1 U24044 ( .A(_02188__PTR155), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR155) );
  MUX2_X1 U24045 ( .A(_02188__PTR156), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR156) );
  MUX2_X1 U24046 ( .A(_02188__PTR157), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR157) );
  MUX2_X1 U24047 ( .A(_02188__PTR158), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR158) );
  MUX2_X1 U24048 ( .A(_02188__PTR160), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03106__PTR160) );
  MUX2_X1 U24049 ( .A(1'b0), .B(_02188__PTR320), .S(P2_P1_State2_PTR0), .Z(_03106__PTR256) );
  MUX2_X1 U24050 ( .A(1'b0), .B(_02188__PTR321), .S(P2_P1_State2_PTR0), .Z(_03106__PTR257) );
  MUX2_X1 U24051 ( .A(1'b0), .B(_02188__PTR322), .S(P2_P1_State2_PTR0), .Z(_03106__PTR258) );
  MUX2_X1 U24052 ( .A(1'b0), .B(_02188__PTR323), .S(P2_P1_State2_PTR0), .Z(_03106__PTR259) );
  MUX2_X1 U24053 ( .A(1'b0), .B(_02188__PTR324), .S(P2_P1_State2_PTR0), .Z(_03106__PTR260) );
  MUX2_X1 U24054 ( .A(1'b0), .B(_02188__PTR325), .S(P2_P1_State2_PTR0), .Z(_03106__PTR261) );
  MUX2_X1 U24055 ( .A(1'b0), .B(_02188__PTR326), .S(P2_P1_State2_PTR0), .Z(_03106__PTR262) );
  MUX2_X1 U24056 ( .A(1'b0), .B(_02188__PTR327), .S(P2_P1_State2_PTR0), .Z(_03106__PTR263) );
  MUX2_X1 U24057 ( .A(1'b0), .B(_02188__PTR328), .S(P2_P1_State2_PTR0), .Z(_03106__PTR264) );
  MUX2_X1 U24058 ( .A(1'b0), .B(_02188__PTR329), .S(P2_P1_State2_PTR0), .Z(_03106__PTR265) );
  MUX2_X1 U24059 ( .A(1'b0), .B(_02188__PTR330), .S(P2_P1_State2_PTR0), .Z(_03106__PTR266) );
  MUX2_X1 U24060 ( .A(1'b0), .B(_02188__PTR331), .S(P2_P1_State2_PTR0), .Z(_03106__PTR267) );
  MUX2_X1 U24061 ( .A(1'b0), .B(_02188__PTR332), .S(P2_P1_State2_PTR0), .Z(_03106__PTR268) );
  MUX2_X1 U24062 ( .A(1'b0), .B(_02188__PTR333), .S(P2_P1_State2_PTR0), .Z(_03106__PTR269) );
  MUX2_X1 U24063 ( .A(1'b0), .B(_02188__PTR334), .S(P2_P1_State2_PTR0), .Z(_03106__PTR270) );
  MUX2_X1 U24064 ( .A(1'b0), .B(_02188__PTR335), .S(P2_P1_State2_PTR0), .Z(_03106__PTR271) );
  MUX2_X1 U24065 ( .A(1'b0), .B(_02188__PTR336), .S(P2_P1_State2_PTR0), .Z(_03106__PTR272) );
  MUX2_X1 U24066 ( .A(1'b0), .B(_02188__PTR337), .S(P2_P1_State2_PTR0), .Z(_03106__PTR273) );
  MUX2_X1 U24067 ( .A(1'b0), .B(_02188__PTR338), .S(P2_P1_State2_PTR0), .Z(_03106__PTR274) );
  MUX2_X1 U24068 ( .A(1'b0), .B(_02188__PTR339), .S(P2_P1_State2_PTR0), .Z(_03106__PTR275) );
  MUX2_X1 U24069 ( .A(1'b0), .B(_02188__PTR340), .S(P2_P1_State2_PTR0), .Z(_03106__PTR276) );
  MUX2_X1 U24070 ( .A(1'b0), .B(_02188__PTR341), .S(P2_P1_State2_PTR0), .Z(_03106__PTR277) );
  MUX2_X1 U24071 ( .A(1'b0), .B(_02188__PTR342), .S(P2_P1_State2_PTR0), .Z(_03106__PTR278) );
  MUX2_X1 U24072 ( .A(1'b0), .B(_02188__PTR343), .S(P2_P1_State2_PTR0), .Z(_03106__PTR279) );
  MUX2_X1 U24073 ( .A(1'b0), .B(_02188__PTR344), .S(P2_P1_State2_PTR0), .Z(_03106__PTR280) );
  MUX2_X1 U24074 ( .A(1'b0), .B(_02188__PTR345), .S(P2_P1_State2_PTR0), .Z(_03106__PTR281) );
  MUX2_X1 U24075 ( .A(1'b0), .B(_02188__PTR346), .S(P2_P1_State2_PTR0), .Z(_03106__PTR282) );
  MUX2_X1 U24076 ( .A(1'b0), .B(_02188__PTR347), .S(P2_P1_State2_PTR0), .Z(_03106__PTR283) );
  MUX2_X1 U24077 ( .A(1'b0), .B(_02188__PTR348), .S(P2_P1_State2_PTR0), .Z(_03106__PTR284) );
  MUX2_X1 U24078 ( .A(1'b0), .B(_02188__PTR349), .S(P2_P1_State2_PTR0), .Z(_03106__PTR285) );
  MUX2_X1 U24079 ( .A(1'b0), .B(_02188__PTR350), .S(P2_P1_State2_PTR0), .Z(_03106__PTR286) );
  MUX2_X1 U24080 ( .A(1'b0), .B(_02188__PTR352), .S(P2_P1_State2_PTR0), .Z(_03106__PTR288) );
  MUX2_X1 U24081 ( .A(_03108__PTR0), .B(_03096__PTR0), .S(P2_P1_State2_PTR3), .Z(_02189__PTR0) );
  MUX2_X1 U24082 ( .A(_03108__PTR1), .B(_03096__PTR1), .S(P2_P1_State2_PTR3), .Z(_02189__PTR1) );
  MUX2_X1 U24083 ( .A(_03108__PTR2), .B(_03096__PTR2), .S(P2_P1_State2_PTR3), .Z(_02189__PTR2) );
  MUX2_X1 U24084 ( .A(_03108__PTR3), .B(_03096__PTR3), .S(P2_P1_State2_PTR3), .Z(_02189__PTR3) );
  MUX2_X1 U24085 ( .A(_03108__PTR4), .B(_03096__PTR4), .S(P2_P1_State2_PTR3), .Z(_02189__PTR4) );
  MUX2_X1 U24086 ( .A(_03108__PTR5), .B(_03096__PTR5), .S(P2_P1_State2_PTR3), .Z(_02189__PTR5) );
  MUX2_X1 U24087 ( .A(_03108__PTR6), .B(_03096__PTR6), .S(P2_P1_State2_PTR3), .Z(_02189__PTR6) );
  MUX2_X1 U24088 ( .A(_03108__PTR7), .B(_03096__PTR7), .S(P2_P1_State2_PTR3), .Z(_02189__PTR7) );
  MUX2_X1 U24089 ( .A(_03108__PTR8), .B(_03096__PTR8), .S(P2_P1_State2_PTR3), .Z(_02189__PTR8) );
  MUX2_X1 U24090 ( .A(_03108__PTR9), .B(_03096__PTR9), .S(P2_P1_State2_PTR3), .Z(_02189__PTR9) );
  MUX2_X1 U24091 ( .A(_03108__PTR10), .B(_03096__PTR10), .S(P2_P1_State2_PTR3), .Z(_02189__PTR10) );
  MUX2_X1 U24092 ( .A(_03108__PTR11), .B(_03096__PTR11), .S(P2_P1_State2_PTR3), .Z(_02189__PTR11) );
  MUX2_X1 U24093 ( .A(_03108__PTR12), .B(_03096__PTR12), .S(P2_P1_State2_PTR3), .Z(_02189__PTR12) );
  MUX2_X1 U24094 ( .A(_03108__PTR13), .B(_03096__PTR13), .S(P2_P1_State2_PTR3), .Z(_02189__PTR13) );
  MUX2_X1 U24095 ( .A(_03108__PTR14), .B(_03096__PTR14), .S(P2_P1_State2_PTR3), .Z(_02189__PTR14) );
  MUX2_X1 U24096 ( .A(_03108__PTR15), .B(_03096__PTR15), .S(P2_P1_State2_PTR3), .Z(_02189__PTR15) );
  MUX2_X1 U24097 ( .A(_03108__PTR16), .B(_03096__PTR16), .S(P2_P1_State2_PTR3), .Z(_02189__PTR16) );
  MUX2_X1 U24098 ( .A(_03108__PTR17), .B(_03096__PTR17), .S(P2_P1_State2_PTR3), .Z(_02189__PTR17) );
  MUX2_X1 U24099 ( .A(_03108__PTR18), .B(_03096__PTR18), .S(P2_P1_State2_PTR3), .Z(_02189__PTR18) );
  MUX2_X1 U24100 ( .A(_03108__PTR19), .B(_03096__PTR19), .S(P2_P1_State2_PTR3), .Z(_02189__PTR19) );
  MUX2_X1 U24101 ( .A(_03108__PTR20), .B(_03096__PTR20), .S(P2_P1_State2_PTR3), .Z(_02189__PTR20) );
  MUX2_X1 U24102 ( .A(_03108__PTR21), .B(_03096__PTR21), .S(P2_P1_State2_PTR3), .Z(_02189__PTR21) );
  MUX2_X1 U24103 ( .A(_03108__PTR22), .B(_03096__PTR22), .S(P2_P1_State2_PTR3), .Z(_02189__PTR22) );
  MUX2_X1 U24104 ( .A(_03108__PTR23), .B(_03096__PTR23), .S(P2_P1_State2_PTR3), .Z(_02189__PTR23) );
  MUX2_X1 U24105 ( .A(_03108__PTR24), .B(_03096__PTR24), .S(P2_P1_State2_PTR3), .Z(_02189__PTR24) );
  MUX2_X1 U24106 ( .A(_03108__PTR25), .B(_03096__PTR25), .S(P2_P1_State2_PTR3), .Z(_02189__PTR25) );
  MUX2_X1 U24107 ( .A(_03108__PTR26), .B(_03096__PTR26), .S(P2_P1_State2_PTR3), .Z(_02189__PTR26) );
  MUX2_X1 U24108 ( .A(_03108__PTR27), .B(_03096__PTR27), .S(P2_P1_State2_PTR3), .Z(_02189__PTR27) );
  MUX2_X1 U24109 ( .A(_03108__PTR28), .B(_03096__PTR28), .S(P2_P1_State2_PTR3), .Z(_02189__PTR28) );
  MUX2_X1 U24110 ( .A(_03108__PTR29), .B(_03096__PTR29), .S(P2_P1_State2_PTR3), .Z(_02189__PTR29) );
  MUX2_X1 U24111 ( .A(_03108__PTR30), .B(_03096__PTR30), .S(P2_P1_State2_PTR3), .Z(_02189__PTR30) );
  MUX2_X1 U24112 ( .A(_03108__PTR32), .B(_03096__PTR31), .S(P2_P1_State2_PTR3), .Z(_02189__PTR32) );
  MUX2_X1 U24113 ( .A(_03107__PTR0), .B(_03107__PTR256), .S(P2_P1_State2_PTR2), .Z(_03108__PTR0) );
  MUX2_X1 U24114 ( .A(_03107__PTR1), .B(_03107__PTR257), .S(P2_P1_State2_PTR2), .Z(_03108__PTR1) );
  MUX2_X1 U24115 ( .A(_03107__PTR2), .B(_03107__PTR258), .S(P2_P1_State2_PTR2), .Z(_03108__PTR2) );
  MUX2_X1 U24116 ( .A(_03107__PTR3), .B(_03107__PTR259), .S(P2_P1_State2_PTR2), .Z(_03108__PTR3) );
  MUX2_X1 U24117 ( .A(_03107__PTR4), .B(_03107__PTR260), .S(P2_P1_State2_PTR2), .Z(_03108__PTR4) );
  MUX2_X1 U24118 ( .A(_03107__PTR5), .B(_03107__PTR261), .S(P2_P1_State2_PTR2), .Z(_03108__PTR5) );
  MUX2_X1 U24119 ( .A(_03107__PTR6), .B(_03107__PTR262), .S(P2_P1_State2_PTR2), .Z(_03108__PTR6) );
  MUX2_X1 U24120 ( .A(_03107__PTR7), .B(_03107__PTR263), .S(P2_P1_State2_PTR2), .Z(_03108__PTR7) );
  MUX2_X1 U24121 ( .A(_03107__PTR8), .B(_03107__PTR264), .S(P2_P1_State2_PTR2), .Z(_03108__PTR8) );
  MUX2_X1 U24122 ( .A(_03107__PTR9), .B(_03107__PTR265), .S(P2_P1_State2_PTR2), .Z(_03108__PTR9) );
  MUX2_X1 U24123 ( .A(_03107__PTR10), .B(_03107__PTR266), .S(P2_P1_State2_PTR2), .Z(_03108__PTR10) );
  MUX2_X1 U24124 ( .A(_03107__PTR11), .B(_03107__PTR267), .S(P2_P1_State2_PTR2), .Z(_03108__PTR11) );
  MUX2_X1 U24125 ( .A(_03107__PTR12), .B(_03107__PTR268), .S(P2_P1_State2_PTR2), .Z(_03108__PTR12) );
  MUX2_X1 U24126 ( .A(_03107__PTR13), .B(_03107__PTR269), .S(P2_P1_State2_PTR2), .Z(_03108__PTR13) );
  MUX2_X1 U24127 ( .A(_03107__PTR14), .B(_03107__PTR270), .S(P2_P1_State2_PTR2), .Z(_03108__PTR14) );
  MUX2_X1 U24128 ( .A(_03107__PTR15), .B(_03107__PTR271), .S(P2_P1_State2_PTR2), .Z(_03108__PTR15) );
  MUX2_X1 U24129 ( .A(_03107__PTR16), .B(_03107__PTR272), .S(P2_P1_State2_PTR2), .Z(_03108__PTR16) );
  MUX2_X1 U24130 ( .A(_03107__PTR17), .B(_03107__PTR273), .S(P2_P1_State2_PTR2), .Z(_03108__PTR17) );
  MUX2_X1 U24131 ( .A(_03107__PTR18), .B(_03107__PTR274), .S(P2_P1_State2_PTR2), .Z(_03108__PTR18) );
  MUX2_X1 U24132 ( .A(_03107__PTR19), .B(_03107__PTR275), .S(P2_P1_State2_PTR2), .Z(_03108__PTR19) );
  MUX2_X1 U24133 ( .A(_03107__PTR20), .B(_03107__PTR276), .S(P2_P1_State2_PTR2), .Z(_03108__PTR20) );
  MUX2_X1 U24134 ( .A(_03107__PTR21), .B(_03107__PTR277), .S(P2_P1_State2_PTR2), .Z(_03108__PTR21) );
  MUX2_X1 U24135 ( .A(_03107__PTR22), .B(_03107__PTR278), .S(P2_P1_State2_PTR2), .Z(_03108__PTR22) );
  MUX2_X1 U24136 ( .A(_03107__PTR23), .B(_03107__PTR279), .S(P2_P1_State2_PTR2), .Z(_03108__PTR23) );
  MUX2_X1 U24137 ( .A(_03107__PTR24), .B(_03107__PTR280), .S(P2_P1_State2_PTR2), .Z(_03108__PTR24) );
  MUX2_X1 U24138 ( .A(_03107__PTR25), .B(_03107__PTR281), .S(P2_P1_State2_PTR2), .Z(_03108__PTR25) );
  MUX2_X1 U24139 ( .A(_03107__PTR26), .B(_03107__PTR282), .S(P2_P1_State2_PTR2), .Z(_03108__PTR26) );
  MUX2_X1 U24140 ( .A(_03107__PTR27), .B(_03107__PTR283), .S(P2_P1_State2_PTR2), .Z(_03108__PTR27) );
  MUX2_X1 U24141 ( .A(_03107__PTR28), .B(_03107__PTR284), .S(P2_P1_State2_PTR2), .Z(_03108__PTR28) );
  MUX2_X1 U24142 ( .A(_03107__PTR29), .B(_03107__PTR285), .S(P2_P1_State2_PTR2), .Z(_03108__PTR29) );
  MUX2_X1 U24143 ( .A(_03107__PTR30), .B(_03107__PTR286), .S(P2_P1_State2_PTR2), .Z(_03108__PTR30) );
  MUX2_X1 U24144 ( .A(_03107__PTR32), .B(_03107__PTR288), .S(P2_P1_State2_PTR2), .Z(_03108__PTR32) );
  MUX2_X1 U24145 ( .A(_03111__PTR0), .B(_03109__PTR64), .S(P2_P1_State2_PTR3), .Z(_02191__PTR0) );
  MUX2_X1 U24146 ( .A(_03111__PTR1), .B(_03109__PTR65), .S(P2_P1_State2_PTR3), .Z(_02191__PTR1) );
  MUX2_X1 U24147 ( .A(_03111__PTR2), .B(_03109__PTR66), .S(P2_P1_State2_PTR3), .Z(_02191__PTR2) );
  MUX2_X1 U24148 ( .A(_03111__PTR3), .B(_03109__PTR67), .S(P2_P1_State2_PTR3), .Z(_02191__PTR3) );
  MUX2_X1 U24149 ( .A(_03111__PTR4), .B(_03109__PTR68), .S(P2_P1_State2_PTR3), .Z(_02191__PTR4) );
  MUX2_X1 U24150 ( .A(_03111__PTR5), .B(_03109__PTR69), .S(P2_P1_State2_PTR3), .Z(_02191__PTR5) );
  MUX2_X1 U24151 ( .A(_03111__PTR6), .B(_03109__PTR70), .S(P2_P1_State2_PTR3), .Z(_02191__PTR6) );
  MUX2_X1 U24152 ( .A(_03111__PTR7), .B(_03109__PTR71), .S(P2_P1_State2_PTR3), .Z(_02191__PTR7) );
  MUX2_X1 U24153 ( .A(_03110__PTR0), .B(_03110__PTR32), .S(P2_P1_State2_PTR2), .Z(_03111__PTR0) );
  MUX2_X1 U24154 ( .A(_03110__PTR1), .B(_03110__PTR33), .S(P2_P1_State2_PTR2), .Z(_03111__PTR1) );
  MUX2_X1 U24155 ( .A(_03110__PTR2), .B(_03110__PTR34), .S(P2_P1_State2_PTR2), .Z(_03111__PTR2) );
  MUX2_X1 U24156 ( .A(_03110__PTR3), .B(_03110__PTR35), .S(P2_P1_State2_PTR2), .Z(_03111__PTR3) );
  MUX2_X1 U24157 ( .A(_03110__PTR4), .B(_03110__PTR36), .S(P2_P1_State2_PTR2), .Z(_03111__PTR4) );
  MUX2_X1 U24158 ( .A(_03110__PTR5), .B(_03110__PTR37), .S(P2_P1_State2_PTR2), .Z(_03111__PTR5) );
  MUX2_X1 U24159 ( .A(_03110__PTR6), .B(_03110__PTR38), .S(P2_P1_State2_PTR2), .Z(_03111__PTR6) );
  MUX2_X1 U24160 ( .A(_03110__PTR7), .B(_03110__PTR39), .S(P2_P1_State2_PTR2), .Z(_03111__PTR7) );
  MUX2_X1 U24161 ( .A(1'b0), .B(_03109__PTR16), .S(P2_P1_State2_PTR1), .Z(_03110__PTR0) );
  MUX2_X1 U24162 ( .A(1'b0), .B(_03109__PTR17), .S(P2_P1_State2_PTR1), .Z(_03110__PTR1) );
  MUX2_X1 U24163 ( .A(1'b0), .B(_03109__PTR18), .S(P2_P1_State2_PTR1), .Z(_03110__PTR2) );
  MUX2_X1 U24164 ( .A(1'b0), .B(_03109__PTR19), .S(P2_P1_State2_PTR1), .Z(_03110__PTR3) );
  MUX2_X1 U24165 ( .A(1'b0), .B(_03109__PTR20), .S(P2_P1_State2_PTR1), .Z(_03110__PTR4) );
  MUX2_X1 U24166 ( .A(1'b0), .B(_03109__PTR21), .S(P2_P1_State2_PTR1), .Z(_03110__PTR5) );
  MUX2_X1 U24167 ( .A(1'b0), .B(_03109__PTR22), .S(P2_P1_State2_PTR1), .Z(_03110__PTR6) );
  MUX2_X1 U24168 ( .A(1'b0), .B(_03109__PTR23), .S(P2_P1_State2_PTR1), .Z(_03110__PTR7) );
  MUX2_X1 U24169 ( .A(_03109__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03110__PTR32) );
  MUX2_X1 U24170 ( .A(_03109__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03110__PTR33) );
  MUX2_X1 U24171 ( .A(_03109__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03110__PTR34) );
  MUX2_X1 U24172 ( .A(_03109__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03110__PTR35) );
  MUX2_X1 U24173 ( .A(_03109__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03110__PTR36) );
  MUX2_X1 U24174 ( .A(_03109__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03110__PTR37) );
  MUX2_X1 U24175 ( .A(_03109__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03110__PTR38) );
  MUX2_X1 U24176 ( .A(_03109__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03110__PTR39) );
  MUX2_X1 U24177 ( .A(_02190__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR16) );
  MUX2_X1 U24178 ( .A(_02190__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR17) );
  MUX2_X1 U24179 ( .A(_02190__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR18) );
  MUX2_X1 U24180 ( .A(_02190__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR19) );
  MUX2_X1 U24181 ( .A(_02190__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR20) );
  MUX2_X1 U24182 ( .A(_02190__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR21) );
  MUX2_X1 U24183 ( .A(_02190__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR22) );
  MUX2_X1 U24184 ( .A(_02190__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR23) );
  MUX2_X1 U24185 ( .A(_02190__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR32) );
  MUX2_X1 U24186 ( .A(_02190__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR33) );
  MUX2_X1 U24187 ( .A(_02190__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR34) );
  MUX2_X1 U24188 ( .A(_02190__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR35) );
  MUX2_X1 U24189 ( .A(_02190__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR36) );
  MUX2_X1 U24190 ( .A(_02190__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR37) );
  MUX2_X1 U24191 ( .A(_02190__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR38) );
  MUX2_X1 U24192 ( .A(_02190__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR39) );
  MUX2_X1 U24193 ( .A(_02190__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR64) );
  MUX2_X1 U24194 ( .A(_02190__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR65) );
  MUX2_X1 U24195 ( .A(_02190__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR66) );
  MUX2_X1 U24196 ( .A(_02190__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR67) );
  MUX2_X1 U24197 ( .A(_02190__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR68) );
  MUX2_X1 U24198 ( .A(_02190__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR69) );
  MUX2_X1 U24199 ( .A(_02190__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR70) );
  MUX2_X1 U24200 ( .A(_02190__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03109__PTR71) );
  MUX2_X1 U24201 ( .A(_03114__PTR0), .B(_03112__PTR64), .S(P2_P1_State2_PTR3), .Z(_02193__PTR0) );
  MUX2_X1 U24202 ( .A(_03114__PTR1), .B(_03112__PTR65), .S(P2_P1_State2_PTR3), .Z(_02193__PTR1) );
  MUX2_X1 U24203 ( .A(_03114__PTR2), .B(_03112__PTR66), .S(P2_P1_State2_PTR3), .Z(_02193__PTR2) );
  MUX2_X1 U24204 ( .A(_03114__PTR3), .B(_03112__PTR67), .S(P2_P1_State2_PTR3), .Z(_02193__PTR3) );
  MUX2_X1 U24205 ( .A(_03114__PTR4), .B(_03112__PTR68), .S(P2_P1_State2_PTR3), .Z(_02193__PTR4) );
  MUX2_X1 U24206 ( .A(_03114__PTR5), .B(_03112__PTR69), .S(P2_P1_State2_PTR3), .Z(_02193__PTR5) );
  MUX2_X1 U24207 ( .A(_03114__PTR6), .B(_03112__PTR70), .S(P2_P1_State2_PTR3), .Z(_02193__PTR6) );
  MUX2_X1 U24208 ( .A(_03114__PTR7), .B(_03112__PTR71), .S(P2_P1_State2_PTR3), .Z(_02193__PTR7) );
  MUX2_X1 U24209 ( .A(_03113__PTR0), .B(_03113__PTR32), .S(P2_P1_State2_PTR2), .Z(_03114__PTR0) );
  MUX2_X1 U24210 ( .A(_03113__PTR1), .B(_03113__PTR33), .S(P2_P1_State2_PTR2), .Z(_03114__PTR1) );
  MUX2_X1 U24211 ( .A(_03113__PTR2), .B(_03113__PTR34), .S(P2_P1_State2_PTR2), .Z(_03114__PTR2) );
  MUX2_X1 U24212 ( .A(_03113__PTR3), .B(_03113__PTR35), .S(P2_P1_State2_PTR2), .Z(_03114__PTR3) );
  MUX2_X1 U24213 ( .A(_03113__PTR4), .B(_03113__PTR36), .S(P2_P1_State2_PTR2), .Z(_03114__PTR4) );
  MUX2_X1 U24214 ( .A(_03113__PTR5), .B(_03113__PTR37), .S(P2_P1_State2_PTR2), .Z(_03114__PTR5) );
  MUX2_X1 U24215 ( .A(_03113__PTR6), .B(_03113__PTR38), .S(P2_P1_State2_PTR2), .Z(_03114__PTR6) );
  MUX2_X1 U24216 ( .A(_03113__PTR7), .B(_03113__PTR39), .S(P2_P1_State2_PTR2), .Z(_03114__PTR7) );
  MUX2_X1 U24217 ( .A(1'b0), .B(_03112__PTR16), .S(P2_P1_State2_PTR1), .Z(_03113__PTR0) );
  MUX2_X1 U24218 ( .A(1'b0), .B(_03112__PTR17), .S(P2_P1_State2_PTR1), .Z(_03113__PTR1) );
  MUX2_X1 U24219 ( .A(1'b0), .B(_03112__PTR18), .S(P2_P1_State2_PTR1), .Z(_03113__PTR2) );
  MUX2_X1 U24220 ( .A(1'b0), .B(_03112__PTR19), .S(P2_P1_State2_PTR1), .Z(_03113__PTR3) );
  MUX2_X1 U24221 ( .A(1'b0), .B(_03112__PTR20), .S(P2_P1_State2_PTR1), .Z(_03113__PTR4) );
  MUX2_X1 U24222 ( .A(1'b0), .B(_03112__PTR21), .S(P2_P1_State2_PTR1), .Z(_03113__PTR5) );
  MUX2_X1 U24223 ( .A(1'b0), .B(_03112__PTR22), .S(P2_P1_State2_PTR1), .Z(_03113__PTR6) );
  MUX2_X1 U24224 ( .A(1'b0), .B(_03112__PTR23), .S(P2_P1_State2_PTR1), .Z(_03113__PTR7) );
  MUX2_X1 U24225 ( .A(_03112__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03113__PTR32) );
  MUX2_X1 U24226 ( .A(_03112__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03113__PTR33) );
  MUX2_X1 U24227 ( .A(_03112__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03113__PTR34) );
  MUX2_X1 U24228 ( .A(_03112__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03113__PTR35) );
  MUX2_X1 U24229 ( .A(_03112__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03113__PTR36) );
  MUX2_X1 U24230 ( .A(_03112__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03113__PTR37) );
  MUX2_X1 U24231 ( .A(_03112__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03113__PTR38) );
  MUX2_X1 U24232 ( .A(_03112__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03113__PTR39) );
  MUX2_X1 U24233 ( .A(_02192__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR16) );
  MUX2_X1 U24234 ( .A(_02192__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR17) );
  MUX2_X1 U24235 ( .A(_02192__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR18) );
  MUX2_X1 U24236 ( .A(_02192__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR19) );
  MUX2_X1 U24237 ( .A(_02192__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR20) );
  MUX2_X1 U24238 ( .A(_02192__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR21) );
  MUX2_X1 U24239 ( .A(_02192__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR22) );
  MUX2_X1 U24240 ( .A(_02192__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR23) );
  MUX2_X1 U24241 ( .A(_02192__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR32) );
  MUX2_X1 U24242 ( .A(_02192__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR33) );
  MUX2_X1 U24243 ( .A(_02192__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR34) );
  MUX2_X1 U24244 ( .A(_02192__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR35) );
  MUX2_X1 U24245 ( .A(_02192__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR36) );
  MUX2_X1 U24246 ( .A(_02192__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR37) );
  MUX2_X1 U24247 ( .A(_02192__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR38) );
  MUX2_X1 U24248 ( .A(_02192__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR39) );
  MUX2_X1 U24249 ( .A(_02192__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR64) );
  MUX2_X1 U24250 ( .A(_02192__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR65) );
  MUX2_X1 U24251 ( .A(_02192__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR66) );
  MUX2_X1 U24252 ( .A(_02192__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR67) );
  MUX2_X1 U24253 ( .A(_02192__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR68) );
  MUX2_X1 U24254 ( .A(_02192__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR69) );
  MUX2_X1 U24255 ( .A(_02192__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR70) );
  MUX2_X1 U24256 ( .A(_02192__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03112__PTR71) );
  MUX2_X1 U24257 ( .A(_03117__PTR0), .B(_03115__PTR64), .S(P2_P1_State2_PTR3), .Z(_02195__PTR0) );
  MUX2_X1 U24258 ( .A(_03117__PTR1), .B(_03115__PTR65), .S(P2_P1_State2_PTR3), .Z(_02195__PTR1) );
  MUX2_X1 U24259 ( .A(_03117__PTR2), .B(_03115__PTR66), .S(P2_P1_State2_PTR3), .Z(_02195__PTR2) );
  MUX2_X1 U24260 ( .A(_03117__PTR3), .B(_03115__PTR67), .S(P2_P1_State2_PTR3), .Z(_02195__PTR3) );
  MUX2_X1 U24261 ( .A(_03117__PTR4), .B(_03115__PTR68), .S(P2_P1_State2_PTR3), .Z(_02195__PTR4) );
  MUX2_X1 U24262 ( .A(_03117__PTR5), .B(_03115__PTR69), .S(P2_P1_State2_PTR3), .Z(_02195__PTR5) );
  MUX2_X1 U24263 ( .A(_03117__PTR6), .B(_03115__PTR70), .S(P2_P1_State2_PTR3), .Z(_02195__PTR6) );
  MUX2_X1 U24264 ( .A(_03117__PTR7), .B(_03115__PTR71), .S(P2_P1_State2_PTR3), .Z(_02195__PTR7) );
  MUX2_X1 U24265 ( .A(_03116__PTR0), .B(_03116__PTR32), .S(P2_P1_State2_PTR2), .Z(_03117__PTR0) );
  MUX2_X1 U24266 ( .A(_03116__PTR1), .B(_03116__PTR33), .S(P2_P1_State2_PTR2), .Z(_03117__PTR1) );
  MUX2_X1 U24267 ( .A(_03116__PTR2), .B(_03116__PTR34), .S(P2_P1_State2_PTR2), .Z(_03117__PTR2) );
  MUX2_X1 U24268 ( .A(_03116__PTR3), .B(_03116__PTR35), .S(P2_P1_State2_PTR2), .Z(_03117__PTR3) );
  MUX2_X1 U24269 ( .A(_03116__PTR4), .B(_03116__PTR36), .S(P2_P1_State2_PTR2), .Z(_03117__PTR4) );
  MUX2_X1 U24270 ( .A(_03116__PTR5), .B(_03116__PTR37), .S(P2_P1_State2_PTR2), .Z(_03117__PTR5) );
  MUX2_X1 U24271 ( .A(_03116__PTR6), .B(_03116__PTR38), .S(P2_P1_State2_PTR2), .Z(_03117__PTR6) );
  MUX2_X1 U24272 ( .A(_03116__PTR7), .B(_03116__PTR39), .S(P2_P1_State2_PTR2), .Z(_03117__PTR7) );
  MUX2_X1 U24273 ( .A(1'b0), .B(_03115__PTR16), .S(P2_P1_State2_PTR1), .Z(_03116__PTR0) );
  MUX2_X1 U24274 ( .A(1'b0), .B(_03115__PTR17), .S(P2_P1_State2_PTR1), .Z(_03116__PTR1) );
  MUX2_X1 U24275 ( .A(1'b0), .B(_03115__PTR18), .S(P2_P1_State2_PTR1), .Z(_03116__PTR2) );
  MUX2_X1 U24276 ( .A(1'b0), .B(_03115__PTR19), .S(P2_P1_State2_PTR1), .Z(_03116__PTR3) );
  MUX2_X1 U24277 ( .A(1'b0), .B(_03115__PTR20), .S(P2_P1_State2_PTR1), .Z(_03116__PTR4) );
  MUX2_X1 U24278 ( .A(1'b0), .B(_03115__PTR21), .S(P2_P1_State2_PTR1), .Z(_03116__PTR5) );
  MUX2_X1 U24279 ( .A(1'b0), .B(_03115__PTR22), .S(P2_P1_State2_PTR1), .Z(_03116__PTR6) );
  MUX2_X1 U24280 ( .A(1'b0), .B(_03115__PTR23), .S(P2_P1_State2_PTR1), .Z(_03116__PTR7) );
  MUX2_X1 U24281 ( .A(_03115__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03116__PTR32) );
  MUX2_X1 U24282 ( .A(_03115__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03116__PTR33) );
  MUX2_X1 U24283 ( .A(_03115__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03116__PTR34) );
  MUX2_X1 U24284 ( .A(_03115__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03116__PTR35) );
  MUX2_X1 U24285 ( .A(_03115__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03116__PTR36) );
  MUX2_X1 U24286 ( .A(_03115__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03116__PTR37) );
  MUX2_X1 U24287 ( .A(_03115__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03116__PTR38) );
  MUX2_X1 U24288 ( .A(_03115__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03116__PTR39) );
  MUX2_X1 U24289 ( .A(_02194__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR16) );
  MUX2_X1 U24290 ( .A(_02194__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR17) );
  MUX2_X1 U24291 ( .A(_02194__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR18) );
  MUX2_X1 U24292 ( .A(_02194__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR19) );
  MUX2_X1 U24293 ( .A(_02194__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR20) );
  MUX2_X1 U24294 ( .A(_02194__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR21) );
  MUX2_X1 U24295 ( .A(_02194__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR22) );
  MUX2_X1 U24296 ( .A(_02194__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR23) );
  MUX2_X1 U24297 ( .A(_02194__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR32) );
  MUX2_X1 U24298 ( .A(_02194__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR33) );
  MUX2_X1 U24299 ( .A(_02194__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR34) );
  MUX2_X1 U24300 ( .A(_02194__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR35) );
  MUX2_X1 U24301 ( .A(_02194__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR36) );
  MUX2_X1 U24302 ( .A(_02194__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR37) );
  MUX2_X1 U24303 ( .A(_02194__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR38) );
  MUX2_X1 U24304 ( .A(_02194__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR39) );
  MUX2_X1 U24305 ( .A(_02194__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR64) );
  MUX2_X1 U24306 ( .A(_02194__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR65) );
  MUX2_X1 U24307 ( .A(_02194__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR66) );
  MUX2_X1 U24308 ( .A(_02194__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR67) );
  MUX2_X1 U24309 ( .A(_02194__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR68) );
  MUX2_X1 U24310 ( .A(_02194__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR69) );
  MUX2_X1 U24311 ( .A(_02194__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR70) );
  MUX2_X1 U24312 ( .A(_02194__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03115__PTR71) );
  MUX2_X1 U24313 ( .A(_03120__PTR0), .B(_03118__PTR64), .S(P2_P1_State2_PTR3), .Z(_02197__PTR0) );
  MUX2_X1 U24314 ( .A(_03120__PTR1), .B(_03118__PTR65), .S(P2_P1_State2_PTR3), .Z(_02197__PTR1) );
  MUX2_X1 U24315 ( .A(_03120__PTR2), .B(_03118__PTR66), .S(P2_P1_State2_PTR3), .Z(_02197__PTR2) );
  MUX2_X1 U24316 ( .A(_03120__PTR3), .B(_03118__PTR67), .S(P2_P1_State2_PTR3), .Z(_02197__PTR3) );
  MUX2_X1 U24317 ( .A(_03120__PTR4), .B(_03118__PTR68), .S(P2_P1_State2_PTR3), .Z(_02197__PTR4) );
  MUX2_X1 U24318 ( .A(_03120__PTR5), .B(_03118__PTR69), .S(P2_P1_State2_PTR3), .Z(_02197__PTR5) );
  MUX2_X1 U24319 ( .A(_03120__PTR6), .B(_03118__PTR70), .S(P2_P1_State2_PTR3), .Z(_02197__PTR6) );
  MUX2_X1 U24320 ( .A(_03120__PTR7), .B(_03118__PTR71), .S(P2_P1_State2_PTR3), .Z(_02197__PTR7) );
  MUX2_X1 U24321 ( .A(_03119__PTR0), .B(_03119__PTR32), .S(P2_P1_State2_PTR2), .Z(_03120__PTR0) );
  MUX2_X1 U24322 ( .A(_03119__PTR1), .B(_03119__PTR33), .S(P2_P1_State2_PTR2), .Z(_03120__PTR1) );
  MUX2_X1 U24323 ( .A(_03119__PTR2), .B(_03119__PTR34), .S(P2_P1_State2_PTR2), .Z(_03120__PTR2) );
  MUX2_X1 U24324 ( .A(_03119__PTR3), .B(_03119__PTR35), .S(P2_P1_State2_PTR2), .Z(_03120__PTR3) );
  MUX2_X1 U24325 ( .A(_03119__PTR4), .B(_03119__PTR36), .S(P2_P1_State2_PTR2), .Z(_03120__PTR4) );
  MUX2_X1 U24326 ( .A(_03119__PTR5), .B(_03119__PTR37), .S(P2_P1_State2_PTR2), .Z(_03120__PTR5) );
  MUX2_X1 U24327 ( .A(_03119__PTR6), .B(_03119__PTR38), .S(P2_P1_State2_PTR2), .Z(_03120__PTR6) );
  MUX2_X1 U24328 ( .A(_03119__PTR7), .B(_03119__PTR39), .S(P2_P1_State2_PTR2), .Z(_03120__PTR7) );
  MUX2_X1 U24329 ( .A(1'b0), .B(_03118__PTR16), .S(P2_P1_State2_PTR1), .Z(_03119__PTR0) );
  MUX2_X1 U24330 ( .A(1'b0), .B(_03118__PTR17), .S(P2_P1_State2_PTR1), .Z(_03119__PTR1) );
  MUX2_X1 U24331 ( .A(1'b0), .B(_03118__PTR18), .S(P2_P1_State2_PTR1), .Z(_03119__PTR2) );
  MUX2_X1 U24332 ( .A(1'b0), .B(_03118__PTR19), .S(P2_P1_State2_PTR1), .Z(_03119__PTR3) );
  MUX2_X1 U24333 ( .A(1'b0), .B(_03118__PTR20), .S(P2_P1_State2_PTR1), .Z(_03119__PTR4) );
  MUX2_X1 U24334 ( .A(1'b0), .B(_03118__PTR21), .S(P2_P1_State2_PTR1), .Z(_03119__PTR5) );
  MUX2_X1 U24335 ( .A(1'b0), .B(_03118__PTR22), .S(P2_P1_State2_PTR1), .Z(_03119__PTR6) );
  MUX2_X1 U24336 ( .A(1'b0), .B(_03118__PTR23), .S(P2_P1_State2_PTR1), .Z(_03119__PTR7) );
  MUX2_X1 U24337 ( .A(_03118__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03119__PTR32) );
  MUX2_X1 U24338 ( .A(_03118__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03119__PTR33) );
  MUX2_X1 U24339 ( .A(_03118__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03119__PTR34) );
  MUX2_X1 U24340 ( .A(_03118__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03119__PTR35) );
  MUX2_X1 U24341 ( .A(_03118__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03119__PTR36) );
  MUX2_X1 U24342 ( .A(_03118__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03119__PTR37) );
  MUX2_X1 U24343 ( .A(_03118__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03119__PTR38) );
  MUX2_X1 U24344 ( .A(_03118__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03119__PTR39) );
  MUX2_X1 U24345 ( .A(_02196__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR16) );
  MUX2_X1 U24346 ( .A(_02196__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR17) );
  MUX2_X1 U24347 ( .A(_02196__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR18) );
  MUX2_X1 U24348 ( .A(_02196__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR19) );
  MUX2_X1 U24349 ( .A(_02196__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR20) );
  MUX2_X1 U24350 ( .A(_02196__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR21) );
  MUX2_X1 U24351 ( .A(_02196__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR22) );
  MUX2_X1 U24352 ( .A(_02196__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR23) );
  MUX2_X1 U24353 ( .A(_02196__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR32) );
  MUX2_X1 U24354 ( .A(_02196__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR33) );
  MUX2_X1 U24355 ( .A(_02196__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR34) );
  MUX2_X1 U24356 ( .A(_02196__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR35) );
  MUX2_X1 U24357 ( .A(_02196__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR36) );
  MUX2_X1 U24358 ( .A(_02196__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR37) );
  MUX2_X1 U24359 ( .A(_02196__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR38) );
  MUX2_X1 U24360 ( .A(_02196__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR39) );
  MUX2_X1 U24361 ( .A(_02196__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR64) );
  MUX2_X1 U24362 ( .A(_02196__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR65) );
  MUX2_X1 U24363 ( .A(_02196__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR66) );
  MUX2_X1 U24364 ( .A(_02196__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR67) );
  MUX2_X1 U24365 ( .A(_02196__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR68) );
  MUX2_X1 U24366 ( .A(_02196__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR69) );
  MUX2_X1 U24367 ( .A(_02196__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR70) );
  MUX2_X1 U24368 ( .A(_02196__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03118__PTR71) );
  MUX2_X1 U24369 ( .A(_03123__PTR0), .B(_03121__PTR64), .S(P2_P1_State2_PTR3), .Z(_02199__PTR0) );
  MUX2_X1 U24370 ( .A(_03123__PTR1), .B(_03121__PTR65), .S(P2_P1_State2_PTR3), .Z(_02199__PTR1) );
  MUX2_X1 U24371 ( .A(_03123__PTR2), .B(_03121__PTR66), .S(P2_P1_State2_PTR3), .Z(_02199__PTR2) );
  MUX2_X1 U24372 ( .A(_03123__PTR3), .B(_03121__PTR67), .S(P2_P1_State2_PTR3), .Z(_02199__PTR3) );
  MUX2_X1 U24373 ( .A(_03123__PTR4), .B(_03121__PTR68), .S(P2_P1_State2_PTR3), .Z(_02199__PTR4) );
  MUX2_X1 U24374 ( .A(_03123__PTR5), .B(_03121__PTR69), .S(P2_P1_State2_PTR3), .Z(_02199__PTR5) );
  MUX2_X1 U24375 ( .A(_03123__PTR6), .B(_03121__PTR70), .S(P2_P1_State2_PTR3), .Z(_02199__PTR6) );
  MUX2_X1 U24376 ( .A(_03123__PTR7), .B(_03121__PTR71), .S(P2_P1_State2_PTR3), .Z(_02199__PTR7) );
  MUX2_X1 U24377 ( .A(_03122__PTR0), .B(_03122__PTR32), .S(P2_P1_State2_PTR2), .Z(_03123__PTR0) );
  MUX2_X1 U24378 ( .A(_03122__PTR1), .B(_03122__PTR33), .S(P2_P1_State2_PTR2), .Z(_03123__PTR1) );
  MUX2_X1 U24379 ( .A(_03122__PTR2), .B(_03122__PTR34), .S(P2_P1_State2_PTR2), .Z(_03123__PTR2) );
  MUX2_X1 U24380 ( .A(_03122__PTR3), .B(_03122__PTR35), .S(P2_P1_State2_PTR2), .Z(_03123__PTR3) );
  MUX2_X1 U24381 ( .A(_03122__PTR4), .B(_03122__PTR36), .S(P2_P1_State2_PTR2), .Z(_03123__PTR4) );
  MUX2_X1 U24382 ( .A(_03122__PTR5), .B(_03122__PTR37), .S(P2_P1_State2_PTR2), .Z(_03123__PTR5) );
  MUX2_X1 U24383 ( .A(_03122__PTR6), .B(_03122__PTR38), .S(P2_P1_State2_PTR2), .Z(_03123__PTR6) );
  MUX2_X1 U24384 ( .A(_03122__PTR7), .B(_03122__PTR39), .S(P2_P1_State2_PTR2), .Z(_03123__PTR7) );
  MUX2_X1 U24385 ( .A(1'b0), .B(_03121__PTR16), .S(P2_P1_State2_PTR1), .Z(_03122__PTR0) );
  MUX2_X1 U24386 ( .A(1'b0), .B(_03121__PTR17), .S(P2_P1_State2_PTR1), .Z(_03122__PTR1) );
  MUX2_X1 U24387 ( .A(1'b0), .B(_03121__PTR18), .S(P2_P1_State2_PTR1), .Z(_03122__PTR2) );
  MUX2_X1 U24388 ( .A(1'b0), .B(_03121__PTR19), .S(P2_P1_State2_PTR1), .Z(_03122__PTR3) );
  MUX2_X1 U24389 ( .A(1'b0), .B(_03121__PTR20), .S(P2_P1_State2_PTR1), .Z(_03122__PTR4) );
  MUX2_X1 U24390 ( .A(1'b0), .B(_03121__PTR21), .S(P2_P1_State2_PTR1), .Z(_03122__PTR5) );
  MUX2_X1 U24391 ( .A(1'b0), .B(_03121__PTR22), .S(P2_P1_State2_PTR1), .Z(_03122__PTR6) );
  MUX2_X1 U24392 ( .A(1'b0), .B(_03121__PTR23), .S(P2_P1_State2_PTR1), .Z(_03122__PTR7) );
  MUX2_X1 U24393 ( .A(_03121__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03122__PTR32) );
  MUX2_X1 U24394 ( .A(_03121__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03122__PTR33) );
  MUX2_X1 U24395 ( .A(_03121__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03122__PTR34) );
  MUX2_X1 U24396 ( .A(_03121__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03122__PTR35) );
  MUX2_X1 U24397 ( .A(_03121__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03122__PTR36) );
  MUX2_X1 U24398 ( .A(_03121__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03122__PTR37) );
  MUX2_X1 U24399 ( .A(_03121__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03122__PTR38) );
  MUX2_X1 U24400 ( .A(_03121__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03122__PTR39) );
  MUX2_X1 U24401 ( .A(_02198__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR16) );
  MUX2_X1 U24402 ( .A(_02198__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR17) );
  MUX2_X1 U24403 ( .A(_02198__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR18) );
  MUX2_X1 U24404 ( .A(_02198__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR19) );
  MUX2_X1 U24405 ( .A(_02198__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR20) );
  MUX2_X1 U24406 ( .A(_02198__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR21) );
  MUX2_X1 U24407 ( .A(_02198__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR22) );
  MUX2_X1 U24408 ( .A(_02198__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR23) );
  MUX2_X1 U24409 ( .A(_02198__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR32) );
  MUX2_X1 U24410 ( .A(_02198__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR33) );
  MUX2_X1 U24411 ( .A(_02198__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR34) );
  MUX2_X1 U24412 ( .A(_02198__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR35) );
  MUX2_X1 U24413 ( .A(_02198__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR36) );
  MUX2_X1 U24414 ( .A(_02198__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR37) );
  MUX2_X1 U24415 ( .A(_02198__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR38) );
  MUX2_X1 U24416 ( .A(_02198__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR39) );
  MUX2_X1 U24417 ( .A(_02198__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR64) );
  MUX2_X1 U24418 ( .A(_02198__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR65) );
  MUX2_X1 U24419 ( .A(_02198__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR66) );
  MUX2_X1 U24420 ( .A(_02198__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR67) );
  MUX2_X1 U24421 ( .A(_02198__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR68) );
  MUX2_X1 U24422 ( .A(_02198__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR69) );
  MUX2_X1 U24423 ( .A(_02198__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR70) );
  MUX2_X1 U24424 ( .A(_02198__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03121__PTR71) );
  MUX2_X1 U24425 ( .A(_03126__PTR0), .B(_03124__PTR64), .S(P2_P1_State2_PTR3), .Z(_02201__PTR0) );
  MUX2_X1 U24426 ( .A(_03126__PTR1), .B(_03124__PTR65), .S(P2_P1_State2_PTR3), .Z(_02201__PTR1) );
  MUX2_X1 U24427 ( .A(_03126__PTR2), .B(_03124__PTR66), .S(P2_P1_State2_PTR3), .Z(_02201__PTR2) );
  MUX2_X1 U24428 ( .A(_03126__PTR3), .B(_03124__PTR67), .S(P2_P1_State2_PTR3), .Z(_02201__PTR3) );
  MUX2_X1 U24429 ( .A(_03126__PTR4), .B(_03124__PTR68), .S(P2_P1_State2_PTR3), .Z(_02201__PTR4) );
  MUX2_X1 U24430 ( .A(_03126__PTR5), .B(_03124__PTR69), .S(P2_P1_State2_PTR3), .Z(_02201__PTR5) );
  MUX2_X1 U24431 ( .A(_03126__PTR6), .B(_03124__PTR70), .S(P2_P1_State2_PTR3), .Z(_02201__PTR6) );
  MUX2_X1 U24432 ( .A(_03126__PTR7), .B(_03124__PTR71), .S(P2_P1_State2_PTR3), .Z(_02201__PTR7) );
  MUX2_X1 U24433 ( .A(_03125__PTR0), .B(_03125__PTR32), .S(P2_P1_State2_PTR2), .Z(_03126__PTR0) );
  MUX2_X1 U24434 ( .A(_03125__PTR1), .B(_03125__PTR33), .S(P2_P1_State2_PTR2), .Z(_03126__PTR1) );
  MUX2_X1 U24435 ( .A(_03125__PTR2), .B(_03125__PTR34), .S(P2_P1_State2_PTR2), .Z(_03126__PTR2) );
  MUX2_X1 U24436 ( .A(_03125__PTR3), .B(_03125__PTR35), .S(P2_P1_State2_PTR2), .Z(_03126__PTR3) );
  MUX2_X1 U24437 ( .A(_03125__PTR4), .B(_03125__PTR36), .S(P2_P1_State2_PTR2), .Z(_03126__PTR4) );
  MUX2_X1 U24438 ( .A(_03125__PTR5), .B(_03125__PTR37), .S(P2_P1_State2_PTR2), .Z(_03126__PTR5) );
  MUX2_X1 U24439 ( .A(_03125__PTR6), .B(_03125__PTR38), .S(P2_P1_State2_PTR2), .Z(_03126__PTR6) );
  MUX2_X1 U24440 ( .A(_03125__PTR7), .B(_03125__PTR39), .S(P2_P1_State2_PTR2), .Z(_03126__PTR7) );
  MUX2_X1 U24441 ( .A(1'b0), .B(_03124__PTR16), .S(P2_P1_State2_PTR1), .Z(_03125__PTR0) );
  MUX2_X1 U24442 ( .A(1'b0), .B(_03124__PTR17), .S(P2_P1_State2_PTR1), .Z(_03125__PTR1) );
  MUX2_X1 U24443 ( .A(1'b0), .B(_03124__PTR18), .S(P2_P1_State2_PTR1), .Z(_03125__PTR2) );
  MUX2_X1 U24444 ( .A(1'b0), .B(_03124__PTR19), .S(P2_P1_State2_PTR1), .Z(_03125__PTR3) );
  MUX2_X1 U24445 ( .A(1'b0), .B(_03124__PTR20), .S(P2_P1_State2_PTR1), .Z(_03125__PTR4) );
  MUX2_X1 U24446 ( .A(1'b0), .B(_03124__PTR21), .S(P2_P1_State2_PTR1), .Z(_03125__PTR5) );
  MUX2_X1 U24447 ( .A(1'b0), .B(_03124__PTR22), .S(P2_P1_State2_PTR1), .Z(_03125__PTR6) );
  MUX2_X1 U24448 ( .A(1'b0), .B(_03124__PTR23), .S(P2_P1_State2_PTR1), .Z(_03125__PTR7) );
  MUX2_X1 U24449 ( .A(_03124__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03125__PTR32) );
  MUX2_X1 U24450 ( .A(_03124__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03125__PTR33) );
  MUX2_X1 U24451 ( .A(_03124__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03125__PTR34) );
  MUX2_X1 U24452 ( .A(_03124__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03125__PTR35) );
  MUX2_X1 U24453 ( .A(_03124__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03125__PTR36) );
  MUX2_X1 U24454 ( .A(_03124__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03125__PTR37) );
  MUX2_X1 U24455 ( .A(_03124__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03125__PTR38) );
  MUX2_X1 U24456 ( .A(_03124__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03125__PTR39) );
  MUX2_X1 U24457 ( .A(_02200__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR16) );
  MUX2_X1 U24458 ( .A(_02200__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR17) );
  MUX2_X1 U24459 ( .A(_02200__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR18) );
  MUX2_X1 U24460 ( .A(_02200__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR19) );
  MUX2_X1 U24461 ( .A(_02200__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR20) );
  MUX2_X1 U24462 ( .A(_02200__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR21) );
  MUX2_X1 U24463 ( .A(_02200__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR22) );
  MUX2_X1 U24464 ( .A(_02200__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR23) );
  MUX2_X1 U24465 ( .A(_02200__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR32) );
  MUX2_X1 U24466 ( .A(_02200__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR33) );
  MUX2_X1 U24467 ( .A(_02200__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR34) );
  MUX2_X1 U24468 ( .A(_02200__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR35) );
  MUX2_X1 U24469 ( .A(_02200__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR36) );
  MUX2_X1 U24470 ( .A(_02200__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR37) );
  MUX2_X1 U24471 ( .A(_02200__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR38) );
  MUX2_X1 U24472 ( .A(_02200__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR39) );
  MUX2_X1 U24473 ( .A(_02200__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR64) );
  MUX2_X1 U24474 ( .A(_02200__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR65) );
  MUX2_X1 U24475 ( .A(_02200__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR66) );
  MUX2_X1 U24476 ( .A(_02200__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR67) );
  MUX2_X1 U24477 ( .A(_02200__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR68) );
  MUX2_X1 U24478 ( .A(_02200__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR69) );
  MUX2_X1 U24479 ( .A(_02200__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR70) );
  MUX2_X1 U24480 ( .A(_02200__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03124__PTR71) );
  MUX2_X1 U24481 ( .A(_03129__PTR0), .B(_03127__PTR64), .S(P2_P1_State2_PTR3), .Z(_02203__PTR0) );
  MUX2_X1 U24482 ( .A(_03129__PTR1), .B(_03127__PTR65), .S(P2_P1_State2_PTR3), .Z(_02203__PTR1) );
  MUX2_X1 U24483 ( .A(_03129__PTR2), .B(_03127__PTR66), .S(P2_P1_State2_PTR3), .Z(_02203__PTR2) );
  MUX2_X1 U24484 ( .A(_03129__PTR3), .B(_03127__PTR67), .S(P2_P1_State2_PTR3), .Z(_02203__PTR3) );
  MUX2_X1 U24485 ( .A(_03129__PTR4), .B(_03127__PTR68), .S(P2_P1_State2_PTR3), .Z(_02203__PTR4) );
  MUX2_X1 U24486 ( .A(_03129__PTR5), .B(_03127__PTR69), .S(P2_P1_State2_PTR3), .Z(_02203__PTR5) );
  MUX2_X1 U24487 ( .A(_03129__PTR6), .B(_03127__PTR70), .S(P2_P1_State2_PTR3), .Z(_02203__PTR6) );
  MUX2_X1 U24488 ( .A(_03129__PTR7), .B(_03127__PTR71), .S(P2_P1_State2_PTR3), .Z(_02203__PTR7) );
  MUX2_X1 U24489 ( .A(_03128__PTR0), .B(_03128__PTR32), .S(P2_P1_State2_PTR2), .Z(_03129__PTR0) );
  MUX2_X1 U24490 ( .A(_03128__PTR1), .B(_03128__PTR33), .S(P2_P1_State2_PTR2), .Z(_03129__PTR1) );
  MUX2_X1 U24491 ( .A(_03128__PTR2), .B(_03128__PTR34), .S(P2_P1_State2_PTR2), .Z(_03129__PTR2) );
  MUX2_X1 U24492 ( .A(_03128__PTR3), .B(_03128__PTR35), .S(P2_P1_State2_PTR2), .Z(_03129__PTR3) );
  MUX2_X1 U24493 ( .A(_03128__PTR4), .B(_03128__PTR36), .S(P2_P1_State2_PTR2), .Z(_03129__PTR4) );
  MUX2_X1 U24494 ( .A(_03128__PTR5), .B(_03128__PTR37), .S(P2_P1_State2_PTR2), .Z(_03129__PTR5) );
  MUX2_X1 U24495 ( .A(_03128__PTR6), .B(_03128__PTR38), .S(P2_P1_State2_PTR2), .Z(_03129__PTR6) );
  MUX2_X1 U24496 ( .A(_03128__PTR7), .B(_03128__PTR39), .S(P2_P1_State2_PTR2), .Z(_03129__PTR7) );
  MUX2_X1 U24497 ( .A(1'b0), .B(_03127__PTR16), .S(P2_P1_State2_PTR1), .Z(_03128__PTR0) );
  MUX2_X1 U24498 ( .A(1'b0), .B(_03127__PTR17), .S(P2_P1_State2_PTR1), .Z(_03128__PTR1) );
  MUX2_X1 U24499 ( .A(1'b0), .B(_03127__PTR18), .S(P2_P1_State2_PTR1), .Z(_03128__PTR2) );
  MUX2_X1 U24500 ( .A(1'b0), .B(_03127__PTR19), .S(P2_P1_State2_PTR1), .Z(_03128__PTR3) );
  MUX2_X1 U24501 ( .A(1'b0), .B(_03127__PTR20), .S(P2_P1_State2_PTR1), .Z(_03128__PTR4) );
  MUX2_X1 U24502 ( .A(1'b0), .B(_03127__PTR21), .S(P2_P1_State2_PTR1), .Z(_03128__PTR5) );
  MUX2_X1 U24503 ( .A(1'b0), .B(_03127__PTR22), .S(P2_P1_State2_PTR1), .Z(_03128__PTR6) );
  MUX2_X1 U24504 ( .A(1'b0), .B(_03127__PTR23), .S(P2_P1_State2_PTR1), .Z(_03128__PTR7) );
  MUX2_X1 U24505 ( .A(_03127__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03128__PTR32) );
  MUX2_X1 U24506 ( .A(_03127__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03128__PTR33) );
  MUX2_X1 U24507 ( .A(_03127__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03128__PTR34) );
  MUX2_X1 U24508 ( .A(_03127__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03128__PTR35) );
  MUX2_X1 U24509 ( .A(_03127__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03128__PTR36) );
  MUX2_X1 U24510 ( .A(_03127__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03128__PTR37) );
  MUX2_X1 U24511 ( .A(_03127__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03128__PTR38) );
  MUX2_X1 U24512 ( .A(_03127__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03128__PTR39) );
  MUX2_X1 U24513 ( .A(_02202__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR16) );
  MUX2_X1 U24514 ( .A(_02202__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR17) );
  MUX2_X1 U24515 ( .A(_02202__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR18) );
  MUX2_X1 U24516 ( .A(_02202__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR19) );
  MUX2_X1 U24517 ( .A(_02202__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR20) );
  MUX2_X1 U24518 ( .A(_02202__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR21) );
  MUX2_X1 U24519 ( .A(_02202__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR22) );
  MUX2_X1 U24520 ( .A(_02202__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR23) );
  MUX2_X1 U24521 ( .A(_02202__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR32) );
  MUX2_X1 U24522 ( .A(_02202__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR33) );
  MUX2_X1 U24523 ( .A(_02202__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR34) );
  MUX2_X1 U24524 ( .A(_02202__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR35) );
  MUX2_X1 U24525 ( .A(_02202__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR36) );
  MUX2_X1 U24526 ( .A(_02202__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR37) );
  MUX2_X1 U24527 ( .A(_02202__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR38) );
  MUX2_X1 U24528 ( .A(_02202__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR39) );
  MUX2_X1 U24529 ( .A(_02202__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR64) );
  MUX2_X1 U24530 ( .A(_02202__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR65) );
  MUX2_X1 U24531 ( .A(_02202__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR66) );
  MUX2_X1 U24532 ( .A(_02202__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR67) );
  MUX2_X1 U24533 ( .A(_02202__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR68) );
  MUX2_X1 U24534 ( .A(_02202__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR69) );
  MUX2_X1 U24535 ( .A(_02202__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR70) );
  MUX2_X1 U24536 ( .A(_02202__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03127__PTR71) );
  MUX2_X1 U24537 ( .A(_03132__PTR0), .B(_03130__PTR64), .S(P2_P1_State2_PTR3), .Z(_02205__PTR0) );
  MUX2_X1 U24538 ( .A(_03132__PTR1), .B(_03130__PTR65), .S(P2_P1_State2_PTR3), .Z(_02205__PTR1) );
  MUX2_X1 U24539 ( .A(_03132__PTR2), .B(_03130__PTR66), .S(P2_P1_State2_PTR3), .Z(_02205__PTR2) );
  MUX2_X1 U24540 ( .A(_03132__PTR3), .B(_03130__PTR67), .S(P2_P1_State2_PTR3), .Z(_02205__PTR3) );
  MUX2_X1 U24541 ( .A(_03132__PTR4), .B(_03130__PTR68), .S(P2_P1_State2_PTR3), .Z(_02205__PTR4) );
  MUX2_X1 U24542 ( .A(_03132__PTR5), .B(_03130__PTR69), .S(P2_P1_State2_PTR3), .Z(_02205__PTR5) );
  MUX2_X1 U24543 ( .A(_03132__PTR6), .B(_03130__PTR70), .S(P2_P1_State2_PTR3), .Z(_02205__PTR6) );
  MUX2_X1 U24544 ( .A(_03132__PTR7), .B(_03130__PTR71), .S(P2_P1_State2_PTR3), .Z(_02205__PTR7) );
  MUX2_X1 U24545 ( .A(_03131__PTR0), .B(_03131__PTR32), .S(P2_P1_State2_PTR2), .Z(_03132__PTR0) );
  MUX2_X1 U24546 ( .A(_03131__PTR1), .B(_03131__PTR33), .S(P2_P1_State2_PTR2), .Z(_03132__PTR1) );
  MUX2_X1 U24547 ( .A(_03131__PTR2), .B(_03131__PTR34), .S(P2_P1_State2_PTR2), .Z(_03132__PTR2) );
  MUX2_X1 U24548 ( .A(_03131__PTR3), .B(_03131__PTR35), .S(P2_P1_State2_PTR2), .Z(_03132__PTR3) );
  MUX2_X1 U24549 ( .A(_03131__PTR4), .B(_03131__PTR36), .S(P2_P1_State2_PTR2), .Z(_03132__PTR4) );
  MUX2_X1 U24550 ( .A(_03131__PTR5), .B(_03131__PTR37), .S(P2_P1_State2_PTR2), .Z(_03132__PTR5) );
  MUX2_X1 U24551 ( .A(_03131__PTR6), .B(_03131__PTR38), .S(P2_P1_State2_PTR2), .Z(_03132__PTR6) );
  MUX2_X1 U24552 ( .A(_03131__PTR7), .B(_03131__PTR39), .S(P2_P1_State2_PTR2), .Z(_03132__PTR7) );
  MUX2_X1 U24553 ( .A(1'b0), .B(_03130__PTR16), .S(P2_P1_State2_PTR1), .Z(_03131__PTR0) );
  MUX2_X1 U24554 ( .A(1'b0), .B(_03130__PTR17), .S(P2_P1_State2_PTR1), .Z(_03131__PTR1) );
  MUX2_X1 U24555 ( .A(1'b0), .B(_03130__PTR18), .S(P2_P1_State2_PTR1), .Z(_03131__PTR2) );
  MUX2_X1 U24556 ( .A(1'b0), .B(_03130__PTR19), .S(P2_P1_State2_PTR1), .Z(_03131__PTR3) );
  MUX2_X1 U24557 ( .A(1'b0), .B(_03130__PTR20), .S(P2_P1_State2_PTR1), .Z(_03131__PTR4) );
  MUX2_X1 U24558 ( .A(1'b0), .B(_03130__PTR21), .S(P2_P1_State2_PTR1), .Z(_03131__PTR5) );
  MUX2_X1 U24559 ( .A(1'b0), .B(_03130__PTR22), .S(P2_P1_State2_PTR1), .Z(_03131__PTR6) );
  MUX2_X1 U24560 ( .A(1'b0), .B(_03130__PTR23), .S(P2_P1_State2_PTR1), .Z(_03131__PTR7) );
  MUX2_X1 U24561 ( .A(_03130__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03131__PTR32) );
  MUX2_X1 U24562 ( .A(_03130__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03131__PTR33) );
  MUX2_X1 U24563 ( .A(_03130__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03131__PTR34) );
  MUX2_X1 U24564 ( .A(_03130__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03131__PTR35) );
  MUX2_X1 U24565 ( .A(_03130__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03131__PTR36) );
  MUX2_X1 U24566 ( .A(_03130__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03131__PTR37) );
  MUX2_X1 U24567 ( .A(_03130__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03131__PTR38) );
  MUX2_X1 U24568 ( .A(_03130__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03131__PTR39) );
  MUX2_X1 U24569 ( .A(_02204__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR16) );
  MUX2_X1 U24570 ( .A(_02204__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR17) );
  MUX2_X1 U24571 ( .A(_02204__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR18) );
  MUX2_X1 U24572 ( .A(_02204__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR19) );
  MUX2_X1 U24573 ( .A(_02204__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR20) );
  MUX2_X1 U24574 ( .A(_02204__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR21) );
  MUX2_X1 U24575 ( .A(_02204__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR22) );
  MUX2_X1 U24576 ( .A(_02204__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR23) );
  MUX2_X1 U24577 ( .A(_02204__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR32) );
  MUX2_X1 U24578 ( .A(_02204__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR33) );
  MUX2_X1 U24579 ( .A(_02204__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR34) );
  MUX2_X1 U24580 ( .A(_02204__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR35) );
  MUX2_X1 U24581 ( .A(_02204__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR36) );
  MUX2_X1 U24582 ( .A(_02204__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR37) );
  MUX2_X1 U24583 ( .A(_02204__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR38) );
  MUX2_X1 U24584 ( .A(_02204__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR39) );
  MUX2_X1 U24585 ( .A(_02204__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR64) );
  MUX2_X1 U24586 ( .A(_02204__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR65) );
  MUX2_X1 U24587 ( .A(_02204__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR66) );
  MUX2_X1 U24588 ( .A(_02204__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR67) );
  MUX2_X1 U24589 ( .A(_02204__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR68) );
  MUX2_X1 U24590 ( .A(_02204__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR69) );
  MUX2_X1 U24591 ( .A(_02204__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR70) );
  MUX2_X1 U24592 ( .A(_02204__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03130__PTR71) );
  MUX2_X1 U24593 ( .A(_03135__PTR0), .B(_03133__PTR64), .S(P2_P1_State2_PTR3), .Z(_02207__PTR0) );
  MUX2_X1 U24594 ( .A(_03135__PTR1), .B(_03133__PTR65), .S(P2_P1_State2_PTR3), .Z(_02207__PTR1) );
  MUX2_X1 U24595 ( .A(_03135__PTR2), .B(_03133__PTR66), .S(P2_P1_State2_PTR3), .Z(_02207__PTR2) );
  MUX2_X1 U24596 ( .A(_03135__PTR3), .B(_03133__PTR67), .S(P2_P1_State2_PTR3), .Z(_02207__PTR3) );
  MUX2_X1 U24597 ( .A(_03135__PTR4), .B(_03133__PTR68), .S(P2_P1_State2_PTR3), .Z(_02207__PTR4) );
  MUX2_X1 U24598 ( .A(_03135__PTR5), .B(_03133__PTR69), .S(P2_P1_State2_PTR3), .Z(_02207__PTR5) );
  MUX2_X1 U24599 ( .A(_03135__PTR6), .B(_03133__PTR70), .S(P2_P1_State2_PTR3), .Z(_02207__PTR6) );
  MUX2_X1 U24600 ( .A(_03135__PTR7), .B(_03133__PTR71), .S(P2_P1_State2_PTR3), .Z(_02207__PTR7) );
  MUX2_X1 U24601 ( .A(_03134__PTR0), .B(_03134__PTR32), .S(P2_P1_State2_PTR2), .Z(_03135__PTR0) );
  MUX2_X1 U24602 ( .A(_03134__PTR1), .B(_03134__PTR33), .S(P2_P1_State2_PTR2), .Z(_03135__PTR1) );
  MUX2_X1 U24603 ( .A(_03134__PTR2), .B(_03134__PTR34), .S(P2_P1_State2_PTR2), .Z(_03135__PTR2) );
  MUX2_X1 U24604 ( .A(_03134__PTR3), .B(_03134__PTR35), .S(P2_P1_State2_PTR2), .Z(_03135__PTR3) );
  MUX2_X1 U24605 ( .A(_03134__PTR4), .B(_03134__PTR36), .S(P2_P1_State2_PTR2), .Z(_03135__PTR4) );
  MUX2_X1 U24606 ( .A(_03134__PTR5), .B(_03134__PTR37), .S(P2_P1_State2_PTR2), .Z(_03135__PTR5) );
  MUX2_X1 U24607 ( .A(_03134__PTR6), .B(_03134__PTR38), .S(P2_P1_State2_PTR2), .Z(_03135__PTR6) );
  MUX2_X1 U24608 ( .A(_03134__PTR7), .B(_03134__PTR39), .S(P2_P1_State2_PTR2), .Z(_03135__PTR7) );
  MUX2_X1 U24609 ( .A(1'b0), .B(_03133__PTR16), .S(P2_P1_State2_PTR1), .Z(_03134__PTR0) );
  MUX2_X1 U24610 ( .A(1'b0), .B(_03133__PTR17), .S(P2_P1_State2_PTR1), .Z(_03134__PTR1) );
  MUX2_X1 U24611 ( .A(1'b0), .B(_03133__PTR18), .S(P2_P1_State2_PTR1), .Z(_03134__PTR2) );
  MUX2_X1 U24612 ( .A(1'b0), .B(_03133__PTR19), .S(P2_P1_State2_PTR1), .Z(_03134__PTR3) );
  MUX2_X1 U24613 ( .A(1'b0), .B(_03133__PTR20), .S(P2_P1_State2_PTR1), .Z(_03134__PTR4) );
  MUX2_X1 U24614 ( .A(1'b0), .B(_03133__PTR21), .S(P2_P1_State2_PTR1), .Z(_03134__PTR5) );
  MUX2_X1 U24615 ( .A(1'b0), .B(_03133__PTR22), .S(P2_P1_State2_PTR1), .Z(_03134__PTR6) );
  MUX2_X1 U24616 ( .A(1'b0), .B(_03133__PTR23), .S(P2_P1_State2_PTR1), .Z(_03134__PTR7) );
  MUX2_X1 U24617 ( .A(_03133__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03134__PTR32) );
  MUX2_X1 U24618 ( .A(_03133__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03134__PTR33) );
  MUX2_X1 U24619 ( .A(_03133__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03134__PTR34) );
  MUX2_X1 U24620 ( .A(_03133__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03134__PTR35) );
  MUX2_X1 U24621 ( .A(_03133__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03134__PTR36) );
  MUX2_X1 U24622 ( .A(_03133__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03134__PTR37) );
  MUX2_X1 U24623 ( .A(_03133__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03134__PTR38) );
  MUX2_X1 U24624 ( .A(_03133__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03134__PTR39) );
  MUX2_X1 U24625 ( .A(_02206__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR16) );
  MUX2_X1 U24626 ( .A(_02206__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR17) );
  MUX2_X1 U24627 ( .A(_02206__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR18) );
  MUX2_X1 U24628 ( .A(_02206__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR19) );
  MUX2_X1 U24629 ( .A(_02206__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR20) );
  MUX2_X1 U24630 ( .A(_02206__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR21) );
  MUX2_X1 U24631 ( .A(_02206__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR22) );
  MUX2_X1 U24632 ( .A(_02206__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR23) );
  MUX2_X1 U24633 ( .A(_02206__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR32) );
  MUX2_X1 U24634 ( .A(_02206__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR33) );
  MUX2_X1 U24635 ( .A(_02206__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR34) );
  MUX2_X1 U24636 ( .A(_02206__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR35) );
  MUX2_X1 U24637 ( .A(_02206__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR36) );
  MUX2_X1 U24638 ( .A(_02206__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR37) );
  MUX2_X1 U24639 ( .A(_02206__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR38) );
  MUX2_X1 U24640 ( .A(_02206__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR39) );
  MUX2_X1 U24641 ( .A(_02206__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR64) );
  MUX2_X1 U24642 ( .A(_02206__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR65) );
  MUX2_X1 U24643 ( .A(_02206__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR66) );
  MUX2_X1 U24644 ( .A(_02206__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR67) );
  MUX2_X1 U24645 ( .A(_02206__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR68) );
  MUX2_X1 U24646 ( .A(_02206__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR69) );
  MUX2_X1 U24647 ( .A(_02206__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR70) );
  MUX2_X1 U24648 ( .A(_02206__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03133__PTR71) );
  MUX2_X1 U24649 ( .A(_03138__PTR0), .B(_03136__PTR64), .S(P2_P1_State2_PTR3), .Z(_02209__PTR0) );
  MUX2_X1 U24650 ( .A(_03138__PTR1), .B(_03136__PTR65), .S(P2_P1_State2_PTR3), .Z(_02209__PTR1) );
  MUX2_X1 U24651 ( .A(_03138__PTR2), .B(_03136__PTR66), .S(P2_P1_State2_PTR3), .Z(_02209__PTR2) );
  MUX2_X1 U24652 ( .A(_03138__PTR3), .B(_03136__PTR67), .S(P2_P1_State2_PTR3), .Z(_02209__PTR3) );
  MUX2_X1 U24653 ( .A(_03138__PTR4), .B(_03136__PTR68), .S(P2_P1_State2_PTR3), .Z(_02209__PTR4) );
  MUX2_X1 U24654 ( .A(_03138__PTR5), .B(_03136__PTR69), .S(P2_P1_State2_PTR3), .Z(_02209__PTR5) );
  MUX2_X1 U24655 ( .A(_03138__PTR6), .B(_03136__PTR70), .S(P2_P1_State2_PTR3), .Z(_02209__PTR6) );
  MUX2_X1 U24656 ( .A(_03138__PTR7), .B(_03136__PTR71), .S(P2_P1_State2_PTR3), .Z(_02209__PTR7) );
  MUX2_X1 U24657 ( .A(_03137__PTR0), .B(_03137__PTR32), .S(P2_P1_State2_PTR2), .Z(_03138__PTR0) );
  MUX2_X1 U24658 ( .A(_03137__PTR1), .B(_03137__PTR33), .S(P2_P1_State2_PTR2), .Z(_03138__PTR1) );
  MUX2_X1 U24659 ( .A(_03137__PTR2), .B(_03137__PTR34), .S(P2_P1_State2_PTR2), .Z(_03138__PTR2) );
  MUX2_X1 U24660 ( .A(_03137__PTR3), .B(_03137__PTR35), .S(P2_P1_State2_PTR2), .Z(_03138__PTR3) );
  MUX2_X1 U24661 ( .A(_03137__PTR4), .B(_03137__PTR36), .S(P2_P1_State2_PTR2), .Z(_03138__PTR4) );
  MUX2_X1 U24662 ( .A(_03137__PTR5), .B(_03137__PTR37), .S(P2_P1_State2_PTR2), .Z(_03138__PTR5) );
  MUX2_X1 U24663 ( .A(_03137__PTR6), .B(_03137__PTR38), .S(P2_P1_State2_PTR2), .Z(_03138__PTR6) );
  MUX2_X1 U24664 ( .A(_03137__PTR7), .B(_03137__PTR39), .S(P2_P1_State2_PTR2), .Z(_03138__PTR7) );
  MUX2_X1 U24665 ( .A(1'b0), .B(_03136__PTR16), .S(P2_P1_State2_PTR1), .Z(_03137__PTR0) );
  MUX2_X1 U24666 ( .A(1'b0), .B(_03136__PTR17), .S(P2_P1_State2_PTR1), .Z(_03137__PTR1) );
  MUX2_X1 U24667 ( .A(1'b0), .B(_03136__PTR18), .S(P2_P1_State2_PTR1), .Z(_03137__PTR2) );
  MUX2_X1 U24668 ( .A(1'b0), .B(_03136__PTR19), .S(P2_P1_State2_PTR1), .Z(_03137__PTR3) );
  MUX2_X1 U24669 ( .A(1'b0), .B(_03136__PTR20), .S(P2_P1_State2_PTR1), .Z(_03137__PTR4) );
  MUX2_X1 U24670 ( .A(1'b0), .B(_03136__PTR21), .S(P2_P1_State2_PTR1), .Z(_03137__PTR5) );
  MUX2_X1 U24671 ( .A(1'b0), .B(_03136__PTR22), .S(P2_P1_State2_PTR1), .Z(_03137__PTR6) );
  MUX2_X1 U24672 ( .A(1'b0), .B(_03136__PTR23), .S(P2_P1_State2_PTR1), .Z(_03137__PTR7) );
  MUX2_X1 U24673 ( .A(_03136__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03137__PTR32) );
  MUX2_X1 U24674 ( .A(_03136__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03137__PTR33) );
  MUX2_X1 U24675 ( .A(_03136__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03137__PTR34) );
  MUX2_X1 U24676 ( .A(_03136__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03137__PTR35) );
  MUX2_X1 U24677 ( .A(_03136__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03137__PTR36) );
  MUX2_X1 U24678 ( .A(_03136__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03137__PTR37) );
  MUX2_X1 U24679 ( .A(_03136__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03137__PTR38) );
  MUX2_X1 U24680 ( .A(_03136__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03137__PTR39) );
  MUX2_X1 U24681 ( .A(_02208__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR16) );
  MUX2_X1 U24682 ( .A(_02208__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR17) );
  MUX2_X1 U24683 ( .A(_02208__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR18) );
  MUX2_X1 U24684 ( .A(_02208__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR19) );
  MUX2_X1 U24685 ( .A(_02208__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR20) );
  MUX2_X1 U24686 ( .A(_02208__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR21) );
  MUX2_X1 U24687 ( .A(_02208__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR22) );
  MUX2_X1 U24688 ( .A(_02208__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR23) );
  MUX2_X1 U24689 ( .A(_02208__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR32) );
  MUX2_X1 U24690 ( .A(_02208__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR33) );
  MUX2_X1 U24691 ( .A(_02208__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR34) );
  MUX2_X1 U24692 ( .A(_02208__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR35) );
  MUX2_X1 U24693 ( .A(_02208__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR36) );
  MUX2_X1 U24694 ( .A(_02208__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR37) );
  MUX2_X1 U24695 ( .A(_02208__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR38) );
  MUX2_X1 U24696 ( .A(_02208__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR39) );
  MUX2_X1 U24697 ( .A(_02208__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR64) );
  MUX2_X1 U24698 ( .A(_02208__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR65) );
  MUX2_X1 U24699 ( .A(_02208__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR66) );
  MUX2_X1 U24700 ( .A(_02208__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR67) );
  MUX2_X1 U24701 ( .A(_02208__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR68) );
  MUX2_X1 U24702 ( .A(_02208__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR69) );
  MUX2_X1 U24703 ( .A(_02208__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR70) );
  MUX2_X1 U24704 ( .A(_02208__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03136__PTR71) );
  MUX2_X1 U24705 ( .A(_03141__PTR0), .B(_03139__PTR64), .S(P2_P1_State2_PTR3), .Z(_02211__PTR0) );
  MUX2_X1 U24706 ( .A(_03141__PTR1), .B(_03139__PTR65), .S(P2_P1_State2_PTR3), .Z(_02211__PTR1) );
  MUX2_X1 U24707 ( .A(_03141__PTR2), .B(_03139__PTR66), .S(P2_P1_State2_PTR3), .Z(_02211__PTR2) );
  MUX2_X1 U24708 ( .A(_03141__PTR3), .B(_03139__PTR67), .S(P2_P1_State2_PTR3), .Z(_02211__PTR3) );
  MUX2_X1 U24709 ( .A(_03141__PTR4), .B(_03139__PTR68), .S(P2_P1_State2_PTR3), .Z(_02211__PTR4) );
  MUX2_X1 U24710 ( .A(_03141__PTR5), .B(_03139__PTR69), .S(P2_P1_State2_PTR3), .Z(_02211__PTR5) );
  MUX2_X1 U24711 ( .A(_03141__PTR6), .B(_03139__PTR70), .S(P2_P1_State2_PTR3), .Z(_02211__PTR6) );
  MUX2_X1 U24712 ( .A(_03141__PTR7), .B(_03139__PTR71), .S(P2_P1_State2_PTR3), .Z(_02211__PTR7) );
  MUX2_X1 U24713 ( .A(_03140__PTR0), .B(_03140__PTR32), .S(P2_P1_State2_PTR2), .Z(_03141__PTR0) );
  MUX2_X1 U24714 ( .A(_03140__PTR1), .B(_03140__PTR33), .S(P2_P1_State2_PTR2), .Z(_03141__PTR1) );
  MUX2_X1 U24715 ( .A(_03140__PTR2), .B(_03140__PTR34), .S(P2_P1_State2_PTR2), .Z(_03141__PTR2) );
  MUX2_X1 U24716 ( .A(_03140__PTR3), .B(_03140__PTR35), .S(P2_P1_State2_PTR2), .Z(_03141__PTR3) );
  MUX2_X1 U24717 ( .A(_03140__PTR4), .B(_03140__PTR36), .S(P2_P1_State2_PTR2), .Z(_03141__PTR4) );
  MUX2_X1 U24718 ( .A(_03140__PTR5), .B(_03140__PTR37), .S(P2_P1_State2_PTR2), .Z(_03141__PTR5) );
  MUX2_X1 U24719 ( .A(_03140__PTR6), .B(_03140__PTR38), .S(P2_P1_State2_PTR2), .Z(_03141__PTR6) );
  MUX2_X1 U24720 ( .A(_03140__PTR7), .B(_03140__PTR39), .S(P2_P1_State2_PTR2), .Z(_03141__PTR7) );
  MUX2_X1 U24721 ( .A(1'b0), .B(_03139__PTR16), .S(P2_P1_State2_PTR1), .Z(_03140__PTR0) );
  MUX2_X1 U24722 ( .A(1'b0), .B(_03139__PTR17), .S(P2_P1_State2_PTR1), .Z(_03140__PTR1) );
  MUX2_X1 U24723 ( .A(1'b0), .B(_03139__PTR18), .S(P2_P1_State2_PTR1), .Z(_03140__PTR2) );
  MUX2_X1 U24724 ( .A(1'b0), .B(_03139__PTR19), .S(P2_P1_State2_PTR1), .Z(_03140__PTR3) );
  MUX2_X1 U24725 ( .A(1'b0), .B(_03139__PTR20), .S(P2_P1_State2_PTR1), .Z(_03140__PTR4) );
  MUX2_X1 U24726 ( .A(1'b0), .B(_03139__PTR21), .S(P2_P1_State2_PTR1), .Z(_03140__PTR5) );
  MUX2_X1 U24727 ( .A(1'b0), .B(_03139__PTR22), .S(P2_P1_State2_PTR1), .Z(_03140__PTR6) );
  MUX2_X1 U24728 ( .A(1'b0), .B(_03139__PTR23), .S(P2_P1_State2_PTR1), .Z(_03140__PTR7) );
  MUX2_X1 U24729 ( .A(_03139__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03140__PTR32) );
  MUX2_X1 U24730 ( .A(_03139__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03140__PTR33) );
  MUX2_X1 U24731 ( .A(_03139__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03140__PTR34) );
  MUX2_X1 U24732 ( .A(_03139__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03140__PTR35) );
  MUX2_X1 U24733 ( .A(_03139__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03140__PTR36) );
  MUX2_X1 U24734 ( .A(_03139__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03140__PTR37) );
  MUX2_X1 U24735 ( .A(_03139__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03140__PTR38) );
  MUX2_X1 U24736 ( .A(_03139__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03140__PTR39) );
  MUX2_X1 U24737 ( .A(_02210__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR16) );
  MUX2_X1 U24738 ( .A(_02210__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR17) );
  MUX2_X1 U24739 ( .A(_02210__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR18) );
  MUX2_X1 U24740 ( .A(_02210__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR19) );
  MUX2_X1 U24741 ( .A(_02210__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR20) );
  MUX2_X1 U24742 ( .A(_02210__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR21) );
  MUX2_X1 U24743 ( .A(_02210__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR22) );
  MUX2_X1 U24744 ( .A(_02210__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR23) );
  MUX2_X1 U24745 ( .A(_02210__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR32) );
  MUX2_X1 U24746 ( .A(_02210__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR33) );
  MUX2_X1 U24747 ( .A(_02210__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR34) );
  MUX2_X1 U24748 ( .A(_02210__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR35) );
  MUX2_X1 U24749 ( .A(_02210__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR36) );
  MUX2_X1 U24750 ( .A(_02210__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR37) );
  MUX2_X1 U24751 ( .A(_02210__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR38) );
  MUX2_X1 U24752 ( .A(_02210__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR39) );
  MUX2_X1 U24753 ( .A(_02210__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR64) );
  MUX2_X1 U24754 ( .A(_02210__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR65) );
  MUX2_X1 U24755 ( .A(_02210__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR66) );
  MUX2_X1 U24756 ( .A(_02210__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR67) );
  MUX2_X1 U24757 ( .A(_02210__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR68) );
  MUX2_X1 U24758 ( .A(_02210__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR69) );
  MUX2_X1 U24759 ( .A(_02210__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR70) );
  MUX2_X1 U24760 ( .A(_02210__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03139__PTR71) );
  MUX2_X1 U24761 ( .A(_03144__PTR0), .B(_03142__PTR64), .S(P2_P1_State2_PTR3), .Z(_02213__PTR0) );
  MUX2_X1 U24762 ( .A(_03144__PTR1), .B(_03142__PTR65), .S(P2_P1_State2_PTR3), .Z(_02213__PTR1) );
  MUX2_X1 U24763 ( .A(_03144__PTR2), .B(_03142__PTR66), .S(P2_P1_State2_PTR3), .Z(_02213__PTR2) );
  MUX2_X1 U24764 ( .A(_03144__PTR3), .B(_03142__PTR67), .S(P2_P1_State2_PTR3), .Z(_02213__PTR3) );
  MUX2_X1 U24765 ( .A(_03144__PTR4), .B(_03142__PTR68), .S(P2_P1_State2_PTR3), .Z(_02213__PTR4) );
  MUX2_X1 U24766 ( .A(_03144__PTR5), .B(_03142__PTR69), .S(P2_P1_State2_PTR3), .Z(_02213__PTR5) );
  MUX2_X1 U24767 ( .A(_03144__PTR6), .B(_03142__PTR70), .S(P2_P1_State2_PTR3), .Z(_02213__PTR6) );
  MUX2_X1 U24768 ( .A(_03144__PTR7), .B(_03142__PTR71), .S(P2_P1_State2_PTR3), .Z(_02213__PTR7) );
  MUX2_X1 U24769 ( .A(_03143__PTR0), .B(_03143__PTR32), .S(P2_P1_State2_PTR2), .Z(_03144__PTR0) );
  MUX2_X1 U24770 ( .A(_03143__PTR1), .B(_03143__PTR33), .S(P2_P1_State2_PTR2), .Z(_03144__PTR1) );
  MUX2_X1 U24771 ( .A(_03143__PTR2), .B(_03143__PTR34), .S(P2_P1_State2_PTR2), .Z(_03144__PTR2) );
  MUX2_X1 U24772 ( .A(_03143__PTR3), .B(_03143__PTR35), .S(P2_P1_State2_PTR2), .Z(_03144__PTR3) );
  MUX2_X1 U24773 ( .A(_03143__PTR4), .B(_03143__PTR36), .S(P2_P1_State2_PTR2), .Z(_03144__PTR4) );
  MUX2_X1 U24774 ( .A(_03143__PTR5), .B(_03143__PTR37), .S(P2_P1_State2_PTR2), .Z(_03144__PTR5) );
  MUX2_X1 U24775 ( .A(_03143__PTR6), .B(_03143__PTR38), .S(P2_P1_State2_PTR2), .Z(_03144__PTR6) );
  MUX2_X1 U24776 ( .A(_03143__PTR7), .B(_03143__PTR39), .S(P2_P1_State2_PTR2), .Z(_03144__PTR7) );
  MUX2_X1 U24777 ( .A(1'b0), .B(_03142__PTR16), .S(P2_P1_State2_PTR1), .Z(_03143__PTR0) );
  MUX2_X1 U24778 ( .A(1'b0), .B(_03142__PTR17), .S(P2_P1_State2_PTR1), .Z(_03143__PTR1) );
  MUX2_X1 U24779 ( .A(1'b0), .B(_03142__PTR18), .S(P2_P1_State2_PTR1), .Z(_03143__PTR2) );
  MUX2_X1 U24780 ( .A(1'b0), .B(_03142__PTR19), .S(P2_P1_State2_PTR1), .Z(_03143__PTR3) );
  MUX2_X1 U24781 ( .A(1'b0), .B(_03142__PTR20), .S(P2_P1_State2_PTR1), .Z(_03143__PTR4) );
  MUX2_X1 U24782 ( .A(1'b0), .B(_03142__PTR21), .S(P2_P1_State2_PTR1), .Z(_03143__PTR5) );
  MUX2_X1 U24783 ( .A(1'b0), .B(_03142__PTR22), .S(P2_P1_State2_PTR1), .Z(_03143__PTR6) );
  MUX2_X1 U24784 ( .A(1'b0), .B(_03142__PTR23), .S(P2_P1_State2_PTR1), .Z(_03143__PTR7) );
  MUX2_X1 U24785 ( .A(_03142__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03143__PTR32) );
  MUX2_X1 U24786 ( .A(_03142__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03143__PTR33) );
  MUX2_X1 U24787 ( .A(_03142__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03143__PTR34) );
  MUX2_X1 U24788 ( .A(_03142__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03143__PTR35) );
  MUX2_X1 U24789 ( .A(_03142__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03143__PTR36) );
  MUX2_X1 U24790 ( .A(_03142__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03143__PTR37) );
  MUX2_X1 U24791 ( .A(_03142__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03143__PTR38) );
  MUX2_X1 U24792 ( .A(_03142__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03143__PTR39) );
  MUX2_X1 U24793 ( .A(_02212__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR16) );
  MUX2_X1 U24794 ( .A(_02212__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR17) );
  MUX2_X1 U24795 ( .A(_02212__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR18) );
  MUX2_X1 U24796 ( .A(_02212__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR19) );
  MUX2_X1 U24797 ( .A(_02212__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR20) );
  MUX2_X1 U24798 ( .A(_02212__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR21) );
  MUX2_X1 U24799 ( .A(_02212__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR22) );
  MUX2_X1 U24800 ( .A(_02212__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR23) );
  MUX2_X1 U24801 ( .A(_02212__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR32) );
  MUX2_X1 U24802 ( .A(_02212__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR33) );
  MUX2_X1 U24803 ( .A(_02212__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR34) );
  MUX2_X1 U24804 ( .A(_02212__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR35) );
  MUX2_X1 U24805 ( .A(_02212__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR36) );
  MUX2_X1 U24806 ( .A(_02212__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR37) );
  MUX2_X1 U24807 ( .A(_02212__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR38) );
  MUX2_X1 U24808 ( .A(_02212__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR39) );
  MUX2_X1 U24809 ( .A(_02212__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR64) );
  MUX2_X1 U24810 ( .A(_02212__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR65) );
  MUX2_X1 U24811 ( .A(_02212__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR66) );
  MUX2_X1 U24812 ( .A(_02212__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR67) );
  MUX2_X1 U24813 ( .A(_02212__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR68) );
  MUX2_X1 U24814 ( .A(_02212__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR69) );
  MUX2_X1 U24815 ( .A(_02212__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR70) );
  MUX2_X1 U24816 ( .A(_02212__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03142__PTR71) );
  MUX2_X1 U24817 ( .A(_03147__PTR0), .B(_03145__PTR64), .S(P2_P1_State2_PTR3), .Z(_02215__PTR0) );
  MUX2_X1 U24818 ( .A(_03147__PTR1), .B(_03145__PTR65), .S(P2_P1_State2_PTR3), .Z(_02215__PTR1) );
  MUX2_X1 U24819 ( .A(_03147__PTR2), .B(_03145__PTR66), .S(P2_P1_State2_PTR3), .Z(_02215__PTR2) );
  MUX2_X1 U24820 ( .A(_03147__PTR3), .B(_03145__PTR67), .S(P2_P1_State2_PTR3), .Z(_02215__PTR3) );
  MUX2_X1 U24821 ( .A(_03147__PTR4), .B(_03145__PTR68), .S(P2_P1_State2_PTR3), .Z(_02215__PTR4) );
  MUX2_X1 U24822 ( .A(_03147__PTR5), .B(_03145__PTR69), .S(P2_P1_State2_PTR3), .Z(_02215__PTR5) );
  MUX2_X1 U24823 ( .A(_03147__PTR6), .B(_03145__PTR70), .S(P2_P1_State2_PTR3), .Z(_02215__PTR6) );
  MUX2_X1 U24824 ( .A(_03147__PTR7), .B(_03145__PTR71), .S(P2_P1_State2_PTR3), .Z(_02215__PTR7) );
  MUX2_X1 U24825 ( .A(_03146__PTR0), .B(_03146__PTR32), .S(P2_P1_State2_PTR2), .Z(_03147__PTR0) );
  MUX2_X1 U24826 ( .A(_03146__PTR1), .B(_03146__PTR33), .S(P2_P1_State2_PTR2), .Z(_03147__PTR1) );
  MUX2_X1 U24827 ( .A(_03146__PTR2), .B(_03146__PTR34), .S(P2_P1_State2_PTR2), .Z(_03147__PTR2) );
  MUX2_X1 U24828 ( .A(_03146__PTR3), .B(_03146__PTR35), .S(P2_P1_State2_PTR2), .Z(_03147__PTR3) );
  MUX2_X1 U24829 ( .A(_03146__PTR4), .B(_03146__PTR36), .S(P2_P1_State2_PTR2), .Z(_03147__PTR4) );
  MUX2_X1 U24830 ( .A(_03146__PTR5), .B(_03146__PTR37), .S(P2_P1_State2_PTR2), .Z(_03147__PTR5) );
  MUX2_X1 U24831 ( .A(_03146__PTR6), .B(_03146__PTR38), .S(P2_P1_State2_PTR2), .Z(_03147__PTR6) );
  MUX2_X1 U24832 ( .A(_03146__PTR7), .B(_03146__PTR39), .S(P2_P1_State2_PTR2), .Z(_03147__PTR7) );
  MUX2_X1 U24833 ( .A(1'b0), .B(_03145__PTR16), .S(P2_P1_State2_PTR1), .Z(_03146__PTR0) );
  MUX2_X1 U24834 ( .A(1'b0), .B(_03145__PTR17), .S(P2_P1_State2_PTR1), .Z(_03146__PTR1) );
  MUX2_X1 U24835 ( .A(1'b0), .B(_03145__PTR18), .S(P2_P1_State2_PTR1), .Z(_03146__PTR2) );
  MUX2_X1 U24836 ( .A(1'b0), .B(_03145__PTR19), .S(P2_P1_State2_PTR1), .Z(_03146__PTR3) );
  MUX2_X1 U24837 ( .A(1'b0), .B(_03145__PTR20), .S(P2_P1_State2_PTR1), .Z(_03146__PTR4) );
  MUX2_X1 U24838 ( .A(1'b0), .B(_03145__PTR21), .S(P2_P1_State2_PTR1), .Z(_03146__PTR5) );
  MUX2_X1 U24839 ( .A(1'b0), .B(_03145__PTR22), .S(P2_P1_State2_PTR1), .Z(_03146__PTR6) );
  MUX2_X1 U24840 ( .A(1'b0), .B(_03145__PTR23), .S(P2_P1_State2_PTR1), .Z(_03146__PTR7) );
  MUX2_X1 U24841 ( .A(_03145__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03146__PTR32) );
  MUX2_X1 U24842 ( .A(_03145__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03146__PTR33) );
  MUX2_X1 U24843 ( .A(_03145__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03146__PTR34) );
  MUX2_X1 U24844 ( .A(_03145__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03146__PTR35) );
  MUX2_X1 U24845 ( .A(_03145__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03146__PTR36) );
  MUX2_X1 U24846 ( .A(_03145__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03146__PTR37) );
  MUX2_X1 U24847 ( .A(_03145__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03146__PTR38) );
  MUX2_X1 U24848 ( .A(_03145__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03146__PTR39) );
  MUX2_X1 U24849 ( .A(_02214__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR16) );
  MUX2_X1 U24850 ( .A(_02214__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR17) );
  MUX2_X1 U24851 ( .A(_02214__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR18) );
  MUX2_X1 U24852 ( .A(_02214__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR19) );
  MUX2_X1 U24853 ( .A(_02214__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR20) );
  MUX2_X1 U24854 ( .A(_02214__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR21) );
  MUX2_X1 U24855 ( .A(_02214__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR22) );
  MUX2_X1 U24856 ( .A(_02214__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR23) );
  MUX2_X1 U24857 ( .A(_02214__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR32) );
  MUX2_X1 U24858 ( .A(_02214__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR33) );
  MUX2_X1 U24859 ( .A(_02214__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR34) );
  MUX2_X1 U24860 ( .A(_02214__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR35) );
  MUX2_X1 U24861 ( .A(_02214__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR36) );
  MUX2_X1 U24862 ( .A(_02214__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR37) );
  MUX2_X1 U24863 ( .A(_02214__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR38) );
  MUX2_X1 U24864 ( .A(_02214__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR39) );
  MUX2_X1 U24865 ( .A(_02214__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR64) );
  MUX2_X1 U24866 ( .A(_02214__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR65) );
  MUX2_X1 U24867 ( .A(_02214__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR66) );
  MUX2_X1 U24868 ( .A(_02214__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR67) );
  MUX2_X1 U24869 ( .A(_02214__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR68) );
  MUX2_X1 U24870 ( .A(_02214__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR69) );
  MUX2_X1 U24871 ( .A(_02214__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR70) );
  MUX2_X1 U24872 ( .A(_02214__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03145__PTR71) );
  MUX2_X1 U24873 ( .A(_03150__PTR0), .B(_03148__PTR64), .S(P2_P1_State2_PTR3), .Z(_02217__PTR0) );
  MUX2_X1 U24874 ( .A(_03150__PTR1), .B(_03148__PTR65), .S(P2_P1_State2_PTR3), .Z(_02217__PTR1) );
  MUX2_X1 U24875 ( .A(_03150__PTR2), .B(_03148__PTR66), .S(P2_P1_State2_PTR3), .Z(_02217__PTR2) );
  MUX2_X1 U24876 ( .A(_03150__PTR3), .B(_03148__PTR67), .S(P2_P1_State2_PTR3), .Z(_02217__PTR3) );
  MUX2_X1 U24877 ( .A(_03150__PTR4), .B(_03148__PTR68), .S(P2_P1_State2_PTR3), .Z(_02217__PTR4) );
  MUX2_X1 U24878 ( .A(_03150__PTR5), .B(_03148__PTR69), .S(P2_P1_State2_PTR3), .Z(_02217__PTR5) );
  MUX2_X1 U24879 ( .A(_03150__PTR6), .B(_03148__PTR70), .S(P2_P1_State2_PTR3), .Z(_02217__PTR6) );
  MUX2_X1 U24880 ( .A(_03150__PTR7), .B(_03148__PTR71), .S(P2_P1_State2_PTR3), .Z(_02217__PTR7) );
  MUX2_X1 U24881 ( .A(_03149__PTR0), .B(_03149__PTR32), .S(P2_P1_State2_PTR2), .Z(_03150__PTR0) );
  MUX2_X1 U24882 ( .A(_03149__PTR1), .B(_03149__PTR33), .S(P2_P1_State2_PTR2), .Z(_03150__PTR1) );
  MUX2_X1 U24883 ( .A(_03149__PTR2), .B(_03149__PTR34), .S(P2_P1_State2_PTR2), .Z(_03150__PTR2) );
  MUX2_X1 U24884 ( .A(_03149__PTR3), .B(_03149__PTR35), .S(P2_P1_State2_PTR2), .Z(_03150__PTR3) );
  MUX2_X1 U24885 ( .A(_03149__PTR4), .B(_03149__PTR36), .S(P2_P1_State2_PTR2), .Z(_03150__PTR4) );
  MUX2_X1 U24886 ( .A(_03149__PTR5), .B(_03149__PTR37), .S(P2_P1_State2_PTR2), .Z(_03150__PTR5) );
  MUX2_X1 U24887 ( .A(_03149__PTR6), .B(_03149__PTR38), .S(P2_P1_State2_PTR2), .Z(_03150__PTR6) );
  MUX2_X1 U24888 ( .A(_03149__PTR7), .B(_03149__PTR39), .S(P2_P1_State2_PTR2), .Z(_03150__PTR7) );
  MUX2_X1 U24889 ( .A(1'b0), .B(_03148__PTR16), .S(P2_P1_State2_PTR1), .Z(_03149__PTR0) );
  MUX2_X1 U24890 ( .A(1'b0), .B(_03148__PTR17), .S(P2_P1_State2_PTR1), .Z(_03149__PTR1) );
  MUX2_X1 U24891 ( .A(1'b0), .B(_03148__PTR18), .S(P2_P1_State2_PTR1), .Z(_03149__PTR2) );
  MUX2_X1 U24892 ( .A(1'b0), .B(_03148__PTR19), .S(P2_P1_State2_PTR1), .Z(_03149__PTR3) );
  MUX2_X1 U24893 ( .A(1'b0), .B(_03148__PTR20), .S(P2_P1_State2_PTR1), .Z(_03149__PTR4) );
  MUX2_X1 U24894 ( .A(1'b0), .B(_03148__PTR21), .S(P2_P1_State2_PTR1), .Z(_03149__PTR5) );
  MUX2_X1 U24895 ( .A(1'b0), .B(_03148__PTR22), .S(P2_P1_State2_PTR1), .Z(_03149__PTR6) );
  MUX2_X1 U24896 ( .A(1'b0), .B(_03148__PTR23), .S(P2_P1_State2_PTR1), .Z(_03149__PTR7) );
  MUX2_X1 U24897 ( .A(_03148__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03149__PTR32) );
  MUX2_X1 U24898 ( .A(_03148__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03149__PTR33) );
  MUX2_X1 U24899 ( .A(_03148__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03149__PTR34) );
  MUX2_X1 U24900 ( .A(_03148__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03149__PTR35) );
  MUX2_X1 U24901 ( .A(_03148__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03149__PTR36) );
  MUX2_X1 U24902 ( .A(_03148__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03149__PTR37) );
  MUX2_X1 U24903 ( .A(_03148__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03149__PTR38) );
  MUX2_X1 U24904 ( .A(_03148__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03149__PTR39) );
  MUX2_X1 U24905 ( .A(_02216__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR16) );
  MUX2_X1 U24906 ( .A(_02216__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR17) );
  MUX2_X1 U24907 ( .A(_02216__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR18) );
  MUX2_X1 U24908 ( .A(_02216__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR19) );
  MUX2_X1 U24909 ( .A(_02216__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR20) );
  MUX2_X1 U24910 ( .A(_02216__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR21) );
  MUX2_X1 U24911 ( .A(_02216__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR22) );
  MUX2_X1 U24912 ( .A(_02216__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR23) );
  MUX2_X1 U24913 ( .A(_02216__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR32) );
  MUX2_X1 U24914 ( .A(_02216__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR33) );
  MUX2_X1 U24915 ( .A(_02216__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR34) );
  MUX2_X1 U24916 ( .A(_02216__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR35) );
  MUX2_X1 U24917 ( .A(_02216__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR36) );
  MUX2_X1 U24918 ( .A(_02216__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR37) );
  MUX2_X1 U24919 ( .A(_02216__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR38) );
  MUX2_X1 U24920 ( .A(_02216__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR39) );
  MUX2_X1 U24921 ( .A(_02216__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR64) );
  MUX2_X1 U24922 ( .A(_02216__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR65) );
  MUX2_X1 U24923 ( .A(_02216__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR66) );
  MUX2_X1 U24924 ( .A(_02216__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR67) );
  MUX2_X1 U24925 ( .A(_02216__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR68) );
  MUX2_X1 U24926 ( .A(_02216__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR69) );
  MUX2_X1 U24927 ( .A(_02216__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR70) );
  MUX2_X1 U24928 ( .A(_02216__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03148__PTR71) );
  MUX2_X1 U24929 ( .A(_03153__PTR0), .B(_03151__PTR64), .S(P2_P1_State2_PTR3), .Z(_02219__PTR0) );
  MUX2_X1 U24930 ( .A(_03153__PTR1), .B(_03151__PTR65), .S(P2_P1_State2_PTR3), .Z(_02219__PTR1) );
  MUX2_X1 U24931 ( .A(_03153__PTR2), .B(_03151__PTR66), .S(P2_P1_State2_PTR3), .Z(_02219__PTR2) );
  MUX2_X1 U24932 ( .A(_03153__PTR3), .B(_03151__PTR67), .S(P2_P1_State2_PTR3), .Z(_02219__PTR3) );
  MUX2_X1 U24933 ( .A(_03153__PTR4), .B(_03151__PTR68), .S(P2_P1_State2_PTR3), .Z(_02219__PTR4) );
  MUX2_X1 U24934 ( .A(_03153__PTR5), .B(_03151__PTR69), .S(P2_P1_State2_PTR3), .Z(_02219__PTR5) );
  MUX2_X1 U24935 ( .A(_03153__PTR6), .B(_03151__PTR70), .S(P2_P1_State2_PTR3), .Z(_02219__PTR6) );
  MUX2_X1 U24936 ( .A(_03153__PTR7), .B(_03151__PTR71), .S(P2_P1_State2_PTR3), .Z(_02219__PTR7) );
  MUX2_X1 U24937 ( .A(_03152__PTR0), .B(_03152__PTR32), .S(P2_P1_State2_PTR2), .Z(_03153__PTR0) );
  MUX2_X1 U24938 ( .A(_03152__PTR1), .B(_03152__PTR33), .S(P2_P1_State2_PTR2), .Z(_03153__PTR1) );
  MUX2_X1 U24939 ( .A(_03152__PTR2), .B(_03152__PTR34), .S(P2_P1_State2_PTR2), .Z(_03153__PTR2) );
  MUX2_X1 U24940 ( .A(_03152__PTR3), .B(_03152__PTR35), .S(P2_P1_State2_PTR2), .Z(_03153__PTR3) );
  MUX2_X1 U24941 ( .A(_03152__PTR4), .B(_03152__PTR36), .S(P2_P1_State2_PTR2), .Z(_03153__PTR4) );
  MUX2_X1 U24942 ( .A(_03152__PTR5), .B(_03152__PTR37), .S(P2_P1_State2_PTR2), .Z(_03153__PTR5) );
  MUX2_X1 U24943 ( .A(_03152__PTR6), .B(_03152__PTR38), .S(P2_P1_State2_PTR2), .Z(_03153__PTR6) );
  MUX2_X1 U24944 ( .A(_03152__PTR7), .B(_03152__PTR39), .S(P2_P1_State2_PTR2), .Z(_03153__PTR7) );
  MUX2_X1 U24945 ( .A(1'b0), .B(_03151__PTR16), .S(P2_P1_State2_PTR1), .Z(_03152__PTR0) );
  MUX2_X1 U24946 ( .A(1'b0), .B(_03151__PTR17), .S(P2_P1_State2_PTR1), .Z(_03152__PTR1) );
  MUX2_X1 U24947 ( .A(1'b0), .B(_03151__PTR18), .S(P2_P1_State2_PTR1), .Z(_03152__PTR2) );
  MUX2_X1 U24948 ( .A(1'b0), .B(_03151__PTR19), .S(P2_P1_State2_PTR1), .Z(_03152__PTR3) );
  MUX2_X1 U24949 ( .A(1'b0), .B(_03151__PTR20), .S(P2_P1_State2_PTR1), .Z(_03152__PTR4) );
  MUX2_X1 U24950 ( .A(1'b0), .B(_03151__PTR21), .S(P2_P1_State2_PTR1), .Z(_03152__PTR5) );
  MUX2_X1 U24951 ( .A(1'b0), .B(_03151__PTR22), .S(P2_P1_State2_PTR1), .Z(_03152__PTR6) );
  MUX2_X1 U24952 ( .A(1'b0), .B(_03151__PTR23), .S(P2_P1_State2_PTR1), .Z(_03152__PTR7) );
  MUX2_X1 U24953 ( .A(_03151__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03152__PTR32) );
  MUX2_X1 U24954 ( .A(_03151__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03152__PTR33) );
  MUX2_X1 U24955 ( .A(_03151__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03152__PTR34) );
  MUX2_X1 U24956 ( .A(_03151__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03152__PTR35) );
  MUX2_X1 U24957 ( .A(_03151__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03152__PTR36) );
  MUX2_X1 U24958 ( .A(_03151__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03152__PTR37) );
  MUX2_X1 U24959 ( .A(_03151__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03152__PTR38) );
  MUX2_X1 U24960 ( .A(_03151__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03152__PTR39) );
  MUX2_X1 U24961 ( .A(_02218__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR16) );
  MUX2_X1 U24962 ( .A(_02218__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR17) );
  MUX2_X1 U24963 ( .A(_02218__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR18) );
  MUX2_X1 U24964 ( .A(_02218__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR19) );
  MUX2_X1 U24965 ( .A(_02218__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR20) );
  MUX2_X1 U24966 ( .A(_02218__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR21) );
  MUX2_X1 U24967 ( .A(_02218__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR22) );
  MUX2_X1 U24968 ( .A(_02218__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR23) );
  MUX2_X1 U24969 ( .A(_02218__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR32) );
  MUX2_X1 U24970 ( .A(_02218__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR33) );
  MUX2_X1 U24971 ( .A(_02218__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR34) );
  MUX2_X1 U24972 ( .A(_02218__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR35) );
  MUX2_X1 U24973 ( .A(_02218__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR36) );
  MUX2_X1 U24974 ( .A(_02218__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR37) );
  MUX2_X1 U24975 ( .A(_02218__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR38) );
  MUX2_X1 U24976 ( .A(_02218__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR39) );
  MUX2_X1 U24977 ( .A(_02218__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR64) );
  MUX2_X1 U24978 ( .A(_02218__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR65) );
  MUX2_X1 U24979 ( .A(_02218__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR66) );
  MUX2_X1 U24980 ( .A(_02218__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR67) );
  MUX2_X1 U24981 ( .A(_02218__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR68) );
  MUX2_X1 U24982 ( .A(_02218__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR69) );
  MUX2_X1 U24983 ( .A(_02218__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR70) );
  MUX2_X1 U24984 ( .A(_02218__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03151__PTR71) );
  MUX2_X1 U24985 ( .A(_03156__PTR0), .B(_03154__PTR64), .S(P2_P1_State2_PTR3), .Z(_02221__PTR0) );
  MUX2_X1 U24986 ( .A(_03156__PTR1), .B(_03154__PTR65), .S(P2_P1_State2_PTR3), .Z(_02221__PTR1) );
  MUX2_X1 U24987 ( .A(_03156__PTR2), .B(_03154__PTR66), .S(P2_P1_State2_PTR3), .Z(_02221__PTR2) );
  MUX2_X1 U24988 ( .A(_03156__PTR3), .B(_03154__PTR67), .S(P2_P1_State2_PTR3), .Z(_02221__PTR3) );
  MUX2_X1 U24989 ( .A(_03156__PTR4), .B(_03154__PTR68), .S(P2_P1_State2_PTR3), .Z(_02221__PTR4) );
  MUX2_X1 U24990 ( .A(_03156__PTR5), .B(_03154__PTR69), .S(P2_P1_State2_PTR3), .Z(_02221__PTR5) );
  MUX2_X1 U24991 ( .A(_03156__PTR6), .B(_03154__PTR70), .S(P2_P1_State2_PTR3), .Z(_02221__PTR6) );
  MUX2_X1 U24992 ( .A(_03156__PTR7), .B(_03154__PTR71), .S(P2_P1_State2_PTR3), .Z(_02221__PTR7) );
  MUX2_X1 U24993 ( .A(_03155__PTR0), .B(_03155__PTR32), .S(P2_P1_State2_PTR2), .Z(_03156__PTR0) );
  MUX2_X1 U24994 ( .A(_03155__PTR1), .B(_03155__PTR33), .S(P2_P1_State2_PTR2), .Z(_03156__PTR1) );
  MUX2_X1 U24995 ( .A(_03155__PTR2), .B(_03155__PTR34), .S(P2_P1_State2_PTR2), .Z(_03156__PTR2) );
  MUX2_X1 U24996 ( .A(_03155__PTR3), .B(_03155__PTR35), .S(P2_P1_State2_PTR2), .Z(_03156__PTR3) );
  MUX2_X1 U24997 ( .A(_03155__PTR4), .B(_03155__PTR36), .S(P2_P1_State2_PTR2), .Z(_03156__PTR4) );
  MUX2_X1 U24998 ( .A(_03155__PTR5), .B(_03155__PTR37), .S(P2_P1_State2_PTR2), .Z(_03156__PTR5) );
  MUX2_X1 U24999 ( .A(_03155__PTR6), .B(_03155__PTR38), .S(P2_P1_State2_PTR2), .Z(_03156__PTR6) );
  MUX2_X1 U25000 ( .A(_03155__PTR7), .B(_03155__PTR39), .S(P2_P1_State2_PTR2), .Z(_03156__PTR7) );
  MUX2_X1 U25001 ( .A(1'b0), .B(_03154__PTR16), .S(P2_P1_State2_PTR1), .Z(_03155__PTR0) );
  MUX2_X1 U25002 ( .A(1'b0), .B(_03154__PTR17), .S(P2_P1_State2_PTR1), .Z(_03155__PTR1) );
  MUX2_X1 U25003 ( .A(1'b0), .B(_03154__PTR18), .S(P2_P1_State2_PTR1), .Z(_03155__PTR2) );
  MUX2_X1 U25004 ( .A(1'b0), .B(_03154__PTR19), .S(P2_P1_State2_PTR1), .Z(_03155__PTR3) );
  MUX2_X1 U25005 ( .A(1'b0), .B(_03154__PTR20), .S(P2_P1_State2_PTR1), .Z(_03155__PTR4) );
  MUX2_X1 U25006 ( .A(1'b0), .B(_03154__PTR21), .S(P2_P1_State2_PTR1), .Z(_03155__PTR5) );
  MUX2_X1 U25007 ( .A(1'b0), .B(_03154__PTR22), .S(P2_P1_State2_PTR1), .Z(_03155__PTR6) );
  MUX2_X1 U25008 ( .A(1'b0), .B(_03154__PTR23), .S(P2_P1_State2_PTR1), .Z(_03155__PTR7) );
  MUX2_X1 U25009 ( .A(_03154__PTR32), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03155__PTR32) );
  MUX2_X1 U25010 ( .A(_03154__PTR33), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03155__PTR33) );
  MUX2_X1 U25011 ( .A(_03154__PTR34), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03155__PTR34) );
  MUX2_X1 U25012 ( .A(_03154__PTR35), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03155__PTR35) );
  MUX2_X1 U25013 ( .A(_03154__PTR36), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03155__PTR36) );
  MUX2_X1 U25014 ( .A(_03154__PTR37), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03155__PTR37) );
  MUX2_X1 U25015 ( .A(_03154__PTR38), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03155__PTR38) );
  MUX2_X1 U25016 ( .A(_03154__PTR39), .B(1'b0), .S(P2_P1_State2_PTR1), .Z(_03155__PTR39) );
  MUX2_X1 U25017 ( .A(_02220__PTR16), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR16) );
  MUX2_X1 U25018 ( .A(_02220__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR17) );
  MUX2_X1 U25019 ( .A(_02220__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR18) );
  MUX2_X1 U25020 ( .A(_02220__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR19) );
  MUX2_X1 U25021 ( .A(_02220__PTR20), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR20) );
  MUX2_X1 U25022 ( .A(_02220__PTR21), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR21) );
  MUX2_X1 U25023 ( .A(_02220__PTR22), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR22) );
  MUX2_X1 U25024 ( .A(_02220__PTR23), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR23) );
  MUX2_X1 U25025 ( .A(_02220__PTR32), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR32) );
  MUX2_X1 U25026 ( .A(_02220__PTR33), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR33) );
  MUX2_X1 U25027 ( .A(_02220__PTR34), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR34) );
  MUX2_X1 U25028 ( .A(_02220__PTR35), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR35) );
  MUX2_X1 U25029 ( .A(_02220__PTR36), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR36) );
  MUX2_X1 U25030 ( .A(_02220__PTR37), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR37) );
  MUX2_X1 U25031 ( .A(_02220__PTR38), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR38) );
  MUX2_X1 U25032 ( .A(_02220__PTR39), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR39) );
  MUX2_X1 U25033 ( .A(_02220__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR64) );
  MUX2_X1 U25034 ( .A(_02220__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR65) );
  MUX2_X1 U25035 ( .A(_02220__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR66) );
  MUX2_X1 U25036 ( .A(_02220__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR67) );
  MUX2_X1 U25037 ( .A(_02220__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR68) );
  MUX2_X1 U25038 ( .A(_02220__PTR69), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR69) );
  MUX2_X1 U25039 ( .A(_02220__PTR70), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR70) );
  MUX2_X1 U25040 ( .A(_02220__PTR71), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03154__PTR71) );
  MUX2_X1 U25041 ( .A(_03159__PTR0), .B(_03157__PTR64), .S(P2_P1_State2_PTR3), .Z(_02223__PTR0) );
  MUX2_X1 U25042 ( .A(_03159__PTR1), .B(_03157__PTR65), .S(P2_P1_State2_PTR3), .Z(_02223__PTR1) );
  MUX2_X1 U25043 ( .A(_03159__PTR2), .B(_03157__PTR66), .S(P2_P1_State2_PTR3), .Z(_02223__PTR2) );
  MUX2_X1 U25044 ( .A(_03159__PTR3), .B(_03157__PTR67), .S(P2_P1_State2_PTR3), .Z(_02223__PTR3) );
  MUX2_X1 U25045 ( .A(_03159__PTR4), .B(_03157__PTR68), .S(P2_P1_State2_PTR3), .Z(_02223__PTR4) );
  MUX2_X1 U25046 ( .A(1'b0), .B(_03158__PTR32), .S(P2_P1_State2_PTR2), .Z(_03159__PTR0) );
  MUX2_X1 U25047 ( .A(_03158__PTR1), .B(_03158__PTR33), .S(P2_P1_State2_PTR2), .Z(_03159__PTR1) );
  MUX2_X1 U25048 ( .A(_03158__PTR2), .B(_03158__PTR34), .S(P2_P1_State2_PTR2), .Z(_03159__PTR2) );
  MUX2_X1 U25049 ( .A(_03158__PTR3), .B(_03158__PTR35), .S(P2_P1_State2_PTR2), .Z(_03159__PTR3) );
  MUX2_X1 U25050 ( .A(_03158__PTR4), .B(_03158__PTR36), .S(P2_P1_State2_PTR2), .Z(_03159__PTR4) );
  MUX2_X1 U25051 ( .A(1'b0), .B(_03157__PTR17), .S(P2_P1_State2_PTR1), .Z(_03158__PTR1) );
  MUX2_X1 U25052 ( .A(1'b0), .B(_03157__PTR18), .S(P2_P1_State2_PTR1), .Z(_03158__PTR2) );
  MUX2_X1 U25053 ( .A(1'b0), .B(_03157__PTR19), .S(P2_P1_State2_PTR1), .Z(_03158__PTR3) );
  MUX2_X1 U25054 ( .A(1'b0), .B(_03157__PTR36), .S(P2_P1_State2_PTR1), .Z(_03158__PTR4) );
  MUX2_X1 U25055 ( .A(1'b0), .B(_03157__PTR48), .S(P2_P1_State2_PTR1), .Z(_03158__PTR32) );
  MUX2_X1 U25056 ( .A(_03157__PTR33), .B(_03157__PTR52), .S(P2_P1_State2_PTR1), .Z(_03158__PTR33) );
  MUX2_X1 U25057 ( .A(_03157__PTR34), .B(_03157__PTR52), .S(P2_P1_State2_PTR1), .Z(_03158__PTR34) );
  MUX2_X1 U25058 ( .A(_03157__PTR35), .B(_03157__PTR52), .S(P2_P1_State2_PTR1), .Z(_03158__PTR35) );
  MUX2_X1 U25059 ( .A(_03157__PTR36), .B(_03157__PTR52), .S(P2_P1_State2_PTR1), .Z(_03158__PTR36) );
  MUX2_X1 U25060 ( .A(_02222__PTR17), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03157__PTR17) );
  MUX2_X1 U25061 ( .A(_02222__PTR18), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03157__PTR18) );
  MUX2_X1 U25062 ( .A(_02222__PTR19), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03157__PTR19) );
  MUX2_X1 U25063 ( .A(_02131__PTR1), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03157__PTR33) );
  MUX2_X1 U25064 ( .A(_02131__PTR2), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03157__PTR34) );
  MUX2_X1 U25065 ( .A(_02131__PTR3), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03157__PTR35) );
  MUX2_X1 U25066 ( .A(1'b0), .B(P2_P1_InstQueueWr_Addr_PTR4), .S(P2_P1_State2_PTR0), .Z(_03157__PTR36) );
  MUX2_X1 U25067 ( .A(1'b0), .B(_02222__PTR56), .S(P2_P1_State2_PTR0), .Z(_03157__PTR48) );
  MUX2_X1 U25068 ( .A(1'b0), .B(_02222__PTR60), .S(P2_P1_State2_PTR0), .Z(_03157__PTR52) );
  MUX2_X1 U25069 ( .A(_02222__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03157__PTR64) );
  MUX2_X1 U25070 ( .A(_02222__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03157__PTR65) );
  MUX2_X1 U25071 ( .A(_02222__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03157__PTR66) );
  MUX2_X1 U25072 ( .A(_02222__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03157__PTR67) );
  MUX2_X1 U25073 ( .A(_02222__PTR68), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03157__PTR68) );
  MUX2_X1 U25074 ( .A(_03162__PTR0), .B(_03160__PTR64), .S(P2_P1_State2_PTR3), .Z(_02225__PTR0) );
  MUX2_X1 U25075 ( .A(_03162__PTR1), .B(_03160__PTR65), .S(P2_P1_State2_PTR3), .Z(_02225__PTR1) );
  MUX2_X1 U25076 ( .A(_03162__PTR2), .B(_03160__PTR66), .S(P2_P1_State2_PTR3), .Z(_02225__PTR2) );
  MUX2_X1 U25077 ( .A(_03162__PTR3), .B(_03160__PTR67), .S(P2_P1_State2_PTR3), .Z(_02225__PTR3) );
  MUX2_X1 U25078 ( .A(_03162__PTR4), .B(_03106__PTR32), .S(P2_P1_State2_PTR3), .Z(_02225__PTR4) );
  MUX2_X1 U25079 ( .A(1'b0), .B(_03161__PTR32), .S(P2_P1_State2_PTR2), .Z(_03162__PTR0) );
  MUX2_X1 U25080 ( .A(1'b0), .B(_03161__PTR33), .S(P2_P1_State2_PTR2), .Z(_03162__PTR1) );
  MUX2_X1 U25081 ( .A(1'b0), .B(_03161__PTR34), .S(P2_P1_State2_PTR2), .Z(_03162__PTR2) );
  MUX2_X1 U25082 ( .A(1'b0), .B(_03161__PTR35), .S(P2_P1_State2_PTR2), .Z(_03162__PTR3) );
  MUX2_X1 U25083 ( .A(1'b0), .B(_03161__PTR36), .S(P2_P1_State2_PTR2), .Z(_03162__PTR4) );
  MUX2_X1 U25084 ( .A(_03160__PTR32), .B(_03160__PTR48), .S(P2_P1_State2_PTR1), .Z(_03161__PTR32) );
  MUX2_X1 U25085 ( .A(_03160__PTR33), .B(_03160__PTR49), .S(P2_P1_State2_PTR1), .Z(_03161__PTR33) );
  MUX2_X1 U25086 ( .A(_03160__PTR34), .B(_03160__PTR50), .S(P2_P1_State2_PTR1), .Z(_03161__PTR34) );
  MUX2_X1 U25087 ( .A(_03160__PTR35), .B(_03160__PTR51), .S(P2_P1_State2_PTR1), .Z(_03161__PTR35) );
  MUX2_X1 U25088 ( .A(_03160__PTR36), .B(_03160__PTR52), .S(P2_P1_State2_PTR1), .Z(_03161__PTR36) );
  MUX2_X1 U25089 ( .A(1'b0), .B(_02224__PTR40), .S(P2_P1_State2_PTR0), .Z(_03160__PTR32) );
  MUX2_X1 U25090 ( .A(1'b0), .B(_02224__PTR41), .S(P2_P1_State2_PTR0), .Z(_03160__PTR33) );
  MUX2_X1 U25091 ( .A(1'b0), .B(_02224__PTR42), .S(P2_P1_State2_PTR0), .Z(_03160__PTR34) );
  MUX2_X1 U25092 ( .A(1'b0), .B(_02224__PTR43), .S(P2_P1_State2_PTR0), .Z(_03160__PTR35) );
  MUX2_X1 U25093 ( .A(1'b0), .B(_02224__PTR44), .S(P2_P1_State2_PTR0), .Z(_03160__PTR36) );
  MUX2_X1 U25094 ( .A(1'b0), .B(_02224__PTR56), .S(P2_P1_State2_PTR0), .Z(_03160__PTR48) );
  MUX2_X1 U25095 ( .A(1'b0), .B(_02224__PTR57), .S(P2_P1_State2_PTR0), .Z(_03160__PTR49) );
  MUX2_X1 U25096 ( .A(1'b0), .B(_02224__PTR58), .S(P2_P1_State2_PTR0), .Z(_03160__PTR50) );
  MUX2_X1 U25097 ( .A(1'b0), .B(_02224__PTR59), .S(P2_P1_State2_PTR0), .Z(_03160__PTR51) );
  MUX2_X1 U25098 ( .A(1'b0), .B(_02224__PTR60), .S(P2_P1_State2_PTR0), .Z(_03160__PTR52) );
  MUX2_X1 U25099 ( .A(_02224__PTR64), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03160__PTR64) );
  MUX2_X1 U25100 ( .A(_02224__PTR65), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03160__PTR65) );
  MUX2_X1 U25101 ( .A(_02224__PTR66), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03160__PTR66) );
  MUX2_X1 U25102 ( .A(_02224__PTR67), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03160__PTR67) );
  MUX2_X1 U25103 ( .A(_03163__PTR256), .B(_03163__PTR384), .S(P2_P1_State2_PTR1), .Z(_03164__PTR256) );
  MUX2_X1 U25104 ( .A(_03163__PTR257), .B(_03163__PTR385), .S(P2_P1_State2_PTR1), .Z(_03164__PTR257) );
  MUX2_X1 U25105 ( .A(_03163__PTR258), .B(_03163__PTR386), .S(P2_P1_State2_PTR1), .Z(_03164__PTR258) );
  MUX2_X1 U25106 ( .A(_03163__PTR259), .B(_03163__PTR387), .S(P2_P1_State2_PTR1), .Z(_03164__PTR259) );
  MUX2_X1 U25107 ( .A(_03163__PTR260), .B(_03163__PTR388), .S(P2_P1_State2_PTR1), .Z(_03164__PTR260) );
  MUX2_X1 U25108 ( .A(_03163__PTR261), .B(_03163__PTR389), .S(P2_P1_State2_PTR1), .Z(_03164__PTR261) );
  MUX2_X1 U25109 ( .A(_03163__PTR262), .B(_03163__PTR390), .S(P2_P1_State2_PTR1), .Z(_03164__PTR262) );
  MUX2_X1 U25110 ( .A(_03163__PTR263), .B(_03163__PTR391), .S(P2_P1_State2_PTR1), .Z(_03164__PTR263) );
  MUX2_X1 U25111 ( .A(_03163__PTR264), .B(_03163__PTR392), .S(P2_P1_State2_PTR1), .Z(_03164__PTR264) );
  MUX2_X1 U25112 ( .A(_03163__PTR265), .B(_03163__PTR393), .S(P2_P1_State2_PTR1), .Z(_03164__PTR265) );
  MUX2_X1 U25113 ( .A(_03163__PTR266), .B(_03163__PTR394), .S(P2_P1_State2_PTR1), .Z(_03164__PTR266) );
  MUX2_X1 U25114 ( .A(_03163__PTR267), .B(_03163__PTR395), .S(P2_P1_State2_PTR1), .Z(_03164__PTR267) );
  MUX2_X1 U25115 ( .A(_03163__PTR268), .B(_03163__PTR396), .S(P2_P1_State2_PTR1), .Z(_03164__PTR268) );
  MUX2_X1 U25116 ( .A(_03163__PTR269), .B(_03163__PTR397), .S(P2_P1_State2_PTR1), .Z(_03164__PTR269) );
  MUX2_X1 U25117 ( .A(_03163__PTR270), .B(_03163__PTR398), .S(P2_P1_State2_PTR1), .Z(_03164__PTR270) );
  MUX2_X1 U25118 ( .A(_03163__PTR271), .B(_03163__PTR399), .S(P2_P1_State2_PTR1), .Z(_03164__PTR271) );
  MUX2_X1 U25119 ( .A(_03163__PTR272), .B(_03163__PTR400), .S(P2_P1_State2_PTR1), .Z(_03164__PTR272) );
  MUX2_X1 U25120 ( .A(_03163__PTR273), .B(_03163__PTR401), .S(P2_P1_State2_PTR1), .Z(_03164__PTR273) );
  MUX2_X1 U25121 ( .A(_03163__PTR274), .B(_03163__PTR402), .S(P2_P1_State2_PTR1), .Z(_03164__PTR274) );
  MUX2_X1 U25122 ( .A(_03163__PTR275), .B(_03163__PTR403), .S(P2_P1_State2_PTR1), .Z(_03164__PTR275) );
  MUX2_X1 U25123 ( .A(_03163__PTR276), .B(_03163__PTR404), .S(P2_P1_State2_PTR1), .Z(_03164__PTR276) );
  MUX2_X1 U25124 ( .A(_03163__PTR277), .B(_03163__PTR405), .S(P2_P1_State2_PTR1), .Z(_03164__PTR277) );
  MUX2_X1 U25125 ( .A(_03163__PTR278), .B(_03163__PTR406), .S(P2_P1_State2_PTR1), .Z(_03164__PTR278) );
  MUX2_X1 U25126 ( .A(_03163__PTR279), .B(_03163__PTR407), .S(P2_P1_State2_PTR1), .Z(_03164__PTR279) );
  MUX2_X1 U25127 ( .A(_03163__PTR280), .B(_03163__PTR408), .S(P2_P1_State2_PTR1), .Z(_03164__PTR280) );
  MUX2_X1 U25128 ( .A(_03163__PTR281), .B(_03163__PTR409), .S(P2_P1_State2_PTR1), .Z(_03164__PTR281) );
  MUX2_X1 U25129 ( .A(_03163__PTR282), .B(_03163__PTR410), .S(P2_P1_State2_PTR1), .Z(_03164__PTR282) );
  MUX2_X1 U25130 ( .A(_03163__PTR283), .B(_03163__PTR411), .S(P2_P1_State2_PTR1), .Z(_03164__PTR283) );
  MUX2_X1 U25131 ( .A(_03163__PTR284), .B(_03163__PTR412), .S(P2_P1_State2_PTR1), .Z(_03164__PTR284) );
  MUX2_X1 U25132 ( .A(_03163__PTR285), .B(_03163__PTR413), .S(P2_P1_State2_PTR1), .Z(_03164__PTR285) );
  MUX2_X1 U25133 ( .A(_03163__PTR286), .B(_03163__PTR414), .S(P2_P1_State2_PTR1), .Z(_03164__PTR286) );
  MUX2_X1 U25134 ( .A(_03163__PTR288), .B(_03106__PTR32), .S(P2_P1_State2_PTR1), .Z(_03164__PTR288) );
  MUX2_X1 U25135 ( .A(1'b0), .B(_02230__PTR320), .S(P2_P1_State2_PTR0), .Z(_03163__PTR256) );
  MUX2_X1 U25136 ( .A(1'b0), .B(_02230__PTR321), .S(P2_P1_State2_PTR0), .Z(_03163__PTR257) );
  MUX2_X1 U25137 ( .A(1'b0), .B(_02230__PTR322), .S(P2_P1_State2_PTR0), .Z(_03163__PTR258) );
  MUX2_X1 U25138 ( .A(1'b0), .B(_02230__PTR323), .S(P2_P1_State2_PTR0), .Z(_03163__PTR259) );
  MUX2_X1 U25139 ( .A(1'b0), .B(_02230__PTR324), .S(P2_P1_State2_PTR0), .Z(_03163__PTR260) );
  MUX2_X1 U25140 ( .A(1'b0), .B(_02230__PTR325), .S(P2_P1_State2_PTR0), .Z(_03163__PTR261) );
  MUX2_X1 U25141 ( .A(1'b0), .B(_02230__PTR326), .S(P2_P1_State2_PTR0), .Z(_03163__PTR262) );
  MUX2_X1 U25142 ( .A(1'b0), .B(_02230__PTR327), .S(P2_P1_State2_PTR0), .Z(_03163__PTR263) );
  MUX2_X1 U25143 ( .A(1'b0), .B(_02230__PTR328), .S(P2_P1_State2_PTR0), .Z(_03163__PTR264) );
  MUX2_X1 U25144 ( .A(1'b0), .B(_02230__PTR329), .S(P2_P1_State2_PTR0), .Z(_03163__PTR265) );
  MUX2_X1 U25145 ( .A(1'b0), .B(_02230__PTR330), .S(P2_P1_State2_PTR0), .Z(_03163__PTR266) );
  MUX2_X1 U25146 ( .A(1'b0), .B(_02230__PTR331), .S(P2_P1_State2_PTR0), .Z(_03163__PTR267) );
  MUX2_X1 U25147 ( .A(1'b0), .B(_02230__PTR332), .S(P2_P1_State2_PTR0), .Z(_03163__PTR268) );
  MUX2_X1 U25148 ( .A(1'b0), .B(_02230__PTR333), .S(P2_P1_State2_PTR0), .Z(_03163__PTR269) );
  MUX2_X1 U25149 ( .A(1'b0), .B(_02230__PTR334), .S(P2_P1_State2_PTR0), .Z(_03163__PTR270) );
  MUX2_X1 U25150 ( .A(1'b0), .B(_02230__PTR335), .S(P2_P1_State2_PTR0), .Z(_03163__PTR271) );
  MUX2_X1 U25151 ( .A(1'b0), .B(_02230__PTR336), .S(P2_P1_State2_PTR0), .Z(_03163__PTR272) );
  MUX2_X1 U25152 ( .A(1'b0), .B(_02230__PTR337), .S(P2_P1_State2_PTR0), .Z(_03163__PTR273) );
  MUX2_X1 U25153 ( .A(1'b0), .B(_02230__PTR338), .S(P2_P1_State2_PTR0), .Z(_03163__PTR274) );
  MUX2_X1 U25154 ( .A(1'b0), .B(_02230__PTR339), .S(P2_P1_State2_PTR0), .Z(_03163__PTR275) );
  MUX2_X1 U25155 ( .A(1'b0), .B(_02230__PTR340), .S(P2_P1_State2_PTR0), .Z(_03163__PTR276) );
  MUX2_X1 U25156 ( .A(1'b0), .B(_02230__PTR341), .S(P2_P1_State2_PTR0), .Z(_03163__PTR277) );
  MUX2_X1 U25157 ( .A(1'b0), .B(_02230__PTR342), .S(P2_P1_State2_PTR0), .Z(_03163__PTR278) );
  MUX2_X1 U25158 ( .A(1'b0), .B(_02230__PTR343), .S(P2_P1_State2_PTR0), .Z(_03163__PTR279) );
  MUX2_X1 U25159 ( .A(1'b0), .B(_02230__PTR344), .S(P2_P1_State2_PTR0), .Z(_03163__PTR280) );
  MUX2_X1 U25160 ( .A(1'b0), .B(_02230__PTR345), .S(P2_P1_State2_PTR0), .Z(_03163__PTR281) );
  MUX2_X1 U25161 ( .A(1'b0), .B(_02230__PTR346), .S(P2_P1_State2_PTR0), .Z(_03163__PTR282) );
  MUX2_X1 U25162 ( .A(1'b0), .B(_02230__PTR347), .S(P2_P1_State2_PTR0), .Z(_03163__PTR283) );
  MUX2_X1 U25163 ( .A(1'b0), .B(_02230__PTR348), .S(P2_P1_State2_PTR0), .Z(_03163__PTR284) );
  MUX2_X1 U25164 ( .A(1'b0), .B(_02230__PTR349), .S(P2_P1_State2_PTR0), .Z(_03163__PTR285) );
  MUX2_X1 U25165 ( .A(1'b0), .B(_02230__PTR350), .S(P2_P1_State2_PTR0), .Z(_03163__PTR286) );
  MUX2_X1 U25166 ( .A(1'b0), .B(_02230__PTR352), .S(P2_P1_State2_PTR0), .Z(_03163__PTR288) );
  MUX2_X1 U25167 ( .A(P2_P1_lWord_PTR0), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR384) );
  MUX2_X1 U25168 ( .A(P2_P1_lWord_PTR1), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR385) );
  MUX2_X1 U25169 ( .A(P2_P1_lWord_PTR2), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR386) );
  MUX2_X1 U25170 ( .A(P2_P1_lWord_PTR3), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR387) );
  MUX2_X1 U25171 ( .A(P2_P1_lWord_PTR4), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR388) );
  MUX2_X1 U25172 ( .A(P2_P1_lWord_PTR5), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR389) );
  MUX2_X1 U25173 ( .A(P2_P1_lWord_PTR6), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR390) );
  MUX2_X1 U25174 ( .A(P2_P1_lWord_PTR7), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR391) );
  MUX2_X1 U25175 ( .A(P2_P1_lWord_PTR8), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR392) );
  MUX2_X1 U25176 ( .A(P2_P1_lWord_PTR9), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR393) );
  MUX2_X1 U25177 ( .A(P2_P1_lWord_PTR10), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR394) );
  MUX2_X1 U25178 ( .A(P2_P1_lWord_PTR11), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR395) );
  MUX2_X1 U25179 ( .A(P2_P1_lWord_PTR12), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR396) );
  MUX2_X1 U25180 ( .A(P2_P1_lWord_PTR13), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR397) );
  MUX2_X1 U25181 ( .A(P2_P1_lWord_PTR14), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR398) );
  MUX2_X1 U25182 ( .A(P2_P1_lWord_PTR15), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR399) );
  MUX2_X1 U25183 ( .A(P2_P1_uWord_PTR0), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR400) );
  MUX2_X1 U25184 ( .A(P2_P1_uWord_PTR1), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR401) );
  MUX2_X1 U25185 ( .A(P2_P1_uWord_PTR2), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR402) );
  MUX2_X1 U25186 ( .A(P2_P1_uWord_PTR3), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR403) );
  MUX2_X1 U25187 ( .A(P2_P1_uWord_PTR4), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR404) );
  MUX2_X1 U25188 ( .A(P2_P1_uWord_PTR5), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR405) );
  MUX2_X1 U25189 ( .A(P2_P1_uWord_PTR6), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR406) );
  MUX2_X1 U25190 ( .A(P2_P1_uWord_PTR7), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR407) );
  MUX2_X1 U25191 ( .A(P2_P1_uWord_PTR8), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR408) );
  MUX2_X1 U25192 ( .A(P2_P1_uWord_PTR9), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR409) );
  MUX2_X1 U25193 ( .A(P2_P1_uWord_PTR10), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR410) );
  MUX2_X1 U25194 ( .A(P2_P1_uWord_PTR11), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR411) );
  MUX2_X1 U25195 ( .A(P2_P1_uWord_PTR12), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR412) );
  MUX2_X1 U25196 ( .A(P2_P1_uWord_PTR13), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR413) );
  MUX2_X1 U25197 ( .A(P2_P1_uWord_PTR14), .B(1'b0), .S(P2_P1_State2_PTR0), .Z(_03163__PTR414) );
  MUX2_X1 U25198 ( .A(_03196__PTR0), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR0) );
  MUX2_X1 U25199 ( .A(_03196__PTR1), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR1) );
  MUX2_X1 U25200 ( .A(_03196__PTR2), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR2) );
  MUX2_X1 U25201 ( .A(_03196__PTR3), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR3) );
  MUX2_X1 U25202 ( .A(_03196__PTR4), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR4) );
  MUX2_X1 U25203 ( .A(_03196__PTR5), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR5) );
  MUX2_X1 U25204 ( .A(_03196__PTR6), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR6) );
  MUX2_X1 U25205 ( .A(_03196__PTR7), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR7) );
  MUX2_X1 U25206 ( .A(1'b0), .B(_03196__PTR0), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR8) );
  MUX2_X1 U25207 ( .A(1'b0), .B(_03196__PTR1), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR9) );
  MUX2_X1 U25208 ( .A(1'b0), .B(_03196__PTR2), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR10) );
  MUX2_X1 U25209 ( .A(1'b0), .B(_03196__PTR3), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR11) );
  MUX2_X1 U25210 ( .A(1'b0), .B(_03196__PTR4), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR12) );
  MUX2_X1 U25211 ( .A(1'b0), .B(_03196__PTR5), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR13) );
  MUX2_X1 U25212 ( .A(1'b0), .B(_03196__PTR6), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR14) );
  MUX2_X1 U25213 ( .A(1'b0), .B(_03196__PTR7), .S(P3_P1_InstQueueWr_Addr_PTR3), .Z(_02417__PTR15) );
  MUX2_X1 U25214 ( .A(_03195__PTR0), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR2), .Z(_03196__PTR0) );
  MUX2_X1 U25215 ( .A(_03195__PTR1), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR2), .Z(_03196__PTR1) );
  MUX2_X1 U25216 ( .A(_03195__PTR2), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR2), .Z(_03196__PTR2) );
  MUX2_X1 U25217 ( .A(_03195__PTR3), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR2), .Z(_03196__PTR3) );
  MUX2_X1 U25218 ( .A(1'b0), .B(_03195__PTR0), .S(P3_P1_InstQueueWr_Addr_PTR2), .Z(_03196__PTR4) );
  MUX2_X1 U25219 ( .A(1'b0), .B(_03195__PTR1), .S(P3_P1_InstQueueWr_Addr_PTR2), .Z(_03196__PTR5) );
  MUX2_X1 U25220 ( .A(1'b0), .B(_03195__PTR2), .S(P3_P1_InstQueueWr_Addr_PTR2), .Z(_03196__PTR6) );
  MUX2_X1 U25221 ( .A(1'b0), .B(_03195__PTR3), .S(P3_P1_InstQueueWr_Addr_PTR2), .Z(_03196__PTR7) );
  MUX2_X1 U25222 ( .A(_02418__PTR0), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR1), .Z(_03195__PTR0) );
  MUX2_X1 U25223 ( .A(P3_P1_InstQueueWr_Addr_PTR0), .B(1'b0), .S(P3_P1_InstQueueWr_Addr_PTR1), .Z(_03195__PTR1) );
  MUX2_X1 U25224 ( .A(1'b0), .B(_02418__PTR0), .S(P3_P1_InstQueueWr_Addr_PTR1), .Z(_03195__PTR2) );
  MUX2_X1 U25225 ( .A(1'b0), .B(P3_P1_InstQueueWr_Addr_PTR0), .S(P3_P1_InstQueueWr_Addr_PTR1), .Z(_03195__PTR3) );
  MUX2_X1 U25226 ( .A(_03198__PTR0), .B(1'b0), .S(_02418__PTR3), .Z(_02419__PTR0) );
  MUX2_X1 U25227 ( .A(_03198__PTR1), .B(1'b0), .S(_02418__PTR3), .Z(_02419__PTR1) );
  MUX2_X1 U25228 ( .A(_03198__PTR2), .B(1'b0), .S(_02418__PTR3), .Z(_02419__PTR2) );
  MUX2_X1 U25229 ( .A(_03198__PTR3), .B(1'b0), .S(_02418__PTR3), .Z(_02419__PTR3) );
  MUX2_X1 U25230 ( .A(_03198__PTR4), .B(1'b0), .S(_02418__PTR3), .Z(_02419__PTR4) );
  MUX2_X1 U25231 ( .A(_03198__PTR5), .B(1'b0), .S(_02418__PTR3), .Z(_02419__PTR5) );
  MUX2_X1 U25232 ( .A(_03198__PTR6), .B(1'b0), .S(_02418__PTR3), .Z(_02419__PTR6) );
  MUX2_X1 U25233 ( .A(_03198__PTR7), .B(1'b0), .S(_02418__PTR3), .Z(_02419__PTR7) );
  MUX2_X1 U25234 ( .A(1'b0), .B(_03198__PTR0), .S(_02418__PTR3), .Z(_02419__PTR8) );
  MUX2_X1 U25235 ( .A(1'b0), .B(_03198__PTR1), .S(_02418__PTR3), .Z(_02419__PTR9) );
  MUX2_X1 U25236 ( .A(1'b0), .B(_03198__PTR2), .S(_02418__PTR3), .Z(_02419__PTR10) );
  MUX2_X1 U25237 ( .A(1'b0), .B(_03198__PTR3), .S(_02418__PTR3), .Z(_02419__PTR11) );
  MUX2_X1 U25238 ( .A(1'b0), .B(_03198__PTR4), .S(_02418__PTR3), .Z(_02419__PTR12) );
  MUX2_X1 U25239 ( .A(1'b0), .B(_03198__PTR5), .S(_02418__PTR3), .Z(_02419__PTR13) );
  MUX2_X1 U25240 ( .A(1'b0), .B(_03198__PTR6), .S(_02418__PTR3), .Z(_02419__PTR14) );
  MUX2_X1 U25241 ( .A(1'b0), .B(_03198__PTR7), .S(_02418__PTR3), .Z(_02419__PTR15) );
  MUX2_X1 U25242 ( .A(_03197__PTR0), .B(1'b0), .S(_02418__PTR2), .Z(_03198__PTR0) );
  MUX2_X1 U25243 ( .A(_03197__PTR1), .B(1'b0), .S(_02418__PTR2), .Z(_03198__PTR1) );
  MUX2_X1 U25244 ( .A(_03197__PTR2), .B(1'b0), .S(_02418__PTR2), .Z(_03198__PTR2) );
  MUX2_X1 U25245 ( .A(_03197__PTR3), .B(1'b0), .S(_02418__PTR2), .Z(_03198__PTR3) );
  MUX2_X1 U25246 ( .A(1'b0), .B(_03197__PTR0), .S(_02418__PTR2), .Z(_03198__PTR4) );
  MUX2_X1 U25247 ( .A(1'b0), .B(_03197__PTR1), .S(_02418__PTR2), .Z(_03198__PTR5) );
  MUX2_X1 U25248 ( .A(1'b0), .B(_03197__PTR2), .S(_02418__PTR2), .Z(_03198__PTR6) );
  MUX2_X1 U25249 ( .A(1'b0), .B(_03197__PTR3), .S(_02418__PTR2), .Z(_03198__PTR7) );
  MUX2_X1 U25250 ( .A(P3_P1_InstQueueWr_Addr_PTR0), .B(1'b0), .S(_02418__PTR1), .Z(_03197__PTR0) );
  MUX2_X1 U25251 ( .A(_02418__PTR0), .B(1'b0), .S(_02418__PTR1), .Z(_03197__PTR1) );
  MUX2_X1 U25252 ( .A(1'b0), .B(P3_P1_InstQueueWr_Addr_PTR0), .S(_02418__PTR1), .Z(_03197__PTR2) );
  MUX2_X1 U25253 ( .A(1'b0), .B(_02418__PTR0), .S(_02418__PTR1), .Z(_03197__PTR3) );
  MUX2_X1 U25254 ( .A(_03200__PTR0), .B(1'b0), .S(_02420__PTR3), .Z(_02421__PTR0) );
  MUX2_X1 U25255 ( .A(_03200__PTR1), .B(1'b0), .S(_02420__PTR3), .Z(_02421__PTR1) );
  MUX2_X1 U25256 ( .A(_03200__PTR2), .B(1'b0), .S(_02420__PTR3), .Z(_02421__PTR2) );
  MUX2_X1 U25257 ( .A(_03200__PTR3), .B(1'b0), .S(_02420__PTR3), .Z(_02421__PTR3) );
  MUX2_X1 U25258 ( .A(_03200__PTR4), .B(1'b0), .S(_02420__PTR3), .Z(_02421__PTR4) );
  MUX2_X1 U25259 ( .A(_03200__PTR5), .B(1'b0), .S(_02420__PTR3), .Z(_02421__PTR5) );
  MUX2_X1 U25260 ( .A(_03200__PTR6), .B(1'b0), .S(_02420__PTR3), .Z(_02421__PTR6) );
  MUX2_X1 U25261 ( .A(_03200__PTR7), .B(1'b0), .S(_02420__PTR3), .Z(_02421__PTR7) );
  MUX2_X1 U25262 ( .A(1'b0), .B(_03200__PTR0), .S(_02420__PTR3), .Z(_02421__PTR8) );
  MUX2_X1 U25263 ( .A(1'b0), .B(_03200__PTR1), .S(_02420__PTR3), .Z(_02421__PTR9) );
  MUX2_X1 U25264 ( .A(1'b0), .B(_03200__PTR2), .S(_02420__PTR3), .Z(_02421__PTR10) );
  MUX2_X1 U25265 ( .A(1'b0), .B(_03200__PTR3), .S(_02420__PTR3), .Z(_02421__PTR11) );
  MUX2_X1 U25266 ( .A(1'b0), .B(_03200__PTR4), .S(_02420__PTR3), .Z(_02421__PTR12) );
  MUX2_X1 U25267 ( .A(1'b0), .B(_03200__PTR5), .S(_02420__PTR3), .Z(_02421__PTR13) );
  MUX2_X1 U25268 ( .A(1'b0), .B(_03200__PTR6), .S(_02420__PTR3), .Z(_02421__PTR14) );
  MUX2_X1 U25269 ( .A(1'b0), .B(_03200__PTR7), .S(_02420__PTR3), .Z(_02421__PTR15) );
  MUX2_X1 U25270 ( .A(_03199__PTR0), .B(1'b0), .S(_02420__PTR2), .Z(_03200__PTR0) );
  MUX2_X1 U25271 ( .A(_03199__PTR1), .B(1'b0), .S(_02420__PTR2), .Z(_03200__PTR1) );
  MUX2_X1 U25272 ( .A(_03199__PTR2), .B(1'b0), .S(_02420__PTR2), .Z(_03200__PTR2) );
  MUX2_X1 U25273 ( .A(_03199__PTR3), .B(1'b0), .S(_02420__PTR2), .Z(_03200__PTR3) );
  MUX2_X1 U25274 ( .A(1'b0), .B(_03199__PTR0), .S(_02420__PTR2), .Z(_03200__PTR4) );
  MUX2_X1 U25275 ( .A(1'b0), .B(_03199__PTR1), .S(_02420__PTR2), .Z(_03200__PTR5) );
  MUX2_X1 U25276 ( .A(1'b0), .B(_03199__PTR2), .S(_02420__PTR2), .Z(_03200__PTR6) );
  MUX2_X1 U25277 ( .A(1'b0), .B(_03199__PTR3), .S(_02420__PTR2), .Z(_03200__PTR7) );
  MUX2_X1 U25278 ( .A(_02418__PTR0), .B(1'b0), .S(_02420__PTR1), .Z(_03199__PTR0) );
  MUX2_X1 U25279 ( .A(P3_P1_InstQueueWr_Addr_PTR0), .B(1'b0), .S(_02420__PTR1), .Z(_03199__PTR1) );
  MUX2_X1 U25280 ( .A(1'b0), .B(_02418__PTR0), .S(_02420__PTR1), .Z(_03199__PTR2) );
  MUX2_X1 U25281 ( .A(1'b0), .B(P3_P1_InstQueueWr_Addr_PTR0), .S(_02420__PTR1), .Z(_03199__PTR3) );
  MUX2_X1 U25282 ( .A(_03202__PTR0), .B(1'b0), .S(_02422__PTR3), .Z(_02423__PTR0) );
  MUX2_X1 U25283 ( .A(_03202__PTR1), .B(1'b0), .S(_02422__PTR3), .Z(_02423__PTR1) );
  MUX2_X1 U25284 ( .A(_03202__PTR2), .B(1'b0), .S(_02422__PTR3), .Z(_02423__PTR2) );
  MUX2_X1 U25285 ( .A(_03202__PTR3), .B(1'b0), .S(_02422__PTR3), .Z(_02423__PTR3) );
  MUX2_X1 U25286 ( .A(_03202__PTR4), .B(1'b0), .S(_02422__PTR3), .Z(_02423__PTR4) );
  MUX2_X1 U25287 ( .A(_03202__PTR5), .B(1'b0), .S(_02422__PTR3), .Z(_02423__PTR5) );
  MUX2_X1 U25288 ( .A(_03202__PTR6), .B(1'b0), .S(_02422__PTR3), .Z(_02423__PTR6) );
  MUX2_X1 U25289 ( .A(_03202__PTR7), .B(1'b0), .S(_02422__PTR3), .Z(_02423__PTR7) );
  MUX2_X1 U25290 ( .A(1'b0), .B(_03202__PTR0), .S(_02422__PTR3), .Z(_02423__PTR8) );
  MUX2_X1 U25291 ( .A(1'b0), .B(_03202__PTR1), .S(_02422__PTR3), .Z(_02423__PTR9) );
  MUX2_X1 U25292 ( .A(1'b0), .B(_03202__PTR2), .S(_02422__PTR3), .Z(_02423__PTR10) );
  MUX2_X1 U25293 ( .A(1'b0), .B(_03202__PTR3), .S(_02422__PTR3), .Z(_02423__PTR11) );
  MUX2_X1 U25294 ( .A(1'b0), .B(_03202__PTR4), .S(_02422__PTR3), .Z(_02423__PTR12) );
  MUX2_X1 U25295 ( .A(1'b0), .B(_03202__PTR5), .S(_02422__PTR3), .Z(_02423__PTR13) );
  MUX2_X1 U25296 ( .A(1'b0), .B(_03202__PTR6), .S(_02422__PTR3), .Z(_02423__PTR14) );
  MUX2_X1 U25297 ( .A(1'b0), .B(_03202__PTR7), .S(_02422__PTR3), .Z(_02423__PTR15) );
  MUX2_X1 U25298 ( .A(_03201__PTR0), .B(1'b0), .S(_02422__PTR2), .Z(_03202__PTR0) );
  MUX2_X1 U25299 ( .A(_03201__PTR1), .B(1'b0), .S(_02422__PTR2), .Z(_03202__PTR1) );
  MUX2_X1 U25300 ( .A(_03201__PTR2), .B(1'b0), .S(_02422__PTR2), .Z(_03202__PTR2) );
  MUX2_X1 U25301 ( .A(_03201__PTR3), .B(1'b0), .S(_02422__PTR2), .Z(_03202__PTR3) );
  MUX2_X1 U25302 ( .A(1'b0), .B(_03201__PTR0), .S(_02422__PTR2), .Z(_03202__PTR4) );
  MUX2_X1 U25303 ( .A(1'b0), .B(_03201__PTR1), .S(_02422__PTR2), .Z(_03202__PTR5) );
  MUX2_X1 U25304 ( .A(1'b0), .B(_03201__PTR2), .S(_02422__PTR2), .Z(_03202__PTR6) );
  MUX2_X1 U25305 ( .A(1'b0), .B(_03201__PTR3), .S(_02422__PTR2), .Z(_03202__PTR7) );
  MUX2_X1 U25306 ( .A(P3_P1_InstQueueWr_Addr_PTR0), .B(1'b0), .S(_02422__PTR1), .Z(_03201__PTR0) );
  MUX2_X1 U25307 ( .A(_02418__PTR0), .B(1'b0), .S(_02422__PTR1), .Z(_03201__PTR1) );
  MUX2_X1 U25308 ( .A(1'b0), .B(P3_P1_InstQueueWr_Addr_PTR0), .S(_02422__PTR1), .Z(_03201__PTR2) );
  MUX2_X1 U25309 ( .A(1'b0), .B(_02418__PTR0), .S(_02422__PTR1), .Z(_03201__PTR3) );
  MUX2_X1 U25310 ( .A(_03245__PTR0), .B(_03245__PTR4), .S(P3_State_PTR2), .Z(_02425_) );
  MUX2_X1 U25311 ( .A(_03244__PTR0), .B(_03244__PTR6), .S(P3_State_PTR1), .Z(_03245__PTR0) );
  MUX2_X1 U25312 ( .A(1'b0), .B(_03244__PTR6), .S(P3_State_PTR1), .Z(_03245__PTR4) );
  MUX2_X1 U25313 ( .A(1'b1), .B(1'b0), .S(P3_State_PTR0), .Z(_03244__PTR0) );
  MUX2_X1 U25314 ( .A(_02424__PTR6), .B(P3_D_C_n), .S(P3_State_PTR0), .Z(_03244__PTR6) );
  MUX2_X1 U25315 ( .A(_03247__PTR0), .B(_03247__PTR4), .S(P3_State_PTR2), .Z(_02426_) );
  MUX2_X1 U25316 ( .A(_03246__PTR4), .B(P3_State_PTR0), .S(P3_State_PTR1), .Z(_03247__PTR0) );
  MUX2_X1 U25317 ( .A(_03246__PTR4), .B(_03246__PTR6), .S(P3_State_PTR1), .Z(_03247__PTR4) );
  MUX2_X1 U25318 ( .A(1'b1), .B(P3_ADS_n), .S(P3_State_PTR0), .Z(_03246__PTR4) );
  MUX2_X1 U25319 ( .A(1'b0), .B(1'b0), .S(P3_State_PTR0), .Z(_03246__PTR6) );
  MUX2_X1 U25320 ( .A(_03249__PTR0), .B(_03249__PTR4), .S(P3_State_PTR2), .Z(_02427_) );
  MUX2_X1 U25321 ( .A(_03244__PTR0), .B(_03248__PTR2), .S(P3_State_PTR1), .Z(_03249__PTR0) );
  MUX2_X1 U25322 ( .A(_03248__PTR4), .B(1'b0), .S(P3_State_PTR1), .Z(_03249__PTR4) );
  MUX2_X1 U25323 ( .A(1'b0), .B(bs16), .S(P3_State_PTR0), .Z(_03248__PTR2) );
  MUX2_X1 U25324 ( .A(bs16), .B(1'b0), .S(P3_State_PTR0), .Z(_03248__PTR4) );
  MUX2_X1 U25325 ( .A(_03251__PTR0), .B(_03251__PTR4), .S(P3_P1_State2_PTR2), .Z(_03252__PTR0) );
  MUX2_X1 U25326 ( .A(1'b1), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03251__PTR0) );
  MUX2_X1 U25327 ( .A(_03250__PTR4), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03251__PTR4) );
  MUX2_X1 U25328 ( .A(1'b0), .B(_02429__PTR5), .S(P3_P1_State2_PTR0), .Z(_03250__PTR4) );
  MUX2_X1 U25329 ( .A(_03251__PTR0), .B(_03254__PTR4), .S(P3_P1_State2_PTR2), .Z(_03255__PTR0) );
  MUX2_X1 U25330 ( .A(_03253__PTR4), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03254__PTR4) );
  MUX2_X1 U25331 ( .A(1'b0), .B(_02430__PTR5), .S(P3_P1_State2_PTR0), .Z(_03253__PTR4) );
  MUX2_X1 U25332 ( .A(_03257__PTR0), .B(_03257__PTR4), .S(P3_P1_State2_PTR2), .Z(_03258__PTR0) );
  MUX2_X1 U25333 ( .A(1'b1), .B(P3_P1_State2_PTR0), .S(P3_P1_State2_PTR1), .Z(_03257__PTR0) );
  MUX2_X1 U25334 ( .A(_03256__PTR4), .B(_03256__PTR6), .S(P3_P1_State2_PTR1), .Z(_03257__PTR4) );
  MUX2_X1 U25335 ( .A(1'b0), .B(_02431__PTR5), .S(P3_P1_State2_PTR0), .Z(_03256__PTR4) );
  MUX2_X1 U25336 ( .A(_02431__PTR6), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03256__PTR6) );
  MUX2_X1 U25337 ( .A(_03260__PTR0), .B(_03260__PTR4), .S(P3_P1_State2_PTR2), .Z(_03261__PTR0) );
  MUX2_X1 U25338 ( .A(_03259__PTR0), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03260__PTR0) );
  MUX2_X1 U25339 ( .A(_03259__PTR4), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03260__PTR4) );
  MUX2_X1 U25340 ( .A(1'b0), .B(1'b1), .S(P3_P1_State2_PTR0), .Z(_03259__PTR0) );
  MUX2_X1 U25341 ( .A(1'b0), .B(_02432__PTR5), .S(P3_P1_State2_PTR0), .Z(_03259__PTR4) );
  MUX2_X1 U25342 ( .A(_03322__PTR0), .B(_03322__PTR16), .S(P3_State_PTR2), .Z(_02459__PTR0) );
  MUX2_X1 U25343 ( .A(_03322__PTR1), .B(_03322__PTR17), .S(P3_State_PTR2), .Z(_02459__PTR1) );
  MUX2_X1 U25344 ( .A(_03322__PTR2), .B(_03322__PTR18), .S(P3_State_PTR2), .Z(_02459__PTR2) );
  MUX2_X1 U25345 ( .A(_03324__PTR0), .B(_03323__PTR0), .S(P3_State_PTR1), .Z(_03322__PTR0) );
  MUX2_X1 U25346 ( .A(_03324__PTR1), .B(_03323__PTR1), .S(P3_State_PTR1), .Z(_03322__PTR1) );
  MUX2_X1 U25347 ( .A(_03324__PTR2), .B(_03323__PTR2), .S(P3_State_PTR1), .Z(_03322__PTR2) );
  MUX2_X1 U25348 ( .A(_03323__PTR8), .B(_03323__PTR16), .S(P3_State_PTR1), .Z(_03322__PTR16) );
  MUX2_X1 U25349 ( .A(_03323__PTR9), .B(_03323__PTR17), .S(P3_State_PTR1), .Z(_03322__PTR17) );
  MUX2_X1 U25350 ( .A(_03323__PTR10), .B(_03323__PTR18), .S(P3_State_PTR1), .Z(_03322__PTR18) );
  MUX2_X1 U25351 ( .A(1'b1), .B(_02458__PTR4), .S(P3_State_PTR0), .Z(_03324__PTR0) );
  MUX2_X1 U25352 ( .A(1'b0), .B(P3_RequestPending), .S(P3_State_PTR0), .Z(_03324__PTR1) );
  MUX2_X1 U25353 ( .A(1'b0), .B(_02458__PTR6), .S(P3_State_PTR0), .Z(_03324__PTR2) );
  MUX2_X1 U25354 ( .A(1'b1), .B(_02458__PTR12), .S(P3_State_PTR0), .Z(_03323__PTR0) );
  MUX2_X1 U25355 ( .A(1'b1), .B(_02458__PTR13), .S(P3_State_PTR0), .Z(_03323__PTR1) );
  MUX2_X1 U25356 ( .A(1'b0), .B(_02458__PTR14), .S(P3_State_PTR0), .Z(_03323__PTR2) );
  MUX2_X1 U25357 ( .A(_02458__PTR16), .B(_02458__PTR20), .S(P3_State_PTR0), .Z(_03323__PTR8) );
  MUX2_X1 U25358 ( .A(_02458__PTR17), .B(_02458__PTR21), .S(P3_State_PTR0), .Z(_03323__PTR9) );
  MUX2_X1 U25359 ( .A(_02458__PTR18), .B(_02458__PTR22), .S(P3_State_PTR0), .Z(_03323__PTR10) );
  MUX2_X1 U25360 ( .A(1'b0), .B(_02458__PTR28), .S(P3_State_PTR0), .Z(_03323__PTR16) );
  MUX2_X1 U25361 ( .A(P3_READY_n), .B(_02458__PTR29), .S(P3_State_PTR0), .Z(_03323__PTR17) );
  MUX2_X1 U25362 ( .A(1'b1), .B(_02458__PTR30), .S(P3_State_PTR0), .Z(_03323__PTR18) );
  MUX2_X1 U25363 ( .A(_03326__PTR0), .B(_03326__PTR256), .S(P3_State_PTR2), .Z(_02460__PTR0) );
  MUX2_X1 U25364 ( .A(_03326__PTR2), .B(_03326__PTR258), .S(P3_State_PTR2), .Z(_02460__PTR2) );
  MUX2_X1 U25365 ( .A(_03326__PTR3), .B(_03326__PTR259), .S(P3_State_PTR2), .Z(_02460__PTR3) );
  MUX2_X1 U25366 ( .A(_03326__PTR4), .B(_03326__PTR260), .S(P3_State_PTR2), .Z(_02460__PTR4) );
  MUX2_X1 U25367 ( .A(_03326__PTR5), .B(_03326__PTR261), .S(P3_State_PTR2), .Z(_02460__PTR5) );
  MUX2_X1 U25368 ( .A(_03326__PTR6), .B(_03326__PTR262), .S(P3_State_PTR2), .Z(_02460__PTR6) );
  MUX2_X1 U25369 ( .A(_03326__PTR7), .B(_03326__PTR263), .S(P3_State_PTR2), .Z(_02460__PTR7) );
  MUX2_X1 U25370 ( .A(_03326__PTR8), .B(_03326__PTR264), .S(P3_State_PTR2), .Z(_02460__PTR8) );
  MUX2_X1 U25371 ( .A(_03326__PTR9), .B(_03326__PTR265), .S(P3_State_PTR2), .Z(_02460__PTR9) );
  MUX2_X1 U25372 ( .A(_03326__PTR10), .B(_03326__PTR266), .S(P3_State_PTR2), .Z(_02460__PTR10) );
  MUX2_X1 U25373 ( .A(_03326__PTR11), .B(_03326__PTR267), .S(P3_State_PTR2), .Z(_02460__PTR11) );
  MUX2_X1 U25374 ( .A(_03326__PTR12), .B(_03326__PTR268), .S(P3_State_PTR2), .Z(_02460__PTR12) );
  MUX2_X1 U25375 ( .A(_03326__PTR13), .B(_03326__PTR269), .S(P3_State_PTR2), .Z(_02460__PTR13) );
  MUX2_X1 U25376 ( .A(_03326__PTR14), .B(_03326__PTR270), .S(P3_State_PTR2), .Z(_02460__PTR14) );
  MUX2_X1 U25377 ( .A(_03326__PTR15), .B(_03326__PTR271), .S(P3_State_PTR2), .Z(_02460__PTR15) );
  MUX2_X1 U25378 ( .A(_03326__PTR16), .B(_03326__PTR272), .S(P3_State_PTR2), .Z(_02460__PTR16) );
  MUX2_X1 U25379 ( .A(_03326__PTR17), .B(_03326__PTR273), .S(P3_State_PTR2), .Z(_02460__PTR17) );
  MUX2_X1 U25380 ( .A(_03326__PTR18), .B(_03326__PTR274), .S(P3_State_PTR2), .Z(_02460__PTR18) );
  MUX2_X1 U25381 ( .A(_03326__PTR19), .B(_03326__PTR275), .S(P3_State_PTR2), .Z(_02460__PTR19) );
  MUX2_X1 U25382 ( .A(_03326__PTR20), .B(_03326__PTR276), .S(P3_State_PTR2), .Z(_02460__PTR20) );
  MUX2_X1 U25383 ( .A(_03326__PTR21), .B(_03326__PTR277), .S(P3_State_PTR2), .Z(_02460__PTR21) );
  MUX2_X1 U25384 ( .A(_03326__PTR22), .B(_03326__PTR278), .S(P3_State_PTR2), .Z(_02460__PTR22) );
  MUX2_X1 U25385 ( .A(_03326__PTR23), .B(_03326__PTR279), .S(P3_State_PTR2), .Z(_02460__PTR23) );
  MUX2_X1 U25386 ( .A(_03326__PTR24), .B(_03326__PTR280), .S(P3_State_PTR2), .Z(_02460__PTR24) );
  MUX2_X1 U25387 ( .A(_03326__PTR25), .B(_03326__PTR281), .S(P3_State_PTR2), .Z(_02460__PTR25) );
  MUX2_X1 U25388 ( .A(_03326__PTR26), .B(_03326__PTR282), .S(P3_State_PTR2), .Z(_02460__PTR26) );
  MUX2_X1 U25389 ( .A(_03326__PTR27), .B(_03326__PTR283), .S(P3_State_PTR2), .Z(_02460__PTR27) );
  MUX2_X1 U25390 ( .A(_03326__PTR28), .B(_03326__PTR284), .S(P3_State_PTR2), .Z(_02460__PTR28) );
  MUX2_X1 U25391 ( .A(_03326__PTR29), .B(_03326__PTR285), .S(P3_State_PTR2), .Z(_02460__PTR29) );
  MUX2_X1 U25392 ( .A(_03326__PTR30), .B(_03326__PTR286), .S(P3_State_PTR2), .Z(_02460__PTR30) );
  MUX2_X1 U25393 ( .A(_03326__PTR32), .B(_03326__PTR288), .S(P3_State_PTR2), .Z(_02460__PTR32) );
  MUX2_X1 U25394 ( .A(_03246__PTR6), .B(_03325__PTR128), .S(P3_State_PTR1), .Z(_03326__PTR0) );
  MUX2_X1 U25395 ( .A(_03325__PTR258), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR2) );
  MUX2_X1 U25396 ( .A(_03325__PTR259), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR3) );
  MUX2_X1 U25397 ( .A(_03325__PTR260), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR4) );
  MUX2_X1 U25398 ( .A(_03325__PTR261), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR5) );
  MUX2_X1 U25399 ( .A(_03325__PTR262), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR6) );
  MUX2_X1 U25400 ( .A(_03325__PTR263), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR7) );
  MUX2_X1 U25401 ( .A(_03325__PTR264), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR8) );
  MUX2_X1 U25402 ( .A(_03325__PTR265), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR9) );
  MUX2_X1 U25403 ( .A(_03325__PTR266), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR10) );
  MUX2_X1 U25404 ( .A(_03325__PTR267), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR11) );
  MUX2_X1 U25405 ( .A(_03325__PTR268), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR12) );
  MUX2_X1 U25406 ( .A(_03325__PTR269), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR13) );
  MUX2_X1 U25407 ( .A(_03325__PTR270), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR14) );
  MUX2_X1 U25408 ( .A(_03325__PTR271), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR15) );
  MUX2_X1 U25409 ( .A(_03325__PTR272), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR16) );
  MUX2_X1 U25410 ( .A(_03325__PTR273), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR17) );
  MUX2_X1 U25411 ( .A(_03325__PTR274), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR18) );
  MUX2_X1 U25412 ( .A(_03325__PTR275), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR19) );
  MUX2_X1 U25413 ( .A(_03325__PTR276), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR20) );
  MUX2_X1 U25414 ( .A(_03325__PTR277), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR21) );
  MUX2_X1 U25415 ( .A(_03325__PTR278), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR22) );
  MUX2_X1 U25416 ( .A(_03325__PTR279), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR23) );
  MUX2_X1 U25417 ( .A(_03325__PTR280), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR24) );
  MUX2_X1 U25418 ( .A(_03325__PTR281), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR25) );
  MUX2_X1 U25419 ( .A(_03325__PTR282), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR26) );
  MUX2_X1 U25420 ( .A(_03325__PTR283), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR27) );
  MUX2_X1 U25421 ( .A(_03325__PTR284), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR28) );
  MUX2_X1 U25422 ( .A(_03325__PTR285), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR29) );
  MUX2_X1 U25423 ( .A(_03325__PTR286), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR30) );
  MUX2_X1 U25424 ( .A(_03325__PTR288), .B(_03325__PTR160), .S(P3_State_PTR1), .Z(_03326__PTR32) );
  MUX2_X1 U25425 ( .A(_03325__PTR256), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR256) );
  MUX2_X1 U25426 ( .A(_03325__PTR258), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR258) );
  MUX2_X1 U25427 ( .A(_03325__PTR259), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR259) );
  MUX2_X1 U25428 ( .A(_03325__PTR260), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR260) );
  MUX2_X1 U25429 ( .A(_03325__PTR261), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR261) );
  MUX2_X1 U25430 ( .A(_03325__PTR262), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR262) );
  MUX2_X1 U25431 ( .A(_03325__PTR263), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR263) );
  MUX2_X1 U25432 ( .A(_03325__PTR264), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR264) );
  MUX2_X1 U25433 ( .A(_03325__PTR265), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR265) );
  MUX2_X1 U25434 ( .A(_03325__PTR266), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR266) );
  MUX2_X1 U25435 ( .A(_03325__PTR267), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR267) );
  MUX2_X1 U25436 ( .A(_03325__PTR268), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR268) );
  MUX2_X1 U25437 ( .A(_03325__PTR269), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR269) );
  MUX2_X1 U25438 ( .A(_03325__PTR270), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR270) );
  MUX2_X1 U25439 ( .A(_03325__PTR271), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR271) );
  MUX2_X1 U25440 ( .A(_03325__PTR272), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR272) );
  MUX2_X1 U25441 ( .A(_03325__PTR273), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR273) );
  MUX2_X1 U25442 ( .A(_03325__PTR274), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR274) );
  MUX2_X1 U25443 ( .A(_03325__PTR275), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR275) );
  MUX2_X1 U25444 ( .A(_03325__PTR276), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR276) );
  MUX2_X1 U25445 ( .A(_03325__PTR277), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR277) );
  MUX2_X1 U25446 ( .A(_03325__PTR278), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR278) );
  MUX2_X1 U25447 ( .A(_03325__PTR279), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR279) );
  MUX2_X1 U25448 ( .A(_03325__PTR280), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR280) );
  MUX2_X1 U25449 ( .A(_03325__PTR281), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR281) );
  MUX2_X1 U25450 ( .A(_03325__PTR282), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR282) );
  MUX2_X1 U25451 ( .A(_03325__PTR283), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR283) );
  MUX2_X1 U25452 ( .A(_03325__PTR284), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR284) );
  MUX2_X1 U25453 ( .A(_03325__PTR285), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR285) );
  MUX2_X1 U25454 ( .A(_03325__PTR286), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR286) );
  MUX2_X1 U25455 ( .A(_03325__PTR288), .B(1'b0), .S(P3_State_PTR1), .Z(_03326__PTR288) );
  MUX2_X1 U25456 ( .A(1'b0), .B(_01878__PTR256), .S(P3_State_PTR0), .Z(_03325__PTR128) );
  MUX2_X1 U25457 ( .A(1'b0), .B(1'b0), .S(P3_State_PTR0), .Z(_03325__PTR160) );
  MUX2_X1 U25458 ( .A(_01878__PTR256), .B(1'b0), .S(P3_State_PTR0), .Z(_03325__PTR256) );
  MUX2_X1 U25459 ( .A(1'b0), .B(P3_DataWidth_PTR2), .S(P3_State_PTR0), .Z(_03325__PTR258) );
  MUX2_X1 U25460 ( .A(1'b0), .B(P3_DataWidth_PTR3), .S(P3_State_PTR0), .Z(_03325__PTR259) );
  MUX2_X1 U25461 ( .A(1'b0), .B(P3_DataWidth_PTR4), .S(P3_State_PTR0), .Z(_03325__PTR260) );
  MUX2_X1 U25462 ( .A(1'b0), .B(P3_DataWidth_PTR5), .S(P3_State_PTR0), .Z(_03325__PTR261) );
  MUX2_X1 U25463 ( .A(1'b0), .B(P3_DataWidth_PTR6), .S(P3_State_PTR0), .Z(_03325__PTR262) );
  MUX2_X1 U25464 ( .A(1'b0), .B(P3_DataWidth_PTR7), .S(P3_State_PTR0), .Z(_03325__PTR263) );
  MUX2_X1 U25465 ( .A(1'b0), .B(P3_DataWidth_PTR8), .S(P3_State_PTR0), .Z(_03325__PTR264) );
  MUX2_X1 U25466 ( .A(1'b0), .B(P3_DataWidth_PTR9), .S(P3_State_PTR0), .Z(_03325__PTR265) );
  MUX2_X1 U25467 ( .A(1'b0), .B(P3_DataWidth_PTR10), .S(P3_State_PTR0), .Z(_03325__PTR266) );
  MUX2_X1 U25468 ( .A(1'b0), .B(P3_DataWidth_PTR11), .S(P3_State_PTR0), .Z(_03325__PTR267) );
  MUX2_X1 U25469 ( .A(1'b0), .B(P3_DataWidth_PTR12), .S(P3_State_PTR0), .Z(_03325__PTR268) );
  MUX2_X1 U25470 ( .A(1'b0), .B(P3_DataWidth_PTR13), .S(P3_State_PTR0), .Z(_03325__PTR269) );
  MUX2_X1 U25471 ( .A(1'b0), .B(P3_DataWidth_PTR14), .S(P3_State_PTR0), .Z(_03325__PTR270) );
  MUX2_X1 U25472 ( .A(1'b0), .B(P3_DataWidth_PTR15), .S(P3_State_PTR0), .Z(_03325__PTR271) );
  MUX2_X1 U25473 ( .A(1'b0), .B(P3_DataWidth_PTR16), .S(P3_State_PTR0), .Z(_03325__PTR272) );
  MUX2_X1 U25474 ( .A(1'b0), .B(P3_DataWidth_PTR17), .S(P3_State_PTR0), .Z(_03325__PTR273) );
  MUX2_X1 U25475 ( .A(1'b0), .B(P3_DataWidth_PTR18), .S(P3_State_PTR0), .Z(_03325__PTR274) );
  MUX2_X1 U25476 ( .A(1'b0), .B(P3_DataWidth_PTR19), .S(P3_State_PTR0), .Z(_03325__PTR275) );
  MUX2_X1 U25477 ( .A(1'b0), .B(P3_DataWidth_PTR20), .S(P3_State_PTR0), .Z(_03325__PTR276) );
  MUX2_X1 U25478 ( .A(1'b0), .B(P3_DataWidth_PTR21), .S(P3_State_PTR0), .Z(_03325__PTR277) );
  MUX2_X1 U25479 ( .A(1'b0), .B(P3_DataWidth_PTR22), .S(P3_State_PTR0), .Z(_03325__PTR278) );
  MUX2_X1 U25480 ( .A(1'b0), .B(P3_DataWidth_PTR23), .S(P3_State_PTR0), .Z(_03325__PTR279) );
  MUX2_X1 U25481 ( .A(1'b0), .B(P3_DataWidth_PTR24), .S(P3_State_PTR0), .Z(_03325__PTR280) );
  MUX2_X1 U25482 ( .A(1'b0), .B(P3_DataWidth_PTR25), .S(P3_State_PTR0), .Z(_03325__PTR281) );
  MUX2_X1 U25483 ( .A(1'b0), .B(P3_DataWidth_PTR26), .S(P3_State_PTR0), .Z(_03325__PTR282) );
  MUX2_X1 U25484 ( .A(1'b0), .B(P3_DataWidth_PTR27), .S(P3_State_PTR0), .Z(_03325__PTR283) );
  MUX2_X1 U25485 ( .A(1'b0), .B(P3_DataWidth_PTR28), .S(P3_State_PTR0), .Z(_03325__PTR284) );
  MUX2_X1 U25486 ( .A(1'b0), .B(P3_DataWidth_PTR29), .S(P3_State_PTR0), .Z(_03325__PTR285) );
  MUX2_X1 U25487 ( .A(1'b0), .B(P3_DataWidth_PTR30), .S(P3_State_PTR0), .Z(_03325__PTR286) );
  MUX2_X1 U25488 ( .A(1'b0), .B(P3_DataWidth_PTR31), .S(P3_State_PTR0), .Z(_03325__PTR288) );
  MUX2_X1 U25489 ( .A(_03328__PTR0), .B(_03328__PTR128), .S(P3_State_PTR2), .Z(_02462__PTR0) );
  MUX2_X1 U25490 ( .A(_03328__PTR1), .B(_03328__PTR129), .S(P3_State_PTR2), .Z(_02462__PTR1) );
  MUX2_X1 U25491 ( .A(_03328__PTR2), .B(_03328__PTR130), .S(P3_State_PTR2), .Z(_02462__PTR2) );
  MUX2_X1 U25492 ( .A(_03328__PTR3), .B(_03328__PTR131), .S(P3_State_PTR2), .Z(_02462__PTR3) );
  MUX2_X1 U25493 ( .A(_03328__PTR4), .B(_03328__PTR132), .S(P3_State_PTR2), .Z(_02462__PTR4) );
  MUX2_X1 U25494 ( .A(_03328__PTR5), .B(_03328__PTR133), .S(P3_State_PTR2), .Z(_02462__PTR5) );
  MUX2_X1 U25495 ( .A(_03328__PTR6), .B(_03328__PTR134), .S(P3_State_PTR2), .Z(_02462__PTR6) );
  MUX2_X1 U25496 ( .A(_03328__PTR7), .B(_03328__PTR135), .S(P3_State_PTR2), .Z(_02462__PTR7) );
  MUX2_X1 U25497 ( .A(_03328__PTR8), .B(_03328__PTR136), .S(P3_State_PTR2), .Z(_02462__PTR8) );
  MUX2_X1 U25498 ( .A(_03328__PTR9), .B(_03328__PTR137), .S(P3_State_PTR2), .Z(_02462__PTR9) );
  MUX2_X1 U25499 ( .A(_03328__PTR10), .B(_03328__PTR138), .S(P3_State_PTR2), .Z(_02462__PTR10) );
  MUX2_X1 U25500 ( .A(_03328__PTR11), .B(_03328__PTR139), .S(P3_State_PTR2), .Z(_02462__PTR11) );
  MUX2_X1 U25501 ( .A(_03328__PTR12), .B(_03328__PTR140), .S(P3_State_PTR2), .Z(_02462__PTR12) );
  MUX2_X1 U25502 ( .A(_03328__PTR13), .B(_03328__PTR141), .S(P3_State_PTR2), .Z(_02462__PTR13) );
  MUX2_X1 U25503 ( .A(_03328__PTR14), .B(_03328__PTR142), .S(P3_State_PTR2), .Z(_02462__PTR14) );
  MUX2_X1 U25504 ( .A(_03328__PTR15), .B(_03328__PTR143), .S(P3_State_PTR2), .Z(_02462__PTR15) );
  MUX2_X1 U25505 ( .A(_03328__PTR16), .B(_03328__PTR144), .S(P3_State_PTR2), .Z(_02462__PTR16) );
  MUX2_X1 U25506 ( .A(_03328__PTR17), .B(_03328__PTR145), .S(P3_State_PTR2), .Z(_02462__PTR17) );
  MUX2_X1 U25507 ( .A(_03328__PTR18), .B(_03328__PTR146), .S(P3_State_PTR2), .Z(_02462__PTR18) );
  MUX2_X1 U25508 ( .A(_03328__PTR19), .B(_03328__PTR147), .S(P3_State_PTR2), .Z(_02462__PTR19) );
  MUX2_X1 U25509 ( .A(_03328__PTR20), .B(_03328__PTR148), .S(P3_State_PTR2), .Z(_02462__PTR20) );
  MUX2_X1 U25510 ( .A(_03328__PTR21), .B(_03328__PTR149), .S(P3_State_PTR2), .Z(_02462__PTR21) );
  MUX2_X1 U25511 ( .A(_03328__PTR22), .B(_03328__PTR150), .S(P3_State_PTR2), .Z(_02462__PTR22) );
  MUX2_X1 U25512 ( .A(_03328__PTR23), .B(_03328__PTR151), .S(P3_State_PTR2), .Z(_02462__PTR23) );
  MUX2_X1 U25513 ( .A(_03328__PTR24), .B(_03328__PTR152), .S(P3_State_PTR2), .Z(_02462__PTR24) );
  MUX2_X1 U25514 ( .A(_03328__PTR25), .B(_03328__PTR153), .S(P3_State_PTR2), .Z(_02462__PTR25) );
  MUX2_X1 U25515 ( .A(_03328__PTR26), .B(_03328__PTR154), .S(P3_State_PTR2), .Z(_02462__PTR26) );
  MUX2_X1 U25516 ( .A(_03328__PTR27), .B(_03328__PTR155), .S(P3_State_PTR2), .Z(_02462__PTR27) );
  MUX2_X1 U25517 ( .A(_03328__PTR28), .B(_03328__PTR156), .S(P3_State_PTR2), .Z(_02462__PTR28) );
  MUX2_X1 U25518 ( .A(_03328__PTR29), .B(_03328__PTR157), .S(P3_State_PTR2), .Z(_02462__PTR29) );
  MUX2_X1 U25519 ( .A(1'b0), .B(_03327__PTR64), .S(P3_State_PTR1), .Z(_03328__PTR0) );
  MUX2_X1 U25520 ( .A(1'b0), .B(_03327__PTR65), .S(P3_State_PTR1), .Z(_03328__PTR1) );
  MUX2_X1 U25521 ( .A(1'b0), .B(_03327__PTR66), .S(P3_State_PTR1), .Z(_03328__PTR2) );
  MUX2_X1 U25522 ( .A(1'b0), .B(_03327__PTR67), .S(P3_State_PTR1), .Z(_03328__PTR3) );
  MUX2_X1 U25523 ( .A(1'b0), .B(_03327__PTR68), .S(P3_State_PTR1), .Z(_03328__PTR4) );
  MUX2_X1 U25524 ( .A(1'b0), .B(_03327__PTR69), .S(P3_State_PTR1), .Z(_03328__PTR5) );
  MUX2_X1 U25525 ( .A(1'b0), .B(_03327__PTR70), .S(P3_State_PTR1), .Z(_03328__PTR6) );
  MUX2_X1 U25526 ( .A(1'b0), .B(_03327__PTR71), .S(P3_State_PTR1), .Z(_03328__PTR7) );
  MUX2_X1 U25527 ( .A(1'b0), .B(_03327__PTR72), .S(P3_State_PTR1), .Z(_03328__PTR8) );
  MUX2_X1 U25528 ( .A(1'b0), .B(_03327__PTR73), .S(P3_State_PTR1), .Z(_03328__PTR9) );
  MUX2_X1 U25529 ( .A(1'b0), .B(_03327__PTR74), .S(P3_State_PTR1), .Z(_03328__PTR10) );
  MUX2_X1 U25530 ( .A(1'b0), .B(_03327__PTR75), .S(P3_State_PTR1), .Z(_03328__PTR11) );
  MUX2_X1 U25531 ( .A(1'b0), .B(_03327__PTR76), .S(P3_State_PTR1), .Z(_03328__PTR12) );
  MUX2_X1 U25532 ( .A(1'b0), .B(_03327__PTR77), .S(P3_State_PTR1), .Z(_03328__PTR13) );
  MUX2_X1 U25533 ( .A(1'b0), .B(_03327__PTR78), .S(P3_State_PTR1), .Z(_03328__PTR14) );
  MUX2_X1 U25534 ( .A(1'b0), .B(_03327__PTR79), .S(P3_State_PTR1), .Z(_03328__PTR15) );
  MUX2_X1 U25535 ( .A(1'b0), .B(_03327__PTR80), .S(P3_State_PTR1), .Z(_03328__PTR16) );
  MUX2_X1 U25536 ( .A(1'b0), .B(_03327__PTR81), .S(P3_State_PTR1), .Z(_03328__PTR17) );
  MUX2_X1 U25537 ( .A(1'b0), .B(_03327__PTR82), .S(P3_State_PTR1), .Z(_03328__PTR18) );
  MUX2_X1 U25538 ( .A(1'b0), .B(_03327__PTR83), .S(P3_State_PTR1), .Z(_03328__PTR19) );
  MUX2_X1 U25539 ( .A(1'b0), .B(_03327__PTR84), .S(P3_State_PTR1), .Z(_03328__PTR20) );
  MUX2_X1 U25540 ( .A(1'b0), .B(_03327__PTR85), .S(P3_State_PTR1), .Z(_03328__PTR21) );
  MUX2_X1 U25541 ( .A(1'b0), .B(_03327__PTR86), .S(P3_State_PTR1), .Z(_03328__PTR22) );
  MUX2_X1 U25542 ( .A(1'b0), .B(_03327__PTR87), .S(P3_State_PTR1), .Z(_03328__PTR23) );
  MUX2_X1 U25543 ( .A(1'b0), .B(_03327__PTR88), .S(P3_State_PTR1), .Z(_03328__PTR24) );
  MUX2_X1 U25544 ( .A(1'b0), .B(_03327__PTR89), .S(P3_State_PTR1), .Z(_03328__PTR25) );
  MUX2_X1 U25545 ( .A(1'b0), .B(_03327__PTR90), .S(P3_State_PTR1), .Z(_03328__PTR26) );
  MUX2_X1 U25546 ( .A(1'b0), .B(_03327__PTR91), .S(P3_State_PTR1), .Z(_03328__PTR27) );
  MUX2_X1 U25547 ( .A(1'b0), .B(_03327__PTR92), .S(P3_State_PTR1), .Z(_03328__PTR28) );
  MUX2_X1 U25548 ( .A(1'b0), .B(_03327__PTR93), .S(P3_State_PTR1), .Z(_03328__PTR29) );
  MUX2_X1 U25549 ( .A(1'b0), .B(_03327__PTR192), .S(P3_State_PTR1), .Z(_03328__PTR128) );
  MUX2_X1 U25550 ( .A(1'b0), .B(_03327__PTR193), .S(P3_State_PTR1), .Z(_03328__PTR129) );
  MUX2_X1 U25551 ( .A(1'b0), .B(_03327__PTR194), .S(P3_State_PTR1), .Z(_03328__PTR130) );
  MUX2_X1 U25552 ( .A(1'b0), .B(_03327__PTR195), .S(P3_State_PTR1), .Z(_03328__PTR131) );
  MUX2_X1 U25553 ( .A(1'b0), .B(_03327__PTR196), .S(P3_State_PTR1), .Z(_03328__PTR132) );
  MUX2_X1 U25554 ( .A(1'b0), .B(_03327__PTR197), .S(P3_State_PTR1), .Z(_03328__PTR133) );
  MUX2_X1 U25555 ( .A(1'b0), .B(_03327__PTR198), .S(P3_State_PTR1), .Z(_03328__PTR134) );
  MUX2_X1 U25556 ( .A(1'b0), .B(_03327__PTR199), .S(P3_State_PTR1), .Z(_03328__PTR135) );
  MUX2_X1 U25557 ( .A(1'b0), .B(_03327__PTR200), .S(P3_State_PTR1), .Z(_03328__PTR136) );
  MUX2_X1 U25558 ( .A(1'b0), .B(_03327__PTR201), .S(P3_State_PTR1), .Z(_03328__PTR137) );
  MUX2_X1 U25559 ( .A(1'b0), .B(_03327__PTR202), .S(P3_State_PTR1), .Z(_03328__PTR138) );
  MUX2_X1 U25560 ( .A(1'b0), .B(_03327__PTR203), .S(P3_State_PTR1), .Z(_03328__PTR139) );
  MUX2_X1 U25561 ( .A(1'b0), .B(_03327__PTR204), .S(P3_State_PTR1), .Z(_03328__PTR140) );
  MUX2_X1 U25562 ( .A(1'b0), .B(_03327__PTR205), .S(P3_State_PTR1), .Z(_03328__PTR141) );
  MUX2_X1 U25563 ( .A(1'b0), .B(_03327__PTR206), .S(P3_State_PTR1), .Z(_03328__PTR142) );
  MUX2_X1 U25564 ( .A(1'b0), .B(_03327__PTR207), .S(P3_State_PTR1), .Z(_03328__PTR143) );
  MUX2_X1 U25565 ( .A(1'b0), .B(_03327__PTR208), .S(P3_State_PTR1), .Z(_03328__PTR144) );
  MUX2_X1 U25566 ( .A(1'b0), .B(_03327__PTR209), .S(P3_State_PTR1), .Z(_03328__PTR145) );
  MUX2_X1 U25567 ( .A(1'b0), .B(_03327__PTR210), .S(P3_State_PTR1), .Z(_03328__PTR146) );
  MUX2_X1 U25568 ( .A(1'b0), .B(_03327__PTR211), .S(P3_State_PTR1), .Z(_03328__PTR147) );
  MUX2_X1 U25569 ( .A(1'b0), .B(_03327__PTR212), .S(P3_State_PTR1), .Z(_03328__PTR148) );
  MUX2_X1 U25570 ( .A(1'b0), .B(_03327__PTR213), .S(P3_State_PTR1), .Z(_03328__PTR149) );
  MUX2_X1 U25571 ( .A(1'b0), .B(_03327__PTR214), .S(P3_State_PTR1), .Z(_03328__PTR150) );
  MUX2_X1 U25572 ( .A(1'b0), .B(_03327__PTR215), .S(P3_State_PTR1), .Z(_03328__PTR151) );
  MUX2_X1 U25573 ( .A(1'b0), .B(_03327__PTR216), .S(P3_State_PTR1), .Z(_03328__PTR152) );
  MUX2_X1 U25574 ( .A(1'b0), .B(_03327__PTR217), .S(P3_State_PTR1), .Z(_03328__PTR153) );
  MUX2_X1 U25575 ( .A(1'b0), .B(_03327__PTR218), .S(P3_State_PTR1), .Z(_03328__PTR154) );
  MUX2_X1 U25576 ( .A(1'b0), .B(_03327__PTR219), .S(P3_State_PTR1), .Z(_03328__PTR155) );
  MUX2_X1 U25577 ( .A(1'b0), .B(_03327__PTR220), .S(P3_State_PTR1), .Z(_03328__PTR156) );
  MUX2_X1 U25578 ( .A(1'b0), .B(_03327__PTR221), .S(P3_State_PTR1), .Z(_03328__PTR157) );
  MUX2_X1 U25579 ( .A(_02461__PTR64), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR64) );
  MUX2_X1 U25580 ( .A(_02461__PTR65), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR65) );
  MUX2_X1 U25581 ( .A(_02461__PTR66), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR66) );
  MUX2_X1 U25582 ( .A(_02461__PTR67), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR67) );
  MUX2_X1 U25583 ( .A(_02461__PTR68), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR68) );
  MUX2_X1 U25584 ( .A(_02461__PTR69), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR69) );
  MUX2_X1 U25585 ( .A(_02461__PTR70), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR70) );
  MUX2_X1 U25586 ( .A(_02461__PTR71), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR71) );
  MUX2_X1 U25587 ( .A(_02461__PTR72), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR72) );
  MUX2_X1 U25588 ( .A(_02461__PTR73), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR73) );
  MUX2_X1 U25589 ( .A(_02461__PTR74), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR74) );
  MUX2_X1 U25590 ( .A(_02461__PTR75), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR75) );
  MUX2_X1 U25591 ( .A(_02461__PTR76), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR76) );
  MUX2_X1 U25592 ( .A(_02461__PTR77), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR77) );
  MUX2_X1 U25593 ( .A(_02461__PTR78), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR78) );
  MUX2_X1 U25594 ( .A(_02461__PTR79), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR79) );
  MUX2_X1 U25595 ( .A(_02461__PTR80), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR80) );
  MUX2_X1 U25596 ( .A(_02461__PTR81), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR81) );
  MUX2_X1 U25597 ( .A(_02461__PTR82), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR82) );
  MUX2_X1 U25598 ( .A(_02461__PTR83), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR83) );
  MUX2_X1 U25599 ( .A(_02461__PTR84), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR84) );
  MUX2_X1 U25600 ( .A(_02461__PTR85), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR85) );
  MUX2_X1 U25601 ( .A(_02461__PTR86), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR86) );
  MUX2_X1 U25602 ( .A(_02461__PTR87), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR87) );
  MUX2_X1 U25603 ( .A(_02461__PTR88), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR88) );
  MUX2_X1 U25604 ( .A(_02461__PTR89), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR89) );
  MUX2_X1 U25605 ( .A(_02461__PTR90), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR90) );
  MUX2_X1 U25606 ( .A(_02461__PTR91), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR91) );
  MUX2_X1 U25607 ( .A(_02461__PTR92), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR92) );
  MUX2_X1 U25608 ( .A(_02461__PTR93), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR93) );
  MUX2_X1 U25609 ( .A(_02461__PTR192), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR192) );
  MUX2_X1 U25610 ( .A(_02461__PTR193), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR193) );
  MUX2_X1 U25611 ( .A(_02461__PTR194), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR194) );
  MUX2_X1 U25612 ( .A(_02461__PTR195), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR195) );
  MUX2_X1 U25613 ( .A(_02461__PTR196), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR196) );
  MUX2_X1 U25614 ( .A(_02461__PTR197), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR197) );
  MUX2_X1 U25615 ( .A(_02461__PTR198), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR198) );
  MUX2_X1 U25616 ( .A(_02461__PTR199), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR199) );
  MUX2_X1 U25617 ( .A(_02461__PTR200), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR200) );
  MUX2_X1 U25618 ( .A(_02461__PTR201), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR201) );
  MUX2_X1 U25619 ( .A(_02461__PTR202), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR202) );
  MUX2_X1 U25620 ( .A(_02461__PTR203), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR203) );
  MUX2_X1 U25621 ( .A(_02461__PTR204), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR204) );
  MUX2_X1 U25622 ( .A(_02461__PTR205), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR205) );
  MUX2_X1 U25623 ( .A(_02461__PTR206), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR206) );
  MUX2_X1 U25624 ( .A(_02461__PTR207), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR207) );
  MUX2_X1 U25625 ( .A(_02461__PTR208), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR208) );
  MUX2_X1 U25626 ( .A(_02461__PTR209), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR209) );
  MUX2_X1 U25627 ( .A(_02461__PTR210), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR210) );
  MUX2_X1 U25628 ( .A(_02461__PTR211), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR211) );
  MUX2_X1 U25629 ( .A(_02461__PTR212), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR212) );
  MUX2_X1 U25630 ( .A(_02461__PTR213), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR213) );
  MUX2_X1 U25631 ( .A(_02461__PTR214), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR214) );
  MUX2_X1 U25632 ( .A(_02461__PTR215), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR215) );
  MUX2_X1 U25633 ( .A(_02461__PTR216), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR216) );
  MUX2_X1 U25634 ( .A(_02461__PTR217), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR217) );
  MUX2_X1 U25635 ( .A(_02461__PTR218), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR218) );
  MUX2_X1 U25636 ( .A(_02461__PTR219), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR219) );
  MUX2_X1 U25637 ( .A(_02461__PTR220), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR220) );
  MUX2_X1 U25638 ( .A(_02461__PTR221), .B(1'b0), .S(P3_State_PTR0), .Z(_03327__PTR221) );
  INV_X1 U25639 ( .A(P3_rEIP_PTR0), .ZN(_03329__PTR43) );
  MUX2_X1 U25640 ( .A(1'b0), .B(P3_rEIP_PTR0), .S(P3_rEIP_PTR1), .Z(_02463__PTR2) );
  MUX2_X1 U25641 ( .A(_03329__PTR43), .B(P3_rEIP_PTR0), .S(P3_rEIP_PTR1), .Z(_02463__PTR6) );
  MUX2_X1 U25642 ( .A(P3_rEIP_PTR0), .B(1'b1), .S(P3_rEIP_PTR1), .Z(_02463__PTR8) );
  MUX2_X1 U25643 ( .A(_03329__PTR43), .B(1'b1), .S(P3_rEIP_PTR1), .Z(_02463__PTR9) );
  MUX2_X1 U25644 ( .A(1'b1), .B(P3_rEIP_PTR0), .S(P3_rEIP_PTR1), .Z(_02463__PTR10) );
  MUX2_X1 U25645 ( .A(1'b1), .B(_03329__PTR43), .S(P3_rEIP_PTR1), .Z(_02463__PTR11) );
  MUX2_X1 U25646 ( .A(_03332__PTR0), .B(_03332__PTR64), .S(P3_P1_InstQueueRd_Addr_PTR3), .Z(_02464__PTR0) );
  MUX2_X1 U25647 ( .A(_03332__PTR1), .B(_03332__PTR65), .S(P3_P1_InstQueueRd_Addr_PTR3), .Z(_02464__PTR1) );
  MUX2_X1 U25648 ( .A(_03332__PTR2), .B(_03332__PTR66), .S(P3_P1_InstQueueRd_Addr_PTR3), .Z(_02464__PTR2) );
  MUX2_X1 U25649 ( .A(_03332__PTR3), .B(_03332__PTR67), .S(P3_P1_InstQueueRd_Addr_PTR3), .Z(_02464__PTR3) );
  MUX2_X1 U25650 ( .A(_03332__PTR4), .B(_03332__PTR68), .S(P3_P1_InstQueueRd_Addr_PTR3), .Z(_02464__PTR4) );
  MUX2_X1 U25651 ( .A(_03332__PTR5), .B(_03332__PTR69), .S(P3_P1_InstQueueRd_Addr_PTR3), .Z(_02464__PTR5) );
  MUX2_X1 U25652 ( .A(_03332__PTR6), .B(_03332__PTR70), .S(P3_P1_InstQueueRd_Addr_PTR3), .Z(_02464__PTR6) );
  MUX2_X1 U25653 ( .A(_03332__PTR7), .B(_03332__PTR71), .S(P3_P1_InstQueueRd_Addr_PTR3), .Z(_02464__PTR7) );
  MUX2_X1 U25654 ( .A(_03331__PTR0), .B(_03331__PTR32), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR0) );
  MUX2_X1 U25655 ( .A(_03331__PTR1), .B(_03331__PTR33), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR1) );
  MUX2_X1 U25656 ( .A(_03331__PTR2), .B(_03331__PTR34), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR2) );
  MUX2_X1 U25657 ( .A(_03331__PTR3), .B(_03331__PTR35), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR3) );
  MUX2_X1 U25658 ( .A(_03331__PTR4), .B(_03331__PTR36), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR4) );
  MUX2_X1 U25659 ( .A(_03331__PTR5), .B(_03331__PTR37), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR5) );
  MUX2_X1 U25660 ( .A(_03331__PTR6), .B(_03331__PTR38), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR6) );
  MUX2_X1 U25661 ( .A(_03331__PTR7), .B(_03331__PTR39), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR7) );
  MUX2_X1 U25662 ( .A(_03331__PTR64), .B(_03331__PTR96), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR64) );
  MUX2_X1 U25663 ( .A(_03331__PTR65), .B(_03331__PTR97), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR65) );
  MUX2_X1 U25664 ( .A(_03331__PTR66), .B(_03331__PTR98), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR66) );
  MUX2_X1 U25665 ( .A(_03331__PTR67), .B(_03331__PTR99), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR67) );
  MUX2_X1 U25666 ( .A(_03331__PTR68), .B(_03331__PTR100), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR68) );
  MUX2_X1 U25667 ( .A(_03331__PTR69), .B(_03331__PTR101), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR69) );
  MUX2_X1 U25668 ( .A(_03331__PTR70), .B(_03331__PTR102), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR70) );
  MUX2_X1 U25669 ( .A(_03331__PTR71), .B(_03331__PTR103), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03332__PTR71) );
  MUX2_X1 U25670 ( .A(_03330__PTR0), .B(_03330__PTR16), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR0) );
  MUX2_X1 U25671 ( .A(_03330__PTR1), .B(_03330__PTR17), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR1) );
  MUX2_X1 U25672 ( .A(_03330__PTR2), .B(_03330__PTR18), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR2) );
  MUX2_X1 U25673 ( .A(_03330__PTR3), .B(_03330__PTR19), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR3) );
  MUX2_X1 U25674 ( .A(_03330__PTR4), .B(_03330__PTR20), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR4) );
  MUX2_X1 U25675 ( .A(_03330__PTR5), .B(_03330__PTR21), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR5) );
  MUX2_X1 U25676 ( .A(_03330__PTR6), .B(_03330__PTR22), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR6) );
  MUX2_X1 U25677 ( .A(_03330__PTR7), .B(_03330__PTR23), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR7) );
  MUX2_X1 U25678 ( .A(_03330__PTR32), .B(_03330__PTR48), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR32) );
  MUX2_X1 U25679 ( .A(_03330__PTR33), .B(_03330__PTR49), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR33) );
  MUX2_X1 U25680 ( .A(_03330__PTR34), .B(_03330__PTR50), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR34) );
  MUX2_X1 U25681 ( .A(_03330__PTR35), .B(_03330__PTR51), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR35) );
  MUX2_X1 U25682 ( .A(_03330__PTR36), .B(_03330__PTR52), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR36) );
  MUX2_X1 U25683 ( .A(_03330__PTR37), .B(_03330__PTR53), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR37) );
  MUX2_X1 U25684 ( .A(_03330__PTR38), .B(_03330__PTR54), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR38) );
  MUX2_X1 U25685 ( .A(_03330__PTR39), .B(_03330__PTR55), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR39) );
  MUX2_X1 U25686 ( .A(_03330__PTR64), .B(_03330__PTR80), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR64) );
  MUX2_X1 U25687 ( .A(_03330__PTR65), .B(_03330__PTR81), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR65) );
  MUX2_X1 U25688 ( .A(_03330__PTR66), .B(_03330__PTR82), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR66) );
  MUX2_X1 U25689 ( .A(_03330__PTR67), .B(_03330__PTR83), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR67) );
  MUX2_X1 U25690 ( .A(_03330__PTR68), .B(_03330__PTR84), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR68) );
  MUX2_X1 U25691 ( .A(_03330__PTR69), .B(_03330__PTR85), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR69) );
  MUX2_X1 U25692 ( .A(_03330__PTR70), .B(_03330__PTR86), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR70) );
  MUX2_X1 U25693 ( .A(_03330__PTR71), .B(_03330__PTR87), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR71) );
  MUX2_X1 U25694 ( .A(_03330__PTR96), .B(_03330__PTR112), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR96) );
  MUX2_X1 U25695 ( .A(_03330__PTR97), .B(_03330__PTR113), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR97) );
  MUX2_X1 U25696 ( .A(_03330__PTR98), .B(_03330__PTR114), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR98) );
  MUX2_X1 U25697 ( .A(_03330__PTR99), .B(_03330__PTR115), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR99) );
  MUX2_X1 U25698 ( .A(_03330__PTR100), .B(_03330__PTR116), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR100) );
  MUX2_X1 U25699 ( .A(_03330__PTR101), .B(_03330__PTR117), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR101) );
  MUX2_X1 U25700 ( .A(_03330__PTR102), .B(_03330__PTR118), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR102) );
  MUX2_X1 U25701 ( .A(_03330__PTR103), .B(_03330__PTR119), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03331__PTR103) );
  MUX2_X1 U25702 ( .A(P3_P1_InstQueue_PTR0_PTR0), .B(P3_P1_InstQueue_PTR1_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR0) );
  MUX2_X1 U25703 ( .A(P3_P1_InstQueue_PTR0_PTR1), .B(P3_P1_InstQueue_PTR1_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR1) );
  MUX2_X1 U25704 ( .A(P3_P1_InstQueue_PTR0_PTR2), .B(P3_P1_InstQueue_PTR1_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR2) );
  MUX2_X1 U25705 ( .A(P3_P1_InstQueue_PTR0_PTR3), .B(P3_P1_InstQueue_PTR1_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR3) );
  MUX2_X1 U25706 ( .A(P3_P1_InstQueue_PTR0_PTR4), .B(P3_P1_InstQueue_PTR1_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR4) );
  MUX2_X1 U25707 ( .A(P3_P1_InstQueue_PTR0_PTR5), .B(P3_P1_InstQueue_PTR1_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR5) );
  MUX2_X1 U25708 ( .A(P3_P1_InstQueue_PTR0_PTR6), .B(P3_P1_InstQueue_PTR1_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR6) );
  MUX2_X1 U25709 ( .A(P3_P1_InstQueue_PTR0_PTR7), .B(P3_P1_InstQueue_PTR1_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR7) );
  MUX2_X1 U25710 ( .A(P3_P1_InstQueue_PTR2_PTR0), .B(P3_P1_InstQueue_PTR3_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR16) );
  MUX2_X1 U25711 ( .A(P3_P1_InstQueue_PTR2_PTR1), .B(P3_P1_InstQueue_PTR3_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR17) );
  MUX2_X1 U25712 ( .A(P3_P1_InstQueue_PTR2_PTR2), .B(P3_P1_InstQueue_PTR3_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR18) );
  MUX2_X1 U25713 ( .A(P3_P1_InstQueue_PTR2_PTR3), .B(P3_P1_InstQueue_PTR3_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR19) );
  MUX2_X1 U25714 ( .A(P3_P1_InstQueue_PTR2_PTR4), .B(P3_P1_InstQueue_PTR3_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR20) );
  MUX2_X1 U25715 ( .A(P3_P1_InstQueue_PTR2_PTR5), .B(P3_P1_InstQueue_PTR3_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR21) );
  MUX2_X1 U25716 ( .A(P3_P1_InstQueue_PTR2_PTR6), .B(P3_P1_InstQueue_PTR3_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR22) );
  MUX2_X1 U25717 ( .A(P3_P1_InstQueue_PTR2_PTR7), .B(P3_P1_InstQueue_PTR3_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR23) );
  MUX2_X1 U25718 ( .A(P3_P1_InstQueue_PTR4_PTR0), .B(P3_P1_InstQueue_PTR5_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR32) );
  MUX2_X1 U25719 ( .A(P3_P1_InstQueue_PTR4_PTR1), .B(P3_P1_InstQueue_PTR5_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR33) );
  MUX2_X1 U25720 ( .A(P3_P1_InstQueue_PTR4_PTR2), .B(P3_P1_InstQueue_PTR5_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR34) );
  MUX2_X1 U25721 ( .A(P3_P1_InstQueue_PTR4_PTR3), .B(P3_P1_InstQueue_PTR5_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR35) );
  MUX2_X1 U25722 ( .A(P3_P1_InstQueue_PTR4_PTR4), .B(P3_P1_InstQueue_PTR5_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR36) );
  MUX2_X1 U25723 ( .A(P3_P1_InstQueue_PTR4_PTR5), .B(P3_P1_InstQueue_PTR5_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR37) );
  MUX2_X1 U25724 ( .A(P3_P1_InstQueue_PTR4_PTR6), .B(P3_P1_InstQueue_PTR5_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR38) );
  MUX2_X1 U25725 ( .A(P3_P1_InstQueue_PTR4_PTR7), .B(P3_P1_InstQueue_PTR5_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR39) );
  MUX2_X1 U25726 ( .A(P3_P1_InstQueue_PTR6_PTR0), .B(P3_P1_InstQueue_PTR7_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR48) );
  MUX2_X1 U25727 ( .A(P3_P1_InstQueue_PTR6_PTR1), .B(P3_P1_InstQueue_PTR7_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR49) );
  MUX2_X1 U25728 ( .A(P3_P1_InstQueue_PTR6_PTR2), .B(P3_P1_InstQueue_PTR7_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR50) );
  MUX2_X1 U25729 ( .A(P3_P1_InstQueue_PTR6_PTR3), .B(P3_P1_InstQueue_PTR7_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR51) );
  MUX2_X1 U25730 ( .A(P3_P1_InstQueue_PTR6_PTR4), .B(P3_P1_InstQueue_PTR7_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR52) );
  MUX2_X1 U25731 ( .A(P3_P1_InstQueue_PTR6_PTR5), .B(P3_P1_InstQueue_PTR7_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR53) );
  MUX2_X1 U25732 ( .A(P3_P1_InstQueue_PTR6_PTR6), .B(P3_P1_InstQueue_PTR7_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR54) );
  MUX2_X1 U25733 ( .A(P3_P1_InstQueue_PTR6_PTR7), .B(P3_P1_InstQueue_PTR7_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR55) );
  MUX2_X1 U25734 ( .A(P3_P1_InstQueue_PTR8_PTR0), .B(P3_P1_InstQueue_PTR9_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR64) );
  MUX2_X1 U25735 ( .A(P3_P1_InstQueue_PTR8_PTR1), .B(P3_P1_InstQueue_PTR9_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR65) );
  MUX2_X1 U25736 ( .A(P3_P1_InstQueue_PTR8_PTR2), .B(P3_P1_InstQueue_PTR9_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR66) );
  MUX2_X1 U25737 ( .A(P3_P1_InstQueue_PTR8_PTR3), .B(P3_P1_InstQueue_PTR9_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR67) );
  MUX2_X1 U25738 ( .A(P3_P1_InstQueue_PTR8_PTR4), .B(P3_P1_InstQueue_PTR9_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR68) );
  MUX2_X1 U25739 ( .A(P3_P1_InstQueue_PTR8_PTR5), .B(P3_P1_InstQueue_PTR9_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR69) );
  MUX2_X1 U25740 ( .A(P3_P1_InstQueue_PTR8_PTR6), .B(P3_P1_InstQueue_PTR9_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR70) );
  MUX2_X1 U25741 ( .A(P3_P1_InstQueue_PTR8_PTR7), .B(P3_P1_InstQueue_PTR9_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR71) );
  MUX2_X1 U25742 ( .A(P3_P1_InstQueue_PTR10_PTR0), .B(P3_P1_InstQueue_PTR11_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR80) );
  MUX2_X1 U25743 ( .A(P3_P1_InstQueue_PTR10_PTR1), .B(P3_P1_InstQueue_PTR11_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR81) );
  MUX2_X1 U25744 ( .A(P3_P1_InstQueue_PTR10_PTR2), .B(P3_P1_InstQueue_PTR11_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR82) );
  MUX2_X1 U25745 ( .A(P3_P1_InstQueue_PTR10_PTR3), .B(P3_P1_InstQueue_PTR11_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR83) );
  MUX2_X1 U25746 ( .A(P3_P1_InstQueue_PTR10_PTR4), .B(P3_P1_InstQueue_PTR11_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR84) );
  MUX2_X1 U25747 ( .A(P3_P1_InstQueue_PTR10_PTR5), .B(P3_P1_InstQueue_PTR11_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR85) );
  MUX2_X1 U25748 ( .A(P3_P1_InstQueue_PTR10_PTR6), .B(P3_P1_InstQueue_PTR11_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR86) );
  MUX2_X1 U25749 ( .A(P3_P1_InstQueue_PTR10_PTR7), .B(P3_P1_InstQueue_PTR11_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR87) );
  MUX2_X1 U25750 ( .A(P3_P1_InstQueue_PTR12_PTR0), .B(P3_P1_InstQueue_PTR13_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR96) );
  MUX2_X1 U25751 ( .A(P3_P1_InstQueue_PTR12_PTR1), .B(P3_P1_InstQueue_PTR13_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR97) );
  MUX2_X1 U25752 ( .A(P3_P1_InstQueue_PTR12_PTR2), .B(P3_P1_InstQueue_PTR13_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR98) );
  MUX2_X1 U25753 ( .A(P3_P1_InstQueue_PTR12_PTR3), .B(P3_P1_InstQueue_PTR13_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR99) );
  MUX2_X1 U25754 ( .A(P3_P1_InstQueue_PTR12_PTR4), .B(P3_P1_InstQueue_PTR13_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR100) );
  MUX2_X1 U25755 ( .A(P3_P1_InstQueue_PTR12_PTR5), .B(P3_P1_InstQueue_PTR13_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR101) );
  MUX2_X1 U25756 ( .A(P3_P1_InstQueue_PTR12_PTR6), .B(P3_P1_InstQueue_PTR13_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR102) );
  MUX2_X1 U25757 ( .A(P3_P1_InstQueue_PTR12_PTR7), .B(P3_P1_InstQueue_PTR13_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR103) );
  MUX2_X1 U25758 ( .A(P3_P1_InstQueue_PTR14_PTR0), .B(P3_P1_InstQueue_PTR15_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR112) );
  MUX2_X1 U25759 ( .A(P3_P1_InstQueue_PTR14_PTR1), .B(P3_P1_InstQueue_PTR15_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR113) );
  MUX2_X1 U25760 ( .A(P3_P1_InstQueue_PTR14_PTR2), .B(P3_P1_InstQueue_PTR15_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR114) );
  MUX2_X1 U25761 ( .A(P3_P1_InstQueue_PTR14_PTR3), .B(P3_P1_InstQueue_PTR15_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR115) );
  MUX2_X1 U25762 ( .A(P3_P1_InstQueue_PTR14_PTR4), .B(P3_P1_InstQueue_PTR15_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR116) );
  MUX2_X1 U25763 ( .A(P3_P1_InstQueue_PTR14_PTR5), .B(P3_P1_InstQueue_PTR15_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR117) );
  MUX2_X1 U25764 ( .A(P3_P1_InstQueue_PTR14_PTR6), .B(P3_P1_InstQueue_PTR15_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR118) );
  MUX2_X1 U25765 ( .A(P3_P1_InstQueue_PTR14_PTR7), .B(P3_P1_InstQueue_PTR15_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03330__PTR119) );
  MUX2_X1 U25766 ( .A(_03335__PTR0), .B(_03335__PTR64), .S(_02465__PTR6), .Z(_02466__PTR0) );
  MUX2_X1 U25767 ( .A(_03335__PTR1), .B(_03335__PTR65), .S(_02465__PTR6), .Z(_02466__PTR1) );
  MUX2_X1 U25768 ( .A(_03335__PTR2), .B(_03335__PTR66), .S(_02465__PTR6), .Z(_02466__PTR2) );
  MUX2_X1 U25769 ( .A(_03335__PTR3), .B(_03335__PTR67), .S(_02465__PTR6), .Z(_02466__PTR3) );
  MUX2_X1 U25770 ( .A(_03335__PTR4), .B(_03335__PTR68), .S(_02465__PTR6), .Z(_02466__PTR4) );
  MUX2_X1 U25771 ( .A(_03335__PTR5), .B(_03335__PTR69), .S(_02465__PTR6), .Z(_02466__PTR5) );
  MUX2_X1 U25772 ( .A(_03335__PTR6), .B(_03335__PTR70), .S(_02465__PTR6), .Z(_02466__PTR6) );
  MUX2_X1 U25773 ( .A(_03335__PTR7), .B(_03335__PTR71), .S(_02465__PTR6), .Z(_02466__PTR7) );
  MUX2_X1 U25774 ( .A(_03334__PTR0), .B(_03334__PTR32), .S(_02465__PTR5), .Z(_03335__PTR0) );
  MUX2_X1 U25775 ( .A(_03334__PTR1), .B(_03334__PTR33), .S(_02465__PTR5), .Z(_03335__PTR1) );
  MUX2_X1 U25776 ( .A(_03334__PTR2), .B(_03334__PTR34), .S(_02465__PTR5), .Z(_03335__PTR2) );
  MUX2_X1 U25777 ( .A(_03334__PTR3), .B(_03334__PTR35), .S(_02465__PTR5), .Z(_03335__PTR3) );
  MUX2_X1 U25778 ( .A(_03334__PTR4), .B(_03334__PTR36), .S(_02465__PTR5), .Z(_03335__PTR4) );
  MUX2_X1 U25779 ( .A(_03334__PTR5), .B(_03334__PTR37), .S(_02465__PTR5), .Z(_03335__PTR5) );
  MUX2_X1 U25780 ( .A(_03334__PTR6), .B(_03334__PTR38), .S(_02465__PTR5), .Z(_03335__PTR6) );
  MUX2_X1 U25781 ( .A(_03334__PTR7), .B(_03334__PTR39), .S(_02465__PTR5), .Z(_03335__PTR7) );
  MUX2_X1 U25782 ( .A(_03334__PTR64), .B(_03334__PTR96), .S(_02465__PTR5), .Z(_03335__PTR64) );
  MUX2_X1 U25783 ( .A(_03334__PTR65), .B(_03334__PTR97), .S(_02465__PTR5), .Z(_03335__PTR65) );
  MUX2_X1 U25784 ( .A(_03334__PTR66), .B(_03334__PTR98), .S(_02465__PTR5), .Z(_03335__PTR66) );
  MUX2_X1 U25785 ( .A(_03334__PTR67), .B(_03334__PTR99), .S(_02465__PTR5), .Z(_03335__PTR67) );
  MUX2_X1 U25786 ( .A(_03334__PTR68), .B(_03334__PTR100), .S(_02465__PTR5), .Z(_03335__PTR68) );
  MUX2_X1 U25787 ( .A(_03334__PTR69), .B(_03334__PTR101), .S(_02465__PTR5), .Z(_03335__PTR69) );
  MUX2_X1 U25788 ( .A(_03334__PTR70), .B(_03334__PTR102), .S(_02465__PTR5), .Z(_03335__PTR70) );
  MUX2_X1 U25789 ( .A(_03334__PTR71), .B(_03334__PTR103), .S(_02465__PTR5), .Z(_03335__PTR71) );
  MUX2_X1 U25790 ( .A(_03333__PTR0), .B(_03333__PTR16), .S(_02465__PTR4), .Z(_03334__PTR0) );
  MUX2_X1 U25791 ( .A(_03333__PTR1), .B(_03333__PTR17), .S(_02465__PTR4), .Z(_03334__PTR1) );
  MUX2_X1 U25792 ( .A(_03333__PTR2), .B(_03333__PTR18), .S(_02465__PTR4), .Z(_03334__PTR2) );
  MUX2_X1 U25793 ( .A(_03333__PTR3), .B(_03333__PTR19), .S(_02465__PTR4), .Z(_03334__PTR3) );
  MUX2_X1 U25794 ( .A(_03333__PTR4), .B(_03333__PTR20), .S(_02465__PTR4), .Z(_03334__PTR4) );
  MUX2_X1 U25795 ( .A(_03333__PTR5), .B(_03333__PTR21), .S(_02465__PTR4), .Z(_03334__PTR5) );
  MUX2_X1 U25796 ( .A(_03333__PTR6), .B(_03333__PTR22), .S(_02465__PTR4), .Z(_03334__PTR6) );
  MUX2_X1 U25797 ( .A(_03333__PTR7), .B(_03333__PTR23), .S(_02465__PTR4), .Z(_03334__PTR7) );
  MUX2_X1 U25798 ( .A(_03333__PTR32), .B(_03333__PTR48), .S(_02465__PTR4), .Z(_03334__PTR32) );
  MUX2_X1 U25799 ( .A(_03333__PTR33), .B(_03333__PTR49), .S(_02465__PTR4), .Z(_03334__PTR33) );
  MUX2_X1 U25800 ( .A(_03333__PTR34), .B(_03333__PTR50), .S(_02465__PTR4), .Z(_03334__PTR34) );
  MUX2_X1 U25801 ( .A(_03333__PTR35), .B(_03333__PTR51), .S(_02465__PTR4), .Z(_03334__PTR35) );
  MUX2_X1 U25802 ( .A(_03333__PTR36), .B(_03333__PTR52), .S(_02465__PTR4), .Z(_03334__PTR36) );
  MUX2_X1 U25803 ( .A(_03333__PTR37), .B(_03333__PTR53), .S(_02465__PTR4), .Z(_03334__PTR37) );
  MUX2_X1 U25804 ( .A(_03333__PTR38), .B(_03333__PTR54), .S(_02465__PTR4), .Z(_03334__PTR38) );
  MUX2_X1 U25805 ( .A(_03333__PTR39), .B(_03333__PTR55), .S(_02465__PTR4), .Z(_03334__PTR39) );
  MUX2_X1 U25806 ( .A(_03333__PTR64), .B(_03333__PTR80), .S(_02465__PTR4), .Z(_03334__PTR64) );
  MUX2_X1 U25807 ( .A(_03333__PTR65), .B(_03333__PTR81), .S(_02465__PTR4), .Z(_03334__PTR65) );
  MUX2_X1 U25808 ( .A(_03333__PTR66), .B(_03333__PTR82), .S(_02465__PTR4), .Z(_03334__PTR66) );
  MUX2_X1 U25809 ( .A(_03333__PTR67), .B(_03333__PTR83), .S(_02465__PTR4), .Z(_03334__PTR67) );
  MUX2_X1 U25810 ( .A(_03333__PTR68), .B(_03333__PTR84), .S(_02465__PTR4), .Z(_03334__PTR68) );
  MUX2_X1 U25811 ( .A(_03333__PTR69), .B(_03333__PTR85), .S(_02465__PTR4), .Z(_03334__PTR69) );
  MUX2_X1 U25812 ( .A(_03333__PTR70), .B(_03333__PTR86), .S(_02465__PTR4), .Z(_03334__PTR70) );
  MUX2_X1 U25813 ( .A(_03333__PTR71), .B(_03333__PTR87), .S(_02465__PTR4), .Z(_03334__PTR71) );
  MUX2_X1 U25814 ( .A(_03333__PTR96), .B(_03333__PTR112), .S(_02465__PTR4), .Z(_03334__PTR96) );
  MUX2_X1 U25815 ( .A(_03333__PTR97), .B(_03333__PTR113), .S(_02465__PTR4), .Z(_03334__PTR97) );
  MUX2_X1 U25816 ( .A(_03333__PTR98), .B(_03333__PTR114), .S(_02465__PTR4), .Z(_03334__PTR98) );
  MUX2_X1 U25817 ( .A(_03333__PTR99), .B(_03333__PTR115), .S(_02465__PTR4), .Z(_03334__PTR99) );
  MUX2_X1 U25818 ( .A(_03333__PTR100), .B(_03333__PTR116), .S(_02465__PTR4), .Z(_03334__PTR100) );
  MUX2_X1 U25819 ( .A(_03333__PTR101), .B(_03333__PTR117), .S(_02465__PTR4), .Z(_03334__PTR101) );
  MUX2_X1 U25820 ( .A(_03333__PTR102), .B(_03333__PTR118), .S(_02465__PTR4), .Z(_03334__PTR102) );
  MUX2_X1 U25821 ( .A(_03333__PTR103), .B(_03333__PTR119), .S(_02465__PTR4), .Z(_03334__PTR103) );
  MUX2_X1 U25822 ( .A(P3_P1_InstQueue_PTR1_PTR0), .B(P3_P1_InstQueue_PTR0_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR0) );
  MUX2_X1 U25823 ( .A(P3_P1_InstQueue_PTR1_PTR1), .B(P3_P1_InstQueue_PTR0_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR1) );
  MUX2_X1 U25824 ( .A(P3_P1_InstQueue_PTR1_PTR2), .B(P3_P1_InstQueue_PTR0_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR2) );
  MUX2_X1 U25825 ( .A(P3_P1_InstQueue_PTR1_PTR3), .B(P3_P1_InstQueue_PTR0_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR3) );
  MUX2_X1 U25826 ( .A(P3_P1_InstQueue_PTR1_PTR4), .B(P3_P1_InstQueue_PTR0_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR4) );
  MUX2_X1 U25827 ( .A(P3_P1_InstQueue_PTR1_PTR5), .B(P3_P1_InstQueue_PTR0_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR5) );
  MUX2_X1 U25828 ( .A(P3_P1_InstQueue_PTR1_PTR6), .B(P3_P1_InstQueue_PTR0_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR6) );
  MUX2_X1 U25829 ( .A(P3_P1_InstQueue_PTR1_PTR7), .B(P3_P1_InstQueue_PTR0_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR7) );
  MUX2_X1 U25830 ( .A(P3_P1_InstQueue_PTR3_PTR0), .B(P3_P1_InstQueue_PTR2_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR16) );
  MUX2_X1 U25831 ( .A(P3_P1_InstQueue_PTR3_PTR1), .B(P3_P1_InstQueue_PTR2_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR17) );
  MUX2_X1 U25832 ( .A(P3_P1_InstQueue_PTR3_PTR2), .B(P3_P1_InstQueue_PTR2_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR18) );
  MUX2_X1 U25833 ( .A(P3_P1_InstQueue_PTR3_PTR3), .B(P3_P1_InstQueue_PTR2_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR19) );
  MUX2_X1 U25834 ( .A(P3_P1_InstQueue_PTR3_PTR4), .B(P3_P1_InstQueue_PTR2_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR20) );
  MUX2_X1 U25835 ( .A(P3_P1_InstQueue_PTR3_PTR5), .B(P3_P1_InstQueue_PTR2_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR21) );
  MUX2_X1 U25836 ( .A(P3_P1_InstQueue_PTR3_PTR6), .B(P3_P1_InstQueue_PTR2_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR22) );
  MUX2_X1 U25837 ( .A(P3_P1_InstQueue_PTR3_PTR7), .B(P3_P1_InstQueue_PTR2_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR23) );
  MUX2_X1 U25838 ( .A(P3_P1_InstQueue_PTR5_PTR0), .B(P3_P1_InstQueue_PTR4_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR32) );
  MUX2_X1 U25839 ( .A(P3_P1_InstQueue_PTR5_PTR1), .B(P3_P1_InstQueue_PTR4_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR33) );
  MUX2_X1 U25840 ( .A(P3_P1_InstQueue_PTR5_PTR2), .B(P3_P1_InstQueue_PTR4_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR34) );
  MUX2_X1 U25841 ( .A(P3_P1_InstQueue_PTR5_PTR3), .B(P3_P1_InstQueue_PTR4_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR35) );
  MUX2_X1 U25842 ( .A(P3_P1_InstQueue_PTR5_PTR4), .B(P3_P1_InstQueue_PTR4_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR36) );
  MUX2_X1 U25843 ( .A(P3_P1_InstQueue_PTR5_PTR5), .B(P3_P1_InstQueue_PTR4_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR37) );
  MUX2_X1 U25844 ( .A(P3_P1_InstQueue_PTR5_PTR6), .B(P3_P1_InstQueue_PTR4_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR38) );
  MUX2_X1 U25845 ( .A(P3_P1_InstQueue_PTR5_PTR7), .B(P3_P1_InstQueue_PTR4_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR39) );
  MUX2_X1 U25846 ( .A(P3_P1_InstQueue_PTR7_PTR0), .B(P3_P1_InstQueue_PTR6_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR48) );
  MUX2_X1 U25847 ( .A(P3_P1_InstQueue_PTR7_PTR1), .B(P3_P1_InstQueue_PTR6_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR49) );
  MUX2_X1 U25848 ( .A(P3_P1_InstQueue_PTR7_PTR2), .B(P3_P1_InstQueue_PTR6_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR50) );
  MUX2_X1 U25849 ( .A(P3_P1_InstQueue_PTR7_PTR3), .B(P3_P1_InstQueue_PTR6_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR51) );
  MUX2_X1 U25850 ( .A(P3_P1_InstQueue_PTR7_PTR4), .B(P3_P1_InstQueue_PTR6_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR52) );
  MUX2_X1 U25851 ( .A(P3_P1_InstQueue_PTR7_PTR5), .B(P3_P1_InstQueue_PTR6_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR53) );
  MUX2_X1 U25852 ( .A(P3_P1_InstQueue_PTR7_PTR6), .B(P3_P1_InstQueue_PTR6_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR54) );
  MUX2_X1 U25853 ( .A(P3_P1_InstQueue_PTR7_PTR7), .B(P3_P1_InstQueue_PTR6_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR55) );
  MUX2_X1 U25854 ( .A(P3_P1_InstQueue_PTR9_PTR0), .B(P3_P1_InstQueue_PTR8_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR64) );
  MUX2_X1 U25855 ( .A(P3_P1_InstQueue_PTR9_PTR1), .B(P3_P1_InstQueue_PTR8_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR65) );
  MUX2_X1 U25856 ( .A(P3_P1_InstQueue_PTR9_PTR2), .B(P3_P1_InstQueue_PTR8_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR66) );
  MUX2_X1 U25857 ( .A(P3_P1_InstQueue_PTR9_PTR3), .B(P3_P1_InstQueue_PTR8_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR67) );
  MUX2_X1 U25858 ( .A(P3_P1_InstQueue_PTR9_PTR4), .B(P3_P1_InstQueue_PTR8_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR68) );
  MUX2_X1 U25859 ( .A(P3_P1_InstQueue_PTR9_PTR5), .B(P3_P1_InstQueue_PTR8_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR69) );
  MUX2_X1 U25860 ( .A(P3_P1_InstQueue_PTR9_PTR6), .B(P3_P1_InstQueue_PTR8_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR70) );
  MUX2_X1 U25861 ( .A(P3_P1_InstQueue_PTR9_PTR7), .B(P3_P1_InstQueue_PTR8_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR71) );
  MUX2_X1 U25862 ( .A(P3_P1_InstQueue_PTR11_PTR0), .B(P3_P1_InstQueue_PTR10_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR80) );
  MUX2_X1 U25863 ( .A(P3_P1_InstQueue_PTR11_PTR1), .B(P3_P1_InstQueue_PTR10_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR81) );
  MUX2_X1 U25864 ( .A(P3_P1_InstQueue_PTR11_PTR2), .B(P3_P1_InstQueue_PTR10_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR82) );
  MUX2_X1 U25865 ( .A(P3_P1_InstQueue_PTR11_PTR3), .B(P3_P1_InstQueue_PTR10_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR83) );
  MUX2_X1 U25866 ( .A(P3_P1_InstQueue_PTR11_PTR4), .B(P3_P1_InstQueue_PTR10_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR84) );
  MUX2_X1 U25867 ( .A(P3_P1_InstQueue_PTR11_PTR5), .B(P3_P1_InstQueue_PTR10_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR85) );
  MUX2_X1 U25868 ( .A(P3_P1_InstQueue_PTR11_PTR6), .B(P3_P1_InstQueue_PTR10_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR86) );
  MUX2_X1 U25869 ( .A(P3_P1_InstQueue_PTR11_PTR7), .B(P3_P1_InstQueue_PTR10_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR87) );
  MUX2_X1 U25870 ( .A(P3_P1_InstQueue_PTR13_PTR0), .B(P3_P1_InstQueue_PTR12_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR96) );
  MUX2_X1 U25871 ( .A(P3_P1_InstQueue_PTR13_PTR1), .B(P3_P1_InstQueue_PTR12_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR97) );
  MUX2_X1 U25872 ( .A(P3_P1_InstQueue_PTR13_PTR2), .B(P3_P1_InstQueue_PTR12_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR98) );
  MUX2_X1 U25873 ( .A(P3_P1_InstQueue_PTR13_PTR3), .B(P3_P1_InstQueue_PTR12_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR99) );
  MUX2_X1 U25874 ( .A(P3_P1_InstQueue_PTR13_PTR4), .B(P3_P1_InstQueue_PTR12_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR100) );
  MUX2_X1 U25875 ( .A(P3_P1_InstQueue_PTR13_PTR5), .B(P3_P1_InstQueue_PTR12_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR101) );
  MUX2_X1 U25876 ( .A(P3_P1_InstQueue_PTR13_PTR6), .B(P3_P1_InstQueue_PTR12_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR102) );
  MUX2_X1 U25877 ( .A(P3_P1_InstQueue_PTR13_PTR7), .B(P3_P1_InstQueue_PTR12_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR103) );
  MUX2_X1 U25878 ( .A(P3_P1_InstQueue_PTR15_PTR0), .B(P3_P1_InstQueue_PTR14_PTR0), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR112) );
  MUX2_X1 U25879 ( .A(P3_P1_InstQueue_PTR15_PTR1), .B(P3_P1_InstQueue_PTR14_PTR1), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR113) );
  MUX2_X1 U25880 ( .A(P3_P1_InstQueue_PTR15_PTR2), .B(P3_P1_InstQueue_PTR14_PTR2), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR114) );
  MUX2_X1 U25881 ( .A(P3_P1_InstQueue_PTR15_PTR3), .B(P3_P1_InstQueue_PTR14_PTR3), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR115) );
  MUX2_X1 U25882 ( .A(P3_P1_InstQueue_PTR15_PTR4), .B(P3_P1_InstQueue_PTR14_PTR4), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR116) );
  MUX2_X1 U25883 ( .A(P3_P1_InstQueue_PTR15_PTR5), .B(P3_P1_InstQueue_PTR14_PTR5), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR117) );
  MUX2_X1 U25884 ( .A(P3_P1_InstQueue_PTR15_PTR6), .B(P3_P1_InstQueue_PTR14_PTR6), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR118) );
  MUX2_X1 U25885 ( .A(P3_P1_InstQueue_PTR15_PTR7), .B(P3_P1_InstQueue_PTR14_PTR7), .S(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03333__PTR119) );
  MUX2_X1 U25886 ( .A(_03336__PTR0), .B(_03336__PTR64), .S(_02467__PTR6), .Z(_02468__PTR0) );
  MUX2_X1 U25887 ( .A(_03336__PTR1), .B(_03336__PTR65), .S(_02467__PTR6), .Z(_02468__PTR1) );
  MUX2_X1 U25888 ( .A(_03336__PTR2), .B(_03336__PTR66), .S(_02467__PTR6), .Z(_02468__PTR2) );
  MUX2_X1 U25889 ( .A(_03336__PTR3), .B(_03336__PTR67), .S(_02467__PTR6), .Z(_02468__PTR3) );
  MUX2_X1 U25890 ( .A(_03336__PTR4), .B(_03336__PTR68), .S(_02467__PTR6), .Z(_02468__PTR4) );
  MUX2_X1 U25891 ( .A(_03336__PTR5), .B(_03336__PTR69), .S(_02467__PTR6), .Z(_02468__PTR5) );
  MUX2_X1 U25892 ( .A(_03336__PTR6), .B(_03336__PTR70), .S(_02467__PTR6), .Z(_02468__PTR6) );
  MUX2_X1 U25893 ( .A(_03336__PTR7), .B(_03336__PTR71), .S(_02467__PTR6), .Z(_02468__PTR7) );
  MUX2_X1 U25894 ( .A(_03331__PTR32), .B(_03331__PTR0), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR0) );
  MUX2_X1 U25895 ( .A(_03331__PTR33), .B(_03331__PTR1), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR1) );
  MUX2_X1 U25896 ( .A(_03331__PTR34), .B(_03331__PTR2), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR2) );
  MUX2_X1 U25897 ( .A(_03331__PTR35), .B(_03331__PTR3), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR3) );
  MUX2_X1 U25898 ( .A(_03331__PTR36), .B(_03331__PTR4), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR4) );
  MUX2_X1 U25899 ( .A(_03331__PTR37), .B(_03331__PTR5), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR5) );
  MUX2_X1 U25900 ( .A(_03331__PTR38), .B(_03331__PTR6), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR6) );
  MUX2_X1 U25901 ( .A(_03331__PTR39), .B(_03331__PTR7), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR7) );
  MUX2_X1 U25902 ( .A(_03331__PTR96), .B(_03331__PTR64), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR64) );
  MUX2_X1 U25903 ( .A(_03331__PTR97), .B(_03331__PTR65), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR65) );
  MUX2_X1 U25904 ( .A(_03331__PTR98), .B(_03331__PTR66), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR66) );
  MUX2_X1 U25905 ( .A(_03331__PTR99), .B(_03331__PTR67), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR67) );
  MUX2_X1 U25906 ( .A(_03331__PTR100), .B(_03331__PTR68), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR68) );
  MUX2_X1 U25907 ( .A(_03331__PTR101), .B(_03331__PTR69), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR69) );
  MUX2_X1 U25908 ( .A(_03331__PTR102), .B(_03331__PTR70), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR70) );
  MUX2_X1 U25909 ( .A(_03331__PTR103), .B(_03331__PTR71), .S(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03336__PTR71) );
  MUX2_X1 U25910 ( .A(_03338__PTR0), .B(_03338__PTR64), .S(_02469__PTR6), .Z(_02470__PTR0) );
  MUX2_X1 U25911 ( .A(_03338__PTR1), .B(_03338__PTR65), .S(_02469__PTR6), .Z(_02470__PTR1) );
  MUX2_X1 U25912 ( .A(_03338__PTR2), .B(_03338__PTR66), .S(_02469__PTR6), .Z(_02470__PTR2) );
  MUX2_X1 U25913 ( .A(_03338__PTR3), .B(_03338__PTR67), .S(_02469__PTR6), .Z(_02470__PTR3) );
  MUX2_X1 U25914 ( .A(_03338__PTR4), .B(_03338__PTR68), .S(_02469__PTR6), .Z(_02470__PTR4) );
  MUX2_X1 U25915 ( .A(_03338__PTR5), .B(_03338__PTR69), .S(_02469__PTR6), .Z(_02470__PTR5) );
  MUX2_X1 U25916 ( .A(_03338__PTR6), .B(_03338__PTR70), .S(_02469__PTR6), .Z(_02470__PTR6) );
  MUX2_X1 U25917 ( .A(_03338__PTR7), .B(_03338__PTR71), .S(_02469__PTR6), .Z(_02470__PTR7) );
  MUX2_X1 U25918 ( .A(_03337__PTR0), .B(_03337__PTR32), .S(_02469__PTR5), .Z(_03338__PTR0) );
  MUX2_X1 U25919 ( .A(_03337__PTR1), .B(_03337__PTR33), .S(_02469__PTR5), .Z(_03338__PTR1) );
  MUX2_X1 U25920 ( .A(_03337__PTR2), .B(_03337__PTR34), .S(_02469__PTR5), .Z(_03338__PTR2) );
  MUX2_X1 U25921 ( .A(_03337__PTR3), .B(_03337__PTR35), .S(_02469__PTR5), .Z(_03338__PTR3) );
  MUX2_X1 U25922 ( .A(_03337__PTR4), .B(_03337__PTR36), .S(_02469__PTR5), .Z(_03338__PTR4) );
  MUX2_X1 U25923 ( .A(_03337__PTR5), .B(_03337__PTR37), .S(_02469__PTR5), .Z(_03338__PTR5) );
  MUX2_X1 U25924 ( .A(_03337__PTR6), .B(_03337__PTR38), .S(_02469__PTR5), .Z(_03338__PTR6) );
  MUX2_X1 U25925 ( .A(_03337__PTR7), .B(_03337__PTR39), .S(_02469__PTR5), .Z(_03338__PTR7) );
  MUX2_X1 U25926 ( .A(_03337__PTR64), .B(_03337__PTR96), .S(_02469__PTR5), .Z(_03338__PTR64) );
  MUX2_X1 U25927 ( .A(_03337__PTR65), .B(_03337__PTR97), .S(_02469__PTR5), .Z(_03338__PTR65) );
  MUX2_X1 U25928 ( .A(_03337__PTR66), .B(_03337__PTR98), .S(_02469__PTR5), .Z(_03338__PTR66) );
  MUX2_X1 U25929 ( .A(_03337__PTR67), .B(_03337__PTR99), .S(_02469__PTR5), .Z(_03338__PTR67) );
  MUX2_X1 U25930 ( .A(_03337__PTR68), .B(_03337__PTR100), .S(_02469__PTR5), .Z(_03338__PTR68) );
  MUX2_X1 U25931 ( .A(_03337__PTR69), .B(_03337__PTR101), .S(_02469__PTR5), .Z(_03338__PTR69) );
  MUX2_X1 U25932 ( .A(_03337__PTR70), .B(_03337__PTR102), .S(_02469__PTR5), .Z(_03338__PTR70) );
  MUX2_X1 U25933 ( .A(_03337__PTR71), .B(_03337__PTR103), .S(_02469__PTR5), .Z(_03338__PTR71) );
  MUX2_X1 U25934 ( .A(_03333__PTR0), .B(_03333__PTR16), .S(_02469__PTR4), .Z(_03337__PTR0) );
  MUX2_X1 U25935 ( .A(_03333__PTR1), .B(_03333__PTR17), .S(_02469__PTR4), .Z(_03337__PTR1) );
  MUX2_X1 U25936 ( .A(_03333__PTR2), .B(_03333__PTR18), .S(_02469__PTR4), .Z(_03337__PTR2) );
  MUX2_X1 U25937 ( .A(_03333__PTR3), .B(_03333__PTR19), .S(_02469__PTR4), .Z(_03337__PTR3) );
  MUX2_X1 U25938 ( .A(_03333__PTR4), .B(_03333__PTR20), .S(_02469__PTR4), .Z(_03337__PTR4) );
  MUX2_X1 U25939 ( .A(_03333__PTR5), .B(_03333__PTR21), .S(_02469__PTR4), .Z(_03337__PTR5) );
  MUX2_X1 U25940 ( .A(_03333__PTR6), .B(_03333__PTR22), .S(_02469__PTR4), .Z(_03337__PTR6) );
  MUX2_X1 U25941 ( .A(_03333__PTR7), .B(_03333__PTR23), .S(_02469__PTR4), .Z(_03337__PTR7) );
  MUX2_X1 U25942 ( .A(_03333__PTR32), .B(_03333__PTR48), .S(_02469__PTR4), .Z(_03337__PTR32) );
  MUX2_X1 U25943 ( .A(_03333__PTR33), .B(_03333__PTR49), .S(_02469__PTR4), .Z(_03337__PTR33) );
  MUX2_X1 U25944 ( .A(_03333__PTR34), .B(_03333__PTR50), .S(_02469__PTR4), .Z(_03337__PTR34) );
  MUX2_X1 U25945 ( .A(_03333__PTR35), .B(_03333__PTR51), .S(_02469__PTR4), .Z(_03337__PTR35) );
  MUX2_X1 U25946 ( .A(_03333__PTR36), .B(_03333__PTR52), .S(_02469__PTR4), .Z(_03337__PTR36) );
  MUX2_X1 U25947 ( .A(_03333__PTR37), .B(_03333__PTR53), .S(_02469__PTR4), .Z(_03337__PTR37) );
  MUX2_X1 U25948 ( .A(_03333__PTR38), .B(_03333__PTR54), .S(_02469__PTR4), .Z(_03337__PTR38) );
  MUX2_X1 U25949 ( .A(_03333__PTR39), .B(_03333__PTR55), .S(_02469__PTR4), .Z(_03337__PTR39) );
  MUX2_X1 U25950 ( .A(_03333__PTR64), .B(_03333__PTR80), .S(_02469__PTR4), .Z(_03337__PTR64) );
  MUX2_X1 U25951 ( .A(_03333__PTR65), .B(_03333__PTR81), .S(_02469__PTR4), .Z(_03337__PTR65) );
  MUX2_X1 U25952 ( .A(_03333__PTR66), .B(_03333__PTR82), .S(_02469__PTR4), .Z(_03337__PTR66) );
  MUX2_X1 U25953 ( .A(_03333__PTR67), .B(_03333__PTR83), .S(_02469__PTR4), .Z(_03337__PTR67) );
  MUX2_X1 U25954 ( .A(_03333__PTR68), .B(_03333__PTR84), .S(_02469__PTR4), .Z(_03337__PTR68) );
  MUX2_X1 U25955 ( .A(_03333__PTR69), .B(_03333__PTR85), .S(_02469__PTR4), .Z(_03337__PTR69) );
  MUX2_X1 U25956 ( .A(_03333__PTR70), .B(_03333__PTR86), .S(_02469__PTR4), .Z(_03337__PTR70) );
  MUX2_X1 U25957 ( .A(_03333__PTR71), .B(_03333__PTR87), .S(_02469__PTR4), .Z(_03337__PTR71) );
  MUX2_X1 U25958 ( .A(_03333__PTR96), .B(_03333__PTR112), .S(_02469__PTR4), .Z(_03337__PTR96) );
  MUX2_X1 U25959 ( .A(_03333__PTR97), .B(_03333__PTR113), .S(_02469__PTR4), .Z(_03337__PTR97) );
  MUX2_X1 U25960 ( .A(_03333__PTR98), .B(_03333__PTR114), .S(_02469__PTR4), .Z(_03337__PTR98) );
  MUX2_X1 U25961 ( .A(_03333__PTR99), .B(_03333__PTR115), .S(_02469__PTR4), .Z(_03337__PTR99) );
  MUX2_X1 U25962 ( .A(_03333__PTR100), .B(_03333__PTR116), .S(_02469__PTR4), .Z(_03337__PTR100) );
  MUX2_X1 U25963 ( .A(_03333__PTR101), .B(_03333__PTR117), .S(_02469__PTR4), .Z(_03337__PTR101) );
  MUX2_X1 U25964 ( .A(_03333__PTR102), .B(_03333__PTR118), .S(_02469__PTR4), .Z(_03337__PTR102) );
  MUX2_X1 U25965 ( .A(_03333__PTR103), .B(_03333__PTR119), .S(_02469__PTR4), .Z(_03337__PTR103) );
  MUX2_X1 U25966 ( .A(_03340__PTR0), .B(_03340__PTR64), .S(_02471__PTR6), .Z(_02472__PTR0) );
  MUX2_X1 U25967 ( .A(_03340__PTR1), .B(_03340__PTR65), .S(_02471__PTR6), .Z(_02472__PTR1) );
  MUX2_X1 U25968 ( .A(_03340__PTR2), .B(_03340__PTR66), .S(_02471__PTR6), .Z(_02472__PTR2) );
  MUX2_X1 U25969 ( .A(_03340__PTR3), .B(_03340__PTR67), .S(_02471__PTR6), .Z(_02472__PTR3) );
  MUX2_X1 U25970 ( .A(_03340__PTR4), .B(_03340__PTR68), .S(_02471__PTR6), .Z(_02472__PTR4) );
  MUX2_X1 U25971 ( .A(_03340__PTR5), .B(_03340__PTR69), .S(_02471__PTR6), .Z(_02472__PTR5) );
  MUX2_X1 U25972 ( .A(_03340__PTR6), .B(_03340__PTR70), .S(_02471__PTR6), .Z(_02472__PTR6) );
  MUX2_X1 U25973 ( .A(_03340__PTR7), .B(_03340__PTR71), .S(_02471__PTR6), .Z(_02472__PTR7) );
  MUX2_X1 U25974 ( .A(_03339__PTR0), .B(_03339__PTR32), .S(_02471__PTR5), .Z(_03340__PTR0) );
  MUX2_X1 U25975 ( .A(_03339__PTR1), .B(_03339__PTR33), .S(_02471__PTR5), .Z(_03340__PTR1) );
  MUX2_X1 U25976 ( .A(_03339__PTR2), .B(_03339__PTR34), .S(_02471__PTR5), .Z(_03340__PTR2) );
  MUX2_X1 U25977 ( .A(_03339__PTR3), .B(_03339__PTR35), .S(_02471__PTR5), .Z(_03340__PTR3) );
  MUX2_X1 U25978 ( .A(_03339__PTR4), .B(_03339__PTR36), .S(_02471__PTR5), .Z(_03340__PTR4) );
  MUX2_X1 U25979 ( .A(_03339__PTR5), .B(_03339__PTR37), .S(_02471__PTR5), .Z(_03340__PTR5) );
  MUX2_X1 U25980 ( .A(_03339__PTR6), .B(_03339__PTR38), .S(_02471__PTR5), .Z(_03340__PTR6) );
  MUX2_X1 U25981 ( .A(_03339__PTR7), .B(_03339__PTR39), .S(_02471__PTR5), .Z(_03340__PTR7) );
  MUX2_X1 U25982 ( .A(_03339__PTR64), .B(_03339__PTR96), .S(_02471__PTR5), .Z(_03340__PTR64) );
  MUX2_X1 U25983 ( .A(_03339__PTR65), .B(_03339__PTR97), .S(_02471__PTR5), .Z(_03340__PTR65) );
  MUX2_X1 U25984 ( .A(_03339__PTR66), .B(_03339__PTR98), .S(_02471__PTR5), .Z(_03340__PTR66) );
  MUX2_X1 U25985 ( .A(_03339__PTR67), .B(_03339__PTR99), .S(_02471__PTR5), .Z(_03340__PTR67) );
  MUX2_X1 U25986 ( .A(_03339__PTR68), .B(_03339__PTR100), .S(_02471__PTR5), .Z(_03340__PTR68) );
  MUX2_X1 U25987 ( .A(_03339__PTR69), .B(_03339__PTR101), .S(_02471__PTR5), .Z(_03340__PTR69) );
  MUX2_X1 U25988 ( .A(_03339__PTR70), .B(_03339__PTR102), .S(_02471__PTR5), .Z(_03340__PTR70) );
  MUX2_X1 U25989 ( .A(_03339__PTR71), .B(_03339__PTR103), .S(_02471__PTR5), .Z(_03340__PTR71) );
  MUX2_X1 U25990 ( .A(_03330__PTR16), .B(_03330__PTR0), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR0) );
  MUX2_X1 U25991 ( .A(_03330__PTR17), .B(_03330__PTR1), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR1) );
  MUX2_X1 U25992 ( .A(_03330__PTR18), .B(_03330__PTR2), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR2) );
  MUX2_X1 U25993 ( .A(_03330__PTR19), .B(_03330__PTR3), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR3) );
  MUX2_X1 U25994 ( .A(_03330__PTR20), .B(_03330__PTR4), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR4) );
  MUX2_X1 U25995 ( .A(_03330__PTR21), .B(_03330__PTR5), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR5) );
  MUX2_X1 U25996 ( .A(_03330__PTR22), .B(_03330__PTR6), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR6) );
  MUX2_X1 U25997 ( .A(_03330__PTR23), .B(_03330__PTR7), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR7) );
  MUX2_X1 U25998 ( .A(_03330__PTR48), .B(_03330__PTR32), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR32) );
  MUX2_X1 U25999 ( .A(_03330__PTR49), .B(_03330__PTR33), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR33) );
  MUX2_X1 U26000 ( .A(_03330__PTR50), .B(_03330__PTR34), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR34) );
  MUX2_X1 U26001 ( .A(_03330__PTR51), .B(_03330__PTR35), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR35) );
  MUX2_X1 U26002 ( .A(_03330__PTR52), .B(_03330__PTR36), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR36) );
  MUX2_X1 U26003 ( .A(_03330__PTR53), .B(_03330__PTR37), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR37) );
  MUX2_X1 U26004 ( .A(_03330__PTR54), .B(_03330__PTR38), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR38) );
  MUX2_X1 U26005 ( .A(_03330__PTR55), .B(_03330__PTR39), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR39) );
  MUX2_X1 U26006 ( .A(_03330__PTR80), .B(_03330__PTR64), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR64) );
  MUX2_X1 U26007 ( .A(_03330__PTR81), .B(_03330__PTR65), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR65) );
  MUX2_X1 U26008 ( .A(_03330__PTR82), .B(_03330__PTR66), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR66) );
  MUX2_X1 U26009 ( .A(_03330__PTR83), .B(_03330__PTR67), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR67) );
  MUX2_X1 U26010 ( .A(_03330__PTR84), .B(_03330__PTR68), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR68) );
  MUX2_X1 U26011 ( .A(_03330__PTR85), .B(_03330__PTR69), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR69) );
  MUX2_X1 U26012 ( .A(_03330__PTR86), .B(_03330__PTR70), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR70) );
  MUX2_X1 U26013 ( .A(_03330__PTR87), .B(_03330__PTR71), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR71) );
  MUX2_X1 U26014 ( .A(_03330__PTR112), .B(_03330__PTR96), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR96) );
  MUX2_X1 U26015 ( .A(_03330__PTR113), .B(_03330__PTR97), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR97) );
  MUX2_X1 U26016 ( .A(_03330__PTR114), .B(_03330__PTR98), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR98) );
  MUX2_X1 U26017 ( .A(_03330__PTR115), .B(_03330__PTR99), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR99) );
  MUX2_X1 U26018 ( .A(_03330__PTR116), .B(_03330__PTR100), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR100) );
  MUX2_X1 U26019 ( .A(_03330__PTR117), .B(_03330__PTR101), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR101) );
  MUX2_X1 U26020 ( .A(_03330__PTR118), .B(_03330__PTR102), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR102) );
  MUX2_X1 U26021 ( .A(_03330__PTR119), .B(_03330__PTR103), .S(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03339__PTR103) );
  MUX2_X1 U26022 ( .A(_03342__PTR0), .B(_03342__PTR128), .S(P3_P1_State2_PTR2), .Z(_03343__PTR0) );
  MUX2_X1 U26023 ( .A(_03342__PTR1), .B(_03342__PTR129), .S(P3_P1_State2_PTR2), .Z(_03343__PTR1) );
  MUX2_X1 U26024 ( .A(_03342__PTR2), .B(_03342__PTR130), .S(P3_P1_State2_PTR2), .Z(_03343__PTR2) );
  MUX2_X1 U26025 ( .A(_03342__PTR3), .B(_03342__PTR131), .S(P3_P1_State2_PTR2), .Z(_03343__PTR3) );
  MUX2_X1 U26026 ( .A(_03342__PTR4), .B(_03342__PTR132), .S(P3_P1_State2_PTR2), .Z(_03343__PTR4) );
  MUX2_X1 U26027 ( .A(_03342__PTR5), .B(_03342__PTR133), .S(P3_P1_State2_PTR2), .Z(_03343__PTR5) );
  MUX2_X1 U26028 ( .A(_03342__PTR6), .B(_03342__PTR134), .S(P3_P1_State2_PTR2), .Z(_03343__PTR6) );
  MUX2_X1 U26029 ( .A(_03342__PTR7), .B(_03342__PTR135), .S(P3_P1_State2_PTR2), .Z(_03343__PTR7) );
  MUX2_X1 U26030 ( .A(_03342__PTR8), .B(_03342__PTR136), .S(P3_P1_State2_PTR2), .Z(_03343__PTR8) );
  MUX2_X1 U26031 ( .A(_03342__PTR9), .B(_03342__PTR137), .S(P3_P1_State2_PTR2), .Z(_03343__PTR9) );
  MUX2_X1 U26032 ( .A(_03342__PTR10), .B(_03342__PTR138), .S(P3_P1_State2_PTR2), .Z(_03343__PTR10) );
  MUX2_X1 U26033 ( .A(_03342__PTR11), .B(_03342__PTR139), .S(P3_P1_State2_PTR2), .Z(_03343__PTR11) );
  MUX2_X1 U26034 ( .A(_03342__PTR12), .B(_03342__PTR140), .S(P3_P1_State2_PTR2), .Z(_03343__PTR12) );
  MUX2_X1 U26035 ( .A(_03342__PTR13), .B(_03342__PTR141), .S(P3_P1_State2_PTR2), .Z(_03343__PTR13) );
  MUX2_X1 U26036 ( .A(_03342__PTR14), .B(_03342__PTR142), .S(P3_P1_State2_PTR2), .Z(_03343__PTR14) );
  MUX2_X1 U26037 ( .A(_03342__PTR15), .B(_03342__PTR143), .S(P3_P1_State2_PTR2), .Z(_03343__PTR15) );
  MUX2_X1 U26038 ( .A(_03342__PTR16), .B(_03342__PTR144), .S(P3_P1_State2_PTR2), .Z(_03343__PTR16) );
  MUX2_X1 U26039 ( .A(_03342__PTR17), .B(_03342__PTR145), .S(P3_P1_State2_PTR2), .Z(_03343__PTR17) );
  MUX2_X1 U26040 ( .A(_03342__PTR18), .B(_03342__PTR146), .S(P3_P1_State2_PTR2), .Z(_03343__PTR18) );
  MUX2_X1 U26041 ( .A(_03342__PTR19), .B(_03342__PTR147), .S(P3_P1_State2_PTR2), .Z(_03343__PTR19) );
  MUX2_X1 U26042 ( .A(_03342__PTR20), .B(_03342__PTR148), .S(P3_P1_State2_PTR2), .Z(_03343__PTR20) );
  MUX2_X1 U26043 ( .A(_03342__PTR21), .B(_03342__PTR149), .S(P3_P1_State2_PTR2), .Z(_03343__PTR21) );
  MUX2_X1 U26044 ( .A(_03342__PTR22), .B(_03342__PTR150), .S(P3_P1_State2_PTR2), .Z(_03343__PTR22) );
  MUX2_X1 U26045 ( .A(_03342__PTR23), .B(_03342__PTR151), .S(P3_P1_State2_PTR2), .Z(_03343__PTR23) );
  MUX2_X1 U26046 ( .A(_03342__PTR24), .B(_03342__PTR152), .S(P3_P1_State2_PTR2), .Z(_03343__PTR24) );
  MUX2_X1 U26047 ( .A(_03342__PTR25), .B(_03342__PTR153), .S(P3_P1_State2_PTR2), .Z(_03343__PTR25) );
  MUX2_X1 U26048 ( .A(_03342__PTR26), .B(_03342__PTR154), .S(P3_P1_State2_PTR2), .Z(_03343__PTR26) );
  MUX2_X1 U26049 ( .A(_03342__PTR27), .B(_03342__PTR155), .S(P3_P1_State2_PTR2), .Z(_03343__PTR27) );
  MUX2_X1 U26050 ( .A(_03342__PTR28), .B(_03342__PTR156), .S(P3_P1_State2_PTR2), .Z(_03343__PTR28) );
  MUX2_X1 U26051 ( .A(_03342__PTR29), .B(_03342__PTR157), .S(P3_P1_State2_PTR2), .Z(_03343__PTR29) );
  MUX2_X1 U26052 ( .A(_03342__PTR30), .B(_03342__PTR158), .S(P3_P1_State2_PTR2), .Z(_03343__PTR30) );
  MUX2_X1 U26053 ( .A(_03342__PTR31), .B(_03342__PTR159), .S(P3_P1_State2_PTR2), .Z(_03343__PTR31) );
  MUX2_X1 U26054 ( .A(_03341__PTR0), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR0) );
  MUX2_X1 U26055 ( .A(_03341__PTR1), .B(_03341__PTR65), .S(P3_P1_State2_PTR1), .Z(_03342__PTR1) );
  MUX2_X1 U26056 ( .A(_03341__PTR2), .B(_03341__PTR66), .S(P3_P1_State2_PTR1), .Z(_03342__PTR2) );
  MUX2_X1 U26057 ( .A(_03341__PTR3), .B(_03341__PTR67), .S(P3_P1_State2_PTR1), .Z(_03342__PTR3) );
  MUX2_X1 U26058 ( .A(_03341__PTR4), .B(_03341__PTR68), .S(P3_P1_State2_PTR1), .Z(_03342__PTR4) );
  MUX2_X1 U26059 ( .A(_03341__PTR5), .B(_03341__PTR69), .S(P3_P1_State2_PTR1), .Z(_03342__PTR5) );
  MUX2_X1 U26060 ( .A(_03341__PTR6), .B(_03341__PTR70), .S(P3_P1_State2_PTR1), .Z(_03342__PTR6) );
  MUX2_X1 U26061 ( .A(_03341__PTR7), .B(_03341__PTR71), .S(P3_P1_State2_PTR1), .Z(_03342__PTR7) );
  MUX2_X1 U26062 ( .A(_03341__PTR8), .B(_03341__PTR72), .S(P3_P1_State2_PTR1), .Z(_03342__PTR8) );
  MUX2_X1 U26063 ( .A(_03341__PTR9), .B(_03341__PTR73), .S(P3_P1_State2_PTR1), .Z(_03342__PTR9) );
  MUX2_X1 U26064 ( .A(_03341__PTR10), .B(_03341__PTR74), .S(P3_P1_State2_PTR1), .Z(_03342__PTR10) );
  MUX2_X1 U26065 ( .A(_03341__PTR11), .B(_03341__PTR75), .S(P3_P1_State2_PTR1), .Z(_03342__PTR11) );
  MUX2_X1 U26066 ( .A(_03341__PTR12), .B(_03341__PTR76), .S(P3_P1_State2_PTR1), .Z(_03342__PTR12) );
  MUX2_X1 U26067 ( .A(_03341__PTR13), .B(_03341__PTR77), .S(P3_P1_State2_PTR1), .Z(_03342__PTR13) );
  MUX2_X1 U26068 ( .A(_03341__PTR14), .B(_03341__PTR78), .S(P3_P1_State2_PTR1), .Z(_03342__PTR14) );
  MUX2_X1 U26069 ( .A(_03341__PTR15), .B(_03341__PTR79), .S(P3_P1_State2_PTR1), .Z(_03342__PTR15) );
  MUX2_X1 U26070 ( .A(_03341__PTR16), .B(_03341__PTR80), .S(P3_P1_State2_PTR1), .Z(_03342__PTR16) );
  MUX2_X1 U26071 ( .A(_03341__PTR17), .B(_03341__PTR81), .S(P3_P1_State2_PTR1), .Z(_03342__PTR17) );
  MUX2_X1 U26072 ( .A(_03341__PTR18), .B(_03341__PTR82), .S(P3_P1_State2_PTR1), .Z(_03342__PTR18) );
  MUX2_X1 U26073 ( .A(_03341__PTR19), .B(_03341__PTR83), .S(P3_P1_State2_PTR1), .Z(_03342__PTR19) );
  MUX2_X1 U26074 ( .A(_03341__PTR20), .B(_03341__PTR84), .S(P3_P1_State2_PTR1), .Z(_03342__PTR20) );
  MUX2_X1 U26075 ( .A(_03341__PTR21), .B(_03341__PTR85), .S(P3_P1_State2_PTR1), .Z(_03342__PTR21) );
  MUX2_X1 U26076 ( .A(_03341__PTR22), .B(_03341__PTR86), .S(P3_P1_State2_PTR1), .Z(_03342__PTR22) );
  MUX2_X1 U26077 ( .A(_03341__PTR23), .B(_03341__PTR87), .S(P3_P1_State2_PTR1), .Z(_03342__PTR23) );
  MUX2_X1 U26078 ( .A(_03341__PTR24), .B(_03341__PTR88), .S(P3_P1_State2_PTR1), .Z(_03342__PTR24) );
  MUX2_X1 U26079 ( .A(_03341__PTR25), .B(_03341__PTR89), .S(P3_P1_State2_PTR1), .Z(_03342__PTR25) );
  MUX2_X1 U26080 ( .A(_03341__PTR26), .B(_03341__PTR90), .S(P3_P1_State2_PTR1), .Z(_03342__PTR26) );
  MUX2_X1 U26081 ( .A(_03341__PTR27), .B(_03341__PTR91), .S(P3_P1_State2_PTR1), .Z(_03342__PTR27) );
  MUX2_X1 U26082 ( .A(_03341__PTR28), .B(_03341__PTR92), .S(P3_P1_State2_PTR1), .Z(_03342__PTR28) );
  MUX2_X1 U26083 ( .A(_03341__PTR29), .B(_03341__PTR93), .S(P3_P1_State2_PTR1), .Z(_03342__PTR29) );
  MUX2_X1 U26084 ( .A(_03341__PTR30), .B(_03341__PTR94), .S(P3_P1_State2_PTR1), .Z(_03342__PTR30) );
  MUX2_X1 U26085 ( .A(_03341__PTR31), .B(_03341__PTR95), .S(P3_P1_State2_PTR1), .Z(_03342__PTR31) );
  MUX2_X1 U26086 ( .A(_03341__PTR128), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR128) );
  MUX2_X1 U26087 ( .A(_03341__PTR129), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR129) );
  MUX2_X1 U26088 ( .A(_03341__PTR130), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR130) );
  MUX2_X1 U26089 ( .A(_03341__PTR131), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR131) );
  MUX2_X1 U26090 ( .A(_03341__PTR132), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR132) );
  MUX2_X1 U26091 ( .A(_03341__PTR133), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR133) );
  MUX2_X1 U26092 ( .A(_03341__PTR134), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR134) );
  MUX2_X1 U26093 ( .A(_03341__PTR135), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR135) );
  MUX2_X1 U26094 ( .A(_03341__PTR136), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR136) );
  MUX2_X1 U26095 ( .A(_03341__PTR137), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR137) );
  MUX2_X1 U26096 ( .A(_03341__PTR138), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR138) );
  MUX2_X1 U26097 ( .A(_03341__PTR139), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR139) );
  MUX2_X1 U26098 ( .A(_03341__PTR140), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR140) );
  MUX2_X1 U26099 ( .A(_03341__PTR141), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR141) );
  MUX2_X1 U26100 ( .A(_03341__PTR142), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR142) );
  MUX2_X1 U26101 ( .A(_03341__PTR143), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR143) );
  MUX2_X1 U26102 ( .A(_03341__PTR144), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR144) );
  MUX2_X1 U26103 ( .A(_03341__PTR145), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR145) );
  MUX2_X1 U26104 ( .A(_03341__PTR146), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR146) );
  MUX2_X1 U26105 ( .A(_03341__PTR147), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR147) );
  MUX2_X1 U26106 ( .A(_03341__PTR148), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR148) );
  MUX2_X1 U26107 ( .A(_03341__PTR149), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR149) );
  MUX2_X1 U26108 ( .A(_03341__PTR150), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR150) );
  MUX2_X1 U26109 ( .A(_03341__PTR151), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR151) );
  MUX2_X1 U26110 ( .A(_03341__PTR152), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR152) );
  MUX2_X1 U26111 ( .A(_03341__PTR153), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR153) );
  MUX2_X1 U26112 ( .A(_03341__PTR154), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR154) );
  MUX2_X1 U26113 ( .A(_03341__PTR155), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR155) );
  MUX2_X1 U26114 ( .A(_03341__PTR156), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR156) );
  MUX2_X1 U26115 ( .A(_03341__PTR157), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR157) );
  MUX2_X1 U26116 ( .A(_03341__PTR158), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR158) );
  MUX2_X1 U26117 ( .A(_03341__PTR159), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03342__PTR159) );
  MUX2_X1 U26118 ( .A(P3_rEIP_PTR0), .B(P3_P1_PhyAddrPointer_PTR0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR0) );
  MUX2_X1 U26119 ( .A(P3_rEIP_PTR1), .B(P3_P1_PhyAddrPointer_PTR1), .S(P3_P1_State2_PTR0), .Z(_03341__PTR1) );
  MUX2_X1 U26120 ( .A(P3_rEIP_PTR2), .B(P3_P1_PhyAddrPointer_PTR2), .S(P3_P1_State2_PTR0), .Z(_03341__PTR2) );
  MUX2_X1 U26121 ( .A(P3_rEIP_PTR3), .B(P3_P1_PhyAddrPointer_PTR3), .S(P3_P1_State2_PTR0), .Z(_03341__PTR3) );
  MUX2_X1 U26122 ( .A(P3_rEIP_PTR4), .B(P3_P1_PhyAddrPointer_PTR4), .S(P3_P1_State2_PTR0), .Z(_03341__PTR4) );
  MUX2_X1 U26123 ( .A(P3_rEIP_PTR5), .B(P3_P1_PhyAddrPointer_PTR5), .S(P3_P1_State2_PTR0), .Z(_03341__PTR5) );
  MUX2_X1 U26124 ( .A(P3_rEIP_PTR6), .B(P3_P1_PhyAddrPointer_PTR6), .S(P3_P1_State2_PTR0), .Z(_03341__PTR6) );
  MUX2_X1 U26125 ( .A(P3_rEIP_PTR7), .B(P3_P1_PhyAddrPointer_PTR7), .S(P3_P1_State2_PTR0), .Z(_03341__PTR7) );
  MUX2_X1 U26126 ( .A(P3_rEIP_PTR8), .B(P3_P1_PhyAddrPointer_PTR8), .S(P3_P1_State2_PTR0), .Z(_03341__PTR8) );
  MUX2_X1 U26127 ( .A(P3_rEIP_PTR9), .B(P3_P1_PhyAddrPointer_PTR9), .S(P3_P1_State2_PTR0), .Z(_03341__PTR9) );
  MUX2_X1 U26128 ( .A(P3_rEIP_PTR10), .B(P3_P1_PhyAddrPointer_PTR10), .S(P3_P1_State2_PTR0), .Z(_03341__PTR10) );
  MUX2_X1 U26129 ( .A(P3_rEIP_PTR11), .B(P3_P1_PhyAddrPointer_PTR11), .S(P3_P1_State2_PTR0), .Z(_03341__PTR11) );
  MUX2_X1 U26130 ( .A(P3_rEIP_PTR12), .B(P3_P1_PhyAddrPointer_PTR12), .S(P3_P1_State2_PTR0), .Z(_03341__PTR12) );
  MUX2_X1 U26131 ( .A(P3_rEIP_PTR13), .B(P3_P1_PhyAddrPointer_PTR13), .S(P3_P1_State2_PTR0), .Z(_03341__PTR13) );
  MUX2_X1 U26132 ( .A(P3_rEIP_PTR14), .B(P3_P1_PhyAddrPointer_PTR14), .S(P3_P1_State2_PTR0), .Z(_03341__PTR14) );
  MUX2_X1 U26133 ( .A(P3_rEIP_PTR15), .B(P3_P1_PhyAddrPointer_PTR15), .S(P3_P1_State2_PTR0), .Z(_03341__PTR15) );
  MUX2_X1 U26134 ( .A(P3_rEIP_PTR16), .B(P3_P1_PhyAddrPointer_PTR16), .S(P3_P1_State2_PTR0), .Z(_03341__PTR16) );
  MUX2_X1 U26135 ( .A(P3_rEIP_PTR17), .B(P3_P1_PhyAddrPointer_PTR17), .S(P3_P1_State2_PTR0), .Z(_03341__PTR17) );
  MUX2_X1 U26136 ( .A(P3_rEIP_PTR18), .B(P3_P1_PhyAddrPointer_PTR18), .S(P3_P1_State2_PTR0), .Z(_03341__PTR18) );
  MUX2_X1 U26137 ( .A(P3_rEIP_PTR19), .B(P3_P1_PhyAddrPointer_PTR19), .S(P3_P1_State2_PTR0), .Z(_03341__PTR19) );
  MUX2_X1 U26138 ( .A(P3_rEIP_PTR20), .B(P3_P1_PhyAddrPointer_PTR20), .S(P3_P1_State2_PTR0), .Z(_03341__PTR20) );
  MUX2_X1 U26139 ( .A(P3_rEIP_PTR21), .B(P3_P1_PhyAddrPointer_PTR21), .S(P3_P1_State2_PTR0), .Z(_03341__PTR21) );
  MUX2_X1 U26140 ( .A(P3_rEIP_PTR22), .B(P3_P1_PhyAddrPointer_PTR22), .S(P3_P1_State2_PTR0), .Z(_03341__PTR22) );
  MUX2_X1 U26141 ( .A(P3_rEIP_PTR23), .B(P3_P1_PhyAddrPointer_PTR23), .S(P3_P1_State2_PTR0), .Z(_03341__PTR23) );
  MUX2_X1 U26142 ( .A(P3_rEIP_PTR24), .B(P3_P1_PhyAddrPointer_PTR24), .S(P3_P1_State2_PTR0), .Z(_03341__PTR24) );
  MUX2_X1 U26143 ( .A(P3_rEIP_PTR25), .B(P3_P1_PhyAddrPointer_PTR25), .S(P3_P1_State2_PTR0), .Z(_03341__PTR25) );
  MUX2_X1 U26144 ( .A(P3_rEIP_PTR26), .B(P3_P1_PhyAddrPointer_PTR26), .S(P3_P1_State2_PTR0), .Z(_03341__PTR26) );
  MUX2_X1 U26145 ( .A(P3_rEIP_PTR27), .B(P3_P1_PhyAddrPointer_PTR27), .S(P3_P1_State2_PTR0), .Z(_03341__PTR27) );
  MUX2_X1 U26146 ( .A(P3_rEIP_PTR28), .B(P3_P1_PhyAddrPointer_PTR28), .S(P3_P1_State2_PTR0), .Z(_03341__PTR28) );
  MUX2_X1 U26147 ( .A(P3_rEIP_PTR29), .B(P3_P1_PhyAddrPointer_PTR29), .S(P3_P1_State2_PTR0), .Z(_03341__PTR29) );
  MUX2_X1 U26148 ( .A(P3_rEIP_PTR30), .B(P3_P1_PhyAddrPointer_PTR30), .S(P3_P1_State2_PTR0), .Z(_03341__PTR30) );
  MUX2_X1 U26149 ( .A(P3_rEIP_PTR31), .B(P3_P1_PhyAddrPointer_PTR31), .S(P3_P1_State2_PTR0), .Z(_03341__PTR31) );
  MUX2_X1 U26150 ( .A(_02473__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR65) );
  MUX2_X1 U26151 ( .A(_02473__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR66) );
  MUX2_X1 U26152 ( .A(_02473__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR67) );
  MUX2_X1 U26153 ( .A(_02473__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR68) );
  MUX2_X1 U26154 ( .A(_02473__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR69) );
  MUX2_X1 U26155 ( .A(_02473__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR70) );
  MUX2_X1 U26156 ( .A(_02473__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR71) );
  MUX2_X1 U26157 ( .A(_02473__PTR72), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR72) );
  MUX2_X1 U26158 ( .A(_02473__PTR73), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR73) );
  MUX2_X1 U26159 ( .A(_02473__PTR74), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR74) );
  MUX2_X1 U26160 ( .A(_02473__PTR75), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR75) );
  MUX2_X1 U26161 ( .A(_02473__PTR76), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR76) );
  MUX2_X1 U26162 ( .A(_02473__PTR77), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR77) );
  MUX2_X1 U26163 ( .A(_02473__PTR78), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR78) );
  MUX2_X1 U26164 ( .A(_02473__PTR79), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR79) );
  MUX2_X1 U26165 ( .A(_02473__PTR80), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR80) );
  MUX2_X1 U26166 ( .A(_02473__PTR81), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR81) );
  MUX2_X1 U26167 ( .A(_02473__PTR82), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR82) );
  MUX2_X1 U26168 ( .A(_02473__PTR83), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR83) );
  MUX2_X1 U26169 ( .A(_02473__PTR84), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR84) );
  MUX2_X1 U26170 ( .A(_02473__PTR85), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR85) );
  MUX2_X1 U26171 ( .A(_02473__PTR86), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR86) );
  MUX2_X1 U26172 ( .A(_02473__PTR87), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR87) );
  MUX2_X1 U26173 ( .A(_02473__PTR88), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR88) );
  MUX2_X1 U26174 ( .A(_02473__PTR89), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR89) );
  MUX2_X1 U26175 ( .A(_02473__PTR90), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR90) );
  MUX2_X1 U26176 ( .A(_02473__PTR91), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR91) );
  MUX2_X1 U26177 ( .A(_02473__PTR92), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR92) );
  MUX2_X1 U26178 ( .A(_02473__PTR93), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR93) );
  MUX2_X1 U26179 ( .A(_02473__PTR94), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR94) );
  MUX2_X1 U26180 ( .A(_02473__PTR95), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03341__PTR95) );
  MUX2_X1 U26181 ( .A(1'b0), .B(_02473__PTR160), .S(P3_P1_State2_PTR0), .Z(_03341__PTR128) );
  MUX2_X1 U26182 ( .A(_02473__PTR129), .B(_02473__PTR161), .S(P3_P1_State2_PTR0), .Z(_03341__PTR129) );
  MUX2_X1 U26183 ( .A(_02473__PTR130), .B(_02473__PTR162), .S(P3_P1_State2_PTR0), .Z(_03341__PTR130) );
  MUX2_X1 U26184 ( .A(_02473__PTR131), .B(_02473__PTR163), .S(P3_P1_State2_PTR0), .Z(_03341__PTR131) );
  MUX2_X1 U26185 ( .A(_02473__PTR132), .B(_02473__PTR164), .S(P3_P1_State2_PTR0), .Z(_03341__PTR132) );
  MUX2_X1 U26186 ( .A(_02473__PTR133), .B(_02473__PTR165), .S(P3_P1_State2_PTR0), .Z(_03341__PTR133) );
  MUX2_X1 U26187 ( .A(_02473__PTR134), .B(_02473__PTR166), .S(P3_P1_State2_PTR0), .Z(_03341__PTR134) );
  MUX2_X1 U26188 ( .A(_02473__PTR135), .B(_02473__PTR167), .S(P3_P1_State2_PTR0), .Z(_03341__PTR135) );
  MUX2_X1 U26189 ( .A(_02473__PTR136), .B(_02473__PTR168), .S(P3_P1_State2_PTR0), .Z(_03341__PTR136) );
  MUX2_X1 U26190 ( .A(_02473__PTR137), .B(_02473__PTR169), .S(P3_P1_State2_PTR0), .Z(_03341__PTR137) );
  MUX2_X1 U26191 ( .A(_02473__PTR138), .B(_02473__PTR170), .S(P3_P1_State2_PTR0), .Z(_03341__PTR138) );
  MUX2_X1 U26192 ( .A(_02473__PTR139), .B(_02473__PTR171), .S(P3_P1_State2_PTR0), .Z(_03341__PTR139) );
  MUX2_X1 U26193 ( .A(_02473__PTR140), .B(_02473__PTR172), .S(P3_P1_State2_PTR0), .Z(_03341__PTR140) );
  MUX2_X1 U26194 ( .A(_02473__PTR141), .B(_02473__PTR173), .S(P3_P1_State2_PTR0), .Z(_03341__PTR141) );
  MUX2_X1 U26195 ( .A(_02473__PTR142), .B(_02473__PTR174), .S(P3_P1_State2_PTR0), .Z(_03341__PTR142) );
  MUX2_X1 U26196 ( .A(_02473__PTR143), .B(_02473__PTR175), .S(P3_P1_State2_PTR0), .Z(_03341__PTR143) );
  MUX2_X1 U26197 ( .A(_02473__PTR144), .B(_02473__PTR176), .S(P3_P1_State2_PTR0), .Z(_03341__PTR144) );
  MUX2_X1 U26198 ( .A(_02473__PTR145), .B(_02473__PTR177), .S(P3_P1_State2_PTR0), .Z(_03341__PTR145) );
  MUX2_X1 U26199 ( .A(_02473__PTR146), .B(_02473__PTR178), .S(P3_P1_State2_PTR0), .Z(_03341__PTR146) );
  MUX2_X1 U26200 ( .A(_02473__PTR147), .B(_02473__PTR179), .S(P3_P1_State2_PTR0), .Z(_03341__PTR147) );
  MUX2_X1 U26201 ( .A(_02473__PTR148), .B(_02473__PTR180), .S(P3_P1_State2_PTR0), .Z(_03341__PTR148) );
  MUX2_X1 U26202 ( .A(_02473__PTR149), .B(_02473__PTR181), .S(P3_P1_State2_PTR0), .Z(_03341__PTR149) );
  MUX2_X1 U26203 ( .A(_02473__PTR150), .B(_02473__PTR182), .S(P3_P1_State2_PTR0), .Z(_03341__PTR150) );
  MUX2_X1 U26204 ( .A(_02473__PTR151), .B(_02473__PTR183), .S(P3_P1_State2_PTR0), .Z(_03341__PTR151) );
  MUX2_X1 U26205 ( .A(_02473__PTR152), .B(_02473__PTR184), .S(P3_P1_State2_PTR0), .Z(_03341__PTR152) );
  MUX2_X1 U26206 ( .A(_02473__PTR153), .B(_02473__PTR185), .S(P3_P1_State2_PTR0), .Z(_03341__PTR153) );
  MUX2_X1 U26207 ( .A(_02473__PTR154), .B(_02473__PTR186), .S(P3_P1_State2_PTR0), .Z(_03341__PTR154) );
  MUX2_X1 U26208 ( .A(_02473__PTR155), .B(_02473__PTR187), .S(P3_P1_State2_PTR0), .Z(_03341__PTR155) );
  MUX2_X1 U26209 ( .A(_02473__PTR156), .B(_02473__PTR188), .S(P3_P1_State2_PTR0), .Z(_03341__PTR156) );
  MUX2_X1 U26210 ( .A(_02473__PTR157), .B(_02473__PTR189), .S(P3_P1_State2_PTR0), .Z(_03341__PTR157) );
  MUX2_X1 U26211 ( .A(_02473__PTR158), .B(_02473__PTR190), .S(P3_P1_State2_PTR0), .Z(_03341__PTR158) );
  MUX2_X1 U26212 ( .A(_02473__PTR159), .B(_02473__PTR191), .S(P3_P1_State2_PTR0), .Z(_03341__PTR159) );
  MUX2_X1 U26213 ( .A(_03345__PTR0), .B(_03345__PTR128), .S(P3_P1_State2_PTR2), .Z(_03346__PTR0) );
  MUX2_X1 U26214 ( .A(_03345__PTR1), .B(_03345__PTR129), .S(P3_P1_State2_PTR2), .Z(_03346__PTR1) );
  MUX2_X1 U26215 ( .A(_03345__PTR2), .B(_03345__PTR130), .S(P3_P1_State2_PTR2), .Z(_03346__PTR2) );
  MUX2_X1 U26216 ( .A(_03345__PTR3), .B(_03345__PTR131), .S(P3_P1_State2_PTR2), .Z(_03346__PTR3) );
  MUX2_X1 U26217 ( .A(_03345__PTR4), .B(_03345__PTR132), .S(P3_P1_State2_PTR2), .Z(_03346__PTR4) );
  MUX2_X1 U26218 ( .A(_03345__PTR5), .B(_03345__PTR133), .S(P3_P1_State2_PTR2), .Z(_03346__PTR5) );
  MUX2_X1 U26219 ( .A(_03345__PTR6), .B(_03345__PTR134), .S(P3_P1_State2_PTR2), .Z(_03346__PTR6) );
  MUX2_X1 U26220 ( .A(_03345__PTR7), .B(_03345__PTR135), .S(P3_P1_State2_PTR2), .Z(_03346__PTR7) );
  MUX2_X1 U26221 ( .A(_03345__PTR8), .B(_03345__PTR136), .S(P3_P1_State2_PTR2), .Z(_03346__PTR8) );
  MUX2_X1 U26222 ( .A(_03345__PTR9), .B(_03345__PTR137), .S(P3_P1_State2_PTR2), .Z(_03346__PTR9) );
  MUX2_X1 U26223 ( .A(_03345__PTR10), .B(_03345__PTR138), .S(P3_P1_State2_PTR2), .Z(_03346__PTR10) );
  MUX2_X1 U26224 ( .A(_03345__PTR11), .B(_03345__PTR139), .S(P3_P1_State2_PTR2), .Z(_03346__PTR11) );
  MUX2_X1 U26225 ( .A(_03345__PTR12), .B(_03345__PTR140), .S(P3_P1_State2_PTR2), .Z(_03346__PTR12) );
  MUX2_X1 U26226 ( .A(_03345__PTR13), .B(_03345__PTR141), .S(P3_P1_State2_PTR2), .Z(_03346__PTR13) );
  MUX2_X1 U26227 ( .A(_03345__PTR14), .B(_03345__PTR142), .S(P3_P1_State2_PTR2), .Z(_03346__PTR14) );
  MUX2_X1 U26228 ( .A(_03345__PTR15), .B(_03345__PTR143), .S(P3_P1_State2_PTR2), .Z(_03346__PTR15) );
  MUX2_X1 U26229 ( .A(_03345__PTR16), .B(_03345__PTR144), .S(P3_P1_State2_PTR2), .Z(_03346__PTR16) );
  MUX2_X1 U26230 ( .A(_03345__PTR17), .B(_03345__PTR145), .S(P3_P1_State2_PTR2), .Z(_03346__PTR17) );
  MUX2_X1 U26231 ( .A(_03345__PTR18), .B(_03345__PTR146), .S(P3_P1_State2_PTR2), .Z(_03346__PTR18) );
  MUX2_X1 U26232 ( .A(_03345__PTR19), .B(_03345__PTR147), .S(P3_P1_State2_PTR2), .Z(_03346__PTR19) );
  MUX2_X1 U26233 ( .A(_03345__PTR20), .B(_03345__PTR148), .S(P3_P1_State2_PTR2), .Z(_03346__PTR20) );
  MUX2_X1 U26234 ( .A(_03345__PTR21), .B(_03345__PTR149), .S(P3_P1_State2_PTR2), .Z(_03346__PTR21) );
  MUX2_X1 U26235 ( .A(_03345__PTR22), .B(_03345__PTR150), .S(P3_P1_State2_PTR2), .Z(_03346__PTR22) );
  MUX2_X1 U26236 ( .A(_03345__PTR23), .B(_03345__PTR151), .S(P3_P1_State2_PTR2), .Z(_03346__PTR23) );
  MUX2_X1 U26237 ( .A(_03345__PTR24), .B(_03345__PTR152), .S(P3_P1_State2_PTR2), .Z(_03346__PTR24) );
  MUX2_X1 U26238 ( .A(_03345__PTR25), .B(_03345__PTR153), .S(P3_P1_State2_PTR2), .Z(_03346__PTR25) );
  MUX2_X1 U26239 ( .A(_03345__PTR26), .B(_03345__PTR154), .S(P3_P1_State2_PTR2), .Z(_03346__PTR26) );
  MUX2_X1 U26240 ( .A(_03345__PTR27), .B(_03345__PTR155), .S(P3_P1_State2_PTR2), .Z(_03346__PTR27) );
  MUX2_X1 U26241 ( .A(_03345__PTR28), .B(_03345__PTR156), .S(P3_P1_State2_PTR2), .Z(_03346__PTR28) );
  MUX2_X1 U26242 ( .A(_03345__PTR29), .B(_03345__PTR157), .S(P3_P1_State2_PTR2), .Z(_03346__PTR29) );
  MUX2_X1 U26243 ( .A(_03345__PTR30), .B(_03345__PTR158), .S(P3_P1_State2_PTR2), .Z(_03346__PTR30) );
  MUX2_X1 U26244 ( .A(_03345__PTR31), .B(_03345__PTR159), .S(P3_P1_State2_PTR2), .Z(_03346__PTR31) );
  MUX2_X1 U26245 ( .A(_03344__PTR0), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR0) );
  MUX2_X1 U26246 ( .A(_03344__PTR1), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR1) );
  MUX2_X1 U26247 ( .A(_03344__PTR2), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR2) );
  MUX2_X1 U26248 ( .A(_03344__PTR3), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR3) );
  MUX2_X1 U26249 ( .A(_03344__PTR4), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR4) );
  MUX2_X1 U26250 ( .A(_03344__PTR5), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR5) );
  MUX2_X1 U26251 ( .A(_03344__PTR6), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR6) );
  MUX2_X1 U26252 ( .A(_03344__PTR7), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR7) );
  MUX2_X1 U26253 ( .A(_03344__PTR8), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR8) );
  MUX2_X1 U26254 ( .A(_03344__PTR9), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR9) );
  MUX2_X1 U26255 ( .A(_03344__PTR10), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR10) );
  MUX2_X1 U26256 ( .A(_03344__PTR11), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR11) );
  MUX2_X1 U26257 ( .A(_03344__PTR12), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR12) );
  MUX2_X1 U26258 ( .A(_03344__PTR13), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR13) );
  MUX2_X1 U26259 ( .A(_03344__PTR14), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR14) );
  MUX2_X1 U26260 ( .A(_03344__PTR15), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR15) );
  MUX2_X1 U26261 ( .A(_03344__PTR16), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR16) );
  MUX2_X1 U26262 ( .A(_03344__PTR17), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR17) );
  MUX2_X1 U26263 ( .A(_03344__PTR18), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR18) );
  MUX2_X1 U26264 ( .A(_03344__PTR19), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR19) );
  MUX2_X1 U26265 ( .A(_03344__PTR20), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR20) );
  MUX2_X1 U26266 ( .A(_03344__PTR21), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR21) );
  MUX2_X1 U26267 ( .A(_03344__PTR22), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR22) );
  MUX2_X1 U26268 ( .A(_03344__PTR23), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR23) );
  MUX2_X1 U26269 ( .A(_03344__PTR24), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR24) );
  MUX2_X1 U26270 ( .A(_03344__PTR25), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR25) );
  MUX2_X1 U26271 ( .A(_03344__PTR26), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR26) );
  MUX2_X1 U26272 ( .A(_03344__PTR27), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR27) );
  MUX2_X1 U26273 ( .A(_03344__PTR28), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR28) );
  MUX2_X1 U26274 ( .A(_03344__PTR29), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR29) );
  MUX2_X1 U26275 ( .A(_03344__PTR30), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR30) );
  MUX2_X1 U26276 ( .A(_03344__PTR31), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR31) );
  MUX2_X1 U26277 ( .A(_03344__PTR128), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR128) );
  MUX2_X1 U26278 ( .A(_03344__PTR129), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR129) );
  MUX2_X1 U26279 ( .A(_03344__PTR130), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR130) );
  MUX2_X1 U26280 ( .A(_03344__PTR131), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR131) );
  MUX2_X1 U26281 ( .A(_03344__PTR132), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR132) );
  MUX2_X1 U26282 ( .A(_03344__PTR133), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR133) );
  MUX2_X1 U26283 ( .A(_03344__PTR134), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR134) );
  MUX2_X1 U26284 ( .A(_03344__PTR135), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR135) );
  MUX2_X1 U26285 ( .A(_03344__PTR136), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR136) );
  MUX2_X1 U26286 ( .A(_03344__PTR137), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR137) );
  MUX2_X1 U26287 ( .A(_03344__PTR138), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR138) );
  MUX2_X1 U26288 ( .A(_03344__PTR139), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR139) );
  MUX2_X1 U26289 ( .A(_03344__PTR140), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR140) );
  MUX2_X1 U26290 ( .A(_03344__PTR141), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR141) );
  MUX2_X1 U26291 ( .A(_03344__PTR142), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR142) );
  MUX2_X1 U26292 ( .A(_03344__PTR143), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR143) );
  MUX2_X1 U26293 ( .A(_03344__PTR144), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR144) );
  MUX2_X1 U26294 ( .A(_03344__PTR145), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR145) );
  MUX2_X1 U26295 ( .A(_03344__PTR146), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR146) );
  MUX2_X1 U26296 ( .A(_03344__PTR147), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR147) );
  MUX2_X1 U26297 ( .A(_03344__PTR148), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR148) );
  MUX2_X1 U26298 ( .A(_03344__PTR149), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR149) );
  MUX2_X1 U26299 ( .A(_03344__PTR150), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR150) );
  MUX2_X1 U26300 ( .A(_03344__PTR151), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR151) );
  MUX2_X1 U26301 ( .A(_03344__PTR152), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR152) );
  MUX2_X1 U26302 ( .A(_03344__PTR153), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR153) );
  MUX2_X1 U26303 ( .A(_03344__PTR154), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR154) );
  MUX2_X1 U26304 ( .A(_03344__PTR155), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR155) );
  MUX2_X1 U26305 ( .A(_03344__PTR156), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR156) );
  MUX2_X1 U26306 ( .A(_03344__PTR157), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR157) );
  MUX2_X1 U26307 ( .A(_03344__PTR158), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR158) );
  MUX2_X1 U26308 ( .A(_03344__PTR159), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03345__PTR159) );
  MUX2_X1 U26309 ( .A(P3_rEIP_PTR0), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR0) );
  MUX2_X1 U26310 ( .A(P3_rEIP_PTR1), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR1) );
  MUX2_X1 U26311 ( .A(P3_rEIP_PTR2), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR2) );
  MUX2_X1 U26312 ( .A(P3_rEIP_PTR3), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR3) );
  MUX2_X1 U26313 ( .A(P3_rEIP_PTR4), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR4) );
  MUX2_X1 U26314 ( .A(P3_rEIP_PTR5), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR5) );
  MUX2_X1 U26315 ( .A(P3_rEIP_PTR6), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR6) );
  MUX2_X1 U26316 ( .A(P3_rEIP_PTR7), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR7) );
  MUX2_X1 U26317 ( .A(P3_rEIP_PTR8), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR8) );
  MUX2_X1 U26318 ( .A(P3_rEIP_PTR9), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR9) );
  MUX2_X1 U26319 ( .A(P3_rEIP_PTR10), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR10) );
  MUX2_X1 U26320 ( .A(P3_rEIP_PTR11), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR11) );
  MUX2_X1 U26321 ( .A(P3_rEIP_PTR12), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR12) );
  MUX2_X1 U26322 ( .A(P3_rEIP_PTR13), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR13) );
  MUX2_X1 U26323 ( .A(P3_rEIP_PTR14), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR14) );
  MUX2_X1 U26324 ( .A(P3_rEIP_PTR15), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR15) );
  MUX2_X1 U26325 ( .A(P3_rEIP_PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR16) );
  MUX2_X1 U26326 ( .A(P3_rEIP_PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR17) );
  MUX2_X1 U26327 ( .A(P3_rEIP_PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR18) );
  MUX2_X1 U26328 ( .A(P3_rEIP_PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR19) );
  MUX2_X1 U26329 ( .A(P3_rEIP_PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR20) );
  MUX2_X1 U26330 ( .A(P3_rEIP_PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR21) );
  MUX2_X1 U26331 ( .A(P3_rEIP_PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR22) );
  MUX2_X1 U26332 ( .A(P3_rEIP_PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR23) );
  MUX2_X1 U26333 ( .A(P3_rEIP_PTR24), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR24) );
  MUX2_X1 U26334 ( .A(P3_rEIP_PTR25), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR25) );
  MUX2_X1 U26335 ( .A(P3_rEIP_PTR26), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR26) );
  MUX2_X1 U26336 ( .A(P3_rEIP_PTR27), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR27) );
  MUX2_X1 U26337 ( .A(P3_rEIP_PTR28), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR28) );
  MUX2_X1 U26338 ( .A(P3_rEIP_PTR29), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR29) );
  MUX2_X1 U26339 ( .A(P3_rEIP_PTR30), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR30) );
  MUX2_X1 U26340 ( .A(P3_rEIP_PTR31), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03344__PTR31) );
  MUX2_X1 U26341 ( .A(1'b0), .B(_02474__PTR160), .S(P3_P1_State2_PTR0), .Z(_03344__PTR128) );
  MUX2_X1 U26342 ( .A(1'b0), .B(_02474__PTR161), .S(P3_P1_State2_PTR0), .Z(_03344__PTR129) );
  MUX2_X1 U26343 ( .A(1'b0), .B(_02474__PTR162), .S(P3_P1_State2_PTR0), .Z(_03344__PTR130) );
  MUX2_X1 U26344 ( .A(1'b0), .B(_02474__PTR163), .S(P3_P1_State2_PTR0), .Z(_03344__PTR131) );
  MUX2_X1 U26345 ( .A(1'b0), .B(_02474__PTR164), .S(P3_P1_State2_PTR0), .Z(_03344__PTR132) );
  MUX2_X1 U26346 ( .A(1'b0), .B(_02474__PTR165), .S(P3_P1_State2_PTR0), .Z(_03344__PTR133) );
  MUX2_X1 U26347 ( .A(1'b0), .B(_02474__PTR166), .S(P3_P1_State2_PTR0), .Z(_03344__PTR134) );
  MUX2_X1 U26348 ( .A(1'b0), .B(_02474__PTR167), .S(P3_P1_State2_PTR0), .Z(_03344__PTR135) );
  MUX2_X1 U26349 ( .A(1'b0), .B(_02474__PTR168), .S(P3_P1_State2_PTR0), .Z(_03344__PTR136) );
  MUX2_X1 U26350 ( .A(1'b0), .B(_02474__PTR169), .S(P3_P1_State2_PTR0), .Z(_03344__PTR137) );
  MUX2_X1 U26351 ( .A(1'b0), .B(_02474__PTR170), .S(P3_P1_State2_PTR0), .Z(_03344__PTR138) );
  MUX2_X1 U26352 ( .A(1'b0), .B(_02474__PTR171), .S(P3_P1_State2_PTR0), .Z(_03344__PTR139) );
  MUX2_X1 U26353 ( .A(1'b0), .B(_02474__PTR172), .S(P3_P1_State2_PTR0), .Z(_03344__PTR140) );
  MUX2_X1 U26354 ( .A(1'b0), .B(_02474__PTR173), .S(P3_P1_State2_PTR0), .Z(_03344__PTR141) );
  MUX2_X1 U26355 ( .A(1'b0), .B(_02474__PTR174), .S(P3_P1_State2_PTR0), .Z(_03344__PTR142) );
  MUX2_X1 U26356 ( .A(1'b0), .B(_02474__PTR175), .S(P3_P1_State2_PTR0), .Z(_03344__PTR143) );
  MUX2_X1 U26357 ( .A(1'b0), .B(_02474__PTR176), .S(P3_P1_State2_PTR0), .Z(_03344__PTR144) );
  MUX2_X1 U26358 ( .A(1'b0), .B(_02474__PTR177), .S(P3_P1_State2_PTR0), .Z(_03344__PTR145) );
  MUX2_X1 U26359 ( .A(1'b0), .B(_02474__PTR178), .S(P3_P1_State2_PTR0), .Z(_03344__PTR146) );
  MUX2_X1 U26360 ( .A(1'b0), .B(_02474__PTR179), .S(P3_P1_State2_PTR0), .Z(_03344__PTR147) );
  MUX2_X1 U26361 ( .A(1'b0), .B(_02474__PTR180), .S(P3_P1_State2_PTR0), .Z(_03344__PTR148) );
  MUX2_X1 U26362 ( .A(1'b0), .B(_02474__PTR181), .S(P3_P1_State2_PTR0), .Z(_03344__PTR149) );
  MUX2_X1 U26363 ( .A(1'b0), .B(_02474__PTR182), .S(P3_P1_State2_PTR0), .Z(_03344__PTR150) );
  MUX2_X1 U26364 ( .A(1'b0), .B(_02474__PTR183), .S(P3_P1_State2_PTR0), .Z(_03344__PTR151) );
  MUX2_X1 U26365 ( .A(1'b0), .B(_02474__PTR184), .S(P3_P1_State2_PTR0), .Z(_03344__PTR152) );
  MUX2_X1 U26366 ( .A(1'b0), .B(_02474__PTR185), .S(P3_P1_State2_PTR0), .Z(_03344__PTR153) );
  MUX2_X1 U26367 ( .A(1'b0), .B(_02474__PTR186), .S(P3_P1_State2_PTR0), .Z(_03344__PTR154) );
  MUX2_X1 U26368 ( .A(1'b0), .B(_02474__PTR187), .S(P3_P1_State2_PTR0), .Z(_03344__PTR155) );
  MUX2_X1 U26369 ( .A(1'b0), .B(_02474__PTR188), .S(P3_P1_State2_PTR0), .Z(_03344__PTR156) );
  MUX2_X1 U26370 ( .A(1'b0), .B(_02474__PTR189), .S(P3_P1_State2_PTR0), .Z(_03344__PTR157) );
  MUX2_X1 U26371 ( .A(1'b0), .B(_02474__PTR190), .S(P3_P1_State2_PTR0), .Z(_03344__PTR158) );
  MUX2_X1 U26372 ( .A(1'b0), .B(_02474__PTR191), .S(P3_P1_State2_PTR0), .Z(_03344__PTR159) );
  MUX2_X1 U26373 ( .A(_03349__PTR0), .B(_03347__PTR32), .S(P3_P1_State2_PTR3), .Z(_02476__PTR0) );
  MUX2_X1 U26374 ( .A(_03349__PTR1), .B(1'b0), .S(P3_P1_State2_PTR3), .Z(_02476__PTR1) );
  MUX2_X1 U26375 ( .A(_03349__PTR2), .B(1'b0), .S(P3_P1_State2_PTR3), .Z(_02476__PTR2) );
  MUX2_X1 U26376 ( .A(_03349__PTR3), .B(_00298_), .S(P3_P1_State2_PTR3), .Z(_02476__PTR3) );
  MUX2_X1 U26377 ( .A(_03347__PTR0), .B(_03347__PTR16), .S(P3_P1_State2_PTR2), .Z(_03349__PTR0) );
  MUX2_X1 U26378 ( .A(_03347__PTR1), .B(_03347__PTR17), .S(P3_P1_State2_PTR2), .Z(_03349__PTR1) );
  MUX2_X1 U26379 ( .A(_03347__PTR2), .B(_03347__PTR18), .S(P3_P1_State2_PTR2), .Z(_03349__PTR2) );
  MUX2_X1 U26380 ( .A(1'b0), .B(_03347__PTR19), .S(P3_P1_State2_PTR2), .Z(_03349__PTR3) );
  MUX2_X1 U26381 ( .A(_03350__PTR1), .B(_03348__PTR1), .S(P3_P1_State2_PTR1), .Z(_03347__PTR1) );
  MUX2_X1 U26382 ( .A(1'b0), .B(_03348__PTR2), .S(P3_P1_State2_PTR1), .Z(_03347__PTR2) );
  MUX2_X1 U26383 ( .A(_03348__PTR8), .B(_03348__PTR16), .S(P3_P1_State2_PTR1), .Z(_03347__PTR16) );
  MUX2_X1 U26384 ( .A(_03348__PTR9), .B(_03348__PTR17), .S(P3_P1_State2_PTR1), .Z(_03347__PTR17) );
  MUX2_X1 U26385 ( .A(_03348__PTR10), .B(_03348__PTR18), .S(P3_P1_State2_PTR1), .Z(_03347__PTR18) );
  MUX2_X1 U26386 ( .A(_03348__PTR11), .B(_03348__PTR19), .S(P3_P1_State2_PTR1), .Z(_03347__PTR19) );
  MUX2_X1 U26387 ( .A(1'b0), .B(_02475__PTR14), .S(P3_P1_State2_PTR0), .Z(_03350__PTR1) );
  MUX2_X1 U26388 ( .A(1'b1), .B(P3_READY_n), .S(P3_P1_State2_PTR0), .Z(_03347__PTR0) );
  MUX2_X1 U26389 ( .A(_02475__PTR9), .B(P3_READY_n), .S(P3_P1_State2_PTR0), .Z(_03348__PTR1) );
  MUX2_X1 U26390 ( .A(P3_StateBS16), .B(_02475__PTR14), .S(P3_P1_State2_PTR0), .Z(_03348__PTR2) );
  MUX2_X1 U26391 ( .A(1'b1), .B(_02475__PTR20), .S(P3_P1_State2_PTR0), .Z(_03348__PTR8) );
  MUX2_X1 U26392 ( .A(1'b0), .B(_02475__PTR21), .S(P3_P1_State2_PTR0), .Z(_03348__PTR9) );
  MUX2_X1 U26393 ( .A(1'b1), .B(_02475__PTR22), .S(P3_P1_State2_PTR0), .Z(_03348__PTR10) );
  MUX2_X1 U26394 ( .A(1'b0), .B(_02475__PTR23), .S(P3_P1_State2_PTR0), .Z(_03348__PTR11) );
  MUX2_X1 U26395 ( .A(_02475__PTR26), .B(_02475__PTR28), .S(P3_P1_State2_PTR0), .Z(_03348__PTR16) );
  MUX2_X1 U26396 ( .A(_02431__PTR6), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03348__PTR17) );
  MUX2_X1 U26397 ( .A(_02475__PTR26), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03348__PTR18) );
  MUX2_X1 U26398 ( .A(_02431__PTR6), .B(1'b1), .S(P3_P1_State2_PTR0), .Z(_03348__PTR19) );
  MUX2_X1 U26399 ( .A(_02475__PTR32), .B(1'b1), .S(P3_P1_State2_PTR0), .Z(_03347__PTR32) );
  MUX2_X1 U26400 ( .A(_03351__PTR32), .B(_03351__PTR128), .S(P3_P1_State2_PTR1), .Z(_03352__PTR0) );
  MUX2_X1 U26401 ( .A(_03351__PTR32), .B(_03351__PTR129), .S(P3_P1_State2_PTR1), .Z(_03352__PTR1) );
  MUX2_X1 U26402 ( .A(_03351__PTR32), .B(_03351__PTR130), .S(P3_P1_State2_PTR1), .Z(_03352__PTR2) );
  MUX2_X1 U26403 ( .A(_03351__PTR32), .B(_03351__PTR131), .S(P3_P1_State2_PTR1), .Z(_03352__PTR3) );
  MUX2_X1 U26404 ( .A(_03351__PTR19), .B(_03351__PTR132), .S(P3_P1_State2_PTR1), .Z(_03352__PTR4) );
  MUX2_X1 U26405 ( .A(_03351__PTR19), .B(_03351__PTR133), .S(P3_P1_State2_PTR1), .Z(_03352__PTR5) );
  MUX2_X1 U26406 ( .A(_03351__PTR19), .B(_03351__PTR134), .S(P3_P1_State2_PTR1), .Z(_03352__PTR6) );
  MUX2_X1 U26407 ( .A(_03351__PTR19), .B(_03351__PTR135), .S(P3_P1_State2_PTR1), .Z(_03352__PTR7) );
  MUX2_X1 U26408 ( .A(_03351__PTR19), .B(_03351__PTR136), .S(P3_P1_State2_PTR1), .Z(_03352__PTR8) );
  MUX2_X1 U26409 ( .A(_03351__PTR19), .B(_03351__PTR137), .S(P3_P1_State2_PTR1), .Z(_03352__PTR9) );
  MUX2_X1 U26410 ( .A(_03351__PTR19), .B(_03351__PTR138), .S(P3_P1_State2_PTR1), .Z(_03352__PTR10) );
  MUX2_X1 U26411 ( .A(_03351__PTR19), .B(_03351__PTR139), .S(P3_P1_State2_PTR1), .Z(_03352__PTR11) );
  MUX2_X1 U26412 ( .A(_03351__PTR19), .B(_03351__PTR140), .S(P3_P1_State2_PTR1), .Z(_03352__PTR12) );
  MUX2_X1 U26413 ( .A(_03351__PTR19), .B(_03351__PTR141), .S(P3_P1_State2_PTR1), .Z(_03352__PTR13) );
  MUX2_X1 U26414 ( .A(_03351__PTR19), .B(_03351__PTR142), .S(P3_P1_State2_PTR1), .Z(_03352__PTR14) );
  MUX2_X1 U26415 ( .A(_03351__PTR19), .B(_03351__PTR143), .S(P3_P1_State2_PTR1), .Z(_03352__PTR15) );
  MUX2_X1 U26416 ( .A(_03351__PTR19), .B(_03351__PTR144), .S(P3_P1_State2_PTR1), .Z(_03352__PTR16) );
  MUX2_X1 U26417 ( .A(_03351__PTR19), .B(_03351__PTR145), .S(P3_P1_State2_PTR1), .Z(_03352__PTR17) );
  MUX2_X1 U26418 ( .A(_03351__PTR19), .B(_03351__PTR146), .S(P3_P1_State2_PTR1), .Z(_03352__PTR18) );
  MUX2_X1 U26419 ( .A(_03351__PTR19), .B(_03351__PTR147), .S(P3_P1_State2_PTR1), .Z(_03352__PTR19) );
  MUX2_X1 U26420 ( .A(_03351__PTR32), .B(_03351__PTR148), .S(P3_P1_State2_PTR1), .Z(_03352__PTR20) );
  MUX2_X1 U26421 ( .A(_03351__PTR32), .B(_03351__PTR149), .S(P3_P1_State2_PTR1), .Z(_03352__PTR21) );
  MUX2_X1 U26422 ( .A(_03351__PTR32), .B(_03351__PTR150), .S(P3_P1_State2_PTR1), .Z(_03352__PTR22) );
  MUX2_X1 U26423 ( .A(_03351__PTR32), .B(_03351__PTR151), .S(P3_P1_State2_PTR1), .Z(_03352__PTR23) );
  MUX2_X1 U26424 ( .A(_03351__PTR32), .B(_03351__PTR152), .S(P3_P1_State2_PTR1), .Z(_03352__PTR24) );
  MUX2_X1 U26425 ( .A(_03351__PTR32), .B(_03351__PTR153), .S(P3_P1_State2_PTR1), .Z(_03352__PTR25) );
  MUX2_X1 U26426 ( .A(_03351__PTR32), .B(_03351__PTR154), .S(P3_P1_State2_PTR1), .Z(_03352__PTR26) );
  MUX2_X1 U26427 ( .A(_03351__PTR32), .B(_03351__PTR155), .S(P3_P1_State2_PTR1), .Z(_03352__PTR27) );
  MUX2_X1 U26428 ( .A(_03351__PTR32), .B(_03351__PTR156), .S(P3_P1_State2_PTR1), .Z(_03352__PTR28) );
  MUX2_X1 U26429 ( .A(_03351__PTR32), .B(_03351__PTR157), .S(P3_P1_State2_PTR1), .Z(_03352__PTR29) );
  MUX2_X1 U26430 ( .A(_03351__PTR32), .B(_03351__PTR158), .S(P3_P1_State2_PTR1), .Z(_03352__PTR30) );
  MUX2_X1 U26431 ( .A(_03351__PTR32), .B(_03351__PTR160), .S(P3_P1_State2_PTR1), .Z(_03352__PTR32) );
  MUX2_X1 U26432 ( .A(_03351__PTR256), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR256) );
  MUX2_X1 U26433 ( .A(_03351__PTR257), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR257) );
  MUX2_X1 U26434 ( .A(_03351__PTR258), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR258) );
  MUX2_X1 U26435 ( .A(_03351__PTR259), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR259) );
  MUX2_X1 U26436 ( .A(_03351__PTR260), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR260) );
  MUX2_X1 U26437 ( .A(_03351__PTR261), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR261) );
  MUX2_X1 U26438 ( .A(_03351__PTR262), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR262) );
  MUX2_X1 U26439 ( .A(_03351__PTR263), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR263) );
  MUX2_X1 U26440 ( .A(_03351__PTR264), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR264) );
  MUX2_X1 U26441 ( .A(_03351__PTR265), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR265) );
  MUX2_X1 U26442 ( .A(_03351__PTR266), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR266) );
  MUX2_X1 U26443 ( .A(_03351__PTR267), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR267) );
  MUX2_X1 U26444 ( .A(_03351__PTR268), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR268) );
  MUX2_X1 U26445 ( .A(_03351__PTR269), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR269) );
  MUX2_X1 U26446 ( .A(_03351__PTR270), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR270) );
  MUX2_X1 U26447 ( .A(_03351__PTR271), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR271) );
  MUX2_X1 U26448 ( .A(_03351__PTR272), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR272) );
  MUX2_X1 U26449 ( .A(_03351__PTR273), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR273) );
  MUX2_X1 U26450 ( .A(_03351__PTR274), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR274) );
  MUX2_X1 U26451 ( .A(_03351__PTR275), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR275) );
  MUX2_X1 U26452 ( .A(_03351__PTR276), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR276) );
  MUX2_X1 U26453 ( .A(_03351__PTR277), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR277) );
  MUX2_X1 U26454 ( .A(_03351__PTR278), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR278) );
  MUX2_X1 U26455 ( .A(_03351__PTR279), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR279) );
  MUX2_X1 U26456 ( .A(_03351__PTR280), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR280) );
  MUX2_X1 U26457 ( .A(_03351__PTR281), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR281) );
  MUX2_X1 U26458 ( .A(_03351__PTR282), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR282) );
  MUX2_X1 U26459 ( .A(_03351__PTR283), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR283) );
  MUX2_X1 U26460 ( .A(_03351__PTR284), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR284) );
  MUX2_X1 U26461 ( .A(_03351__PTR285), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR285) );
  MUX2_X1 U26462 ( .A(_03351__PTR286), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR286) );
  MUX2_X1 U26463 ( .A(_03351__PTR288), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03352__PTR288) );
  MUX2_X1 U26464 ( .A(1'b0), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR32) );
  MUX2_X1 U26465 ( .A(1'b1), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR19) );
  MUX2_X1 U26466 ( .A(_02477__PTR128), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR128) );
  MUX2_X1 U26467 ( .A(_02477__PTR129), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR129) );
  MUX2_X1 U26468 ( .A(_02477__PTR130), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR130) );
  MUX2_X1 U26469 ( .A(_02477__PTR131), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR131) );
  MUX2_X1 U26470 ( .A(_02477__PTR132), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR132) );
  MUX2_X1 U26471 ( .A(_02477__PTR133), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR133) );
  MUX2_X1 U26472 ( .A(_02477__PTR134), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR134) );
  MUX2_X1 U26473 ( .A(_02477__PTR135), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR135) );
  MUX2_X1 U26474 ( .A(_02477__PTR136), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR136) );
  MUX2_X1 U26475 ( .A(_02477__PTR137), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR137) );
  MUX2_X1 U26476 ( .A(_02477__PTR138), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR138) );
  MUX2_X1 U26477 ( .A(_02477__PTR139), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR139) );
  MUX2_X1 U26478 ( .A(_02477__PTR140), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR140) );
  MUX2_X1 U26479 ( .A(_02477__PTR141), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR141) );
  MUX2_X1 U26480 ( .A(_02477__PTR142), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR142) );
  MUX2_X1 U26481 ( .A(_02477__PTR143), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR143) );
  MUX2_X1 U26482 ( .A(_02477__PTR144), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR144) );
  MUX2_X1 U26483 ( .A(_02477__PTR145), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR145) );
  MUX2_X1 U26484 ( .A(_02477__PTR146), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR146) );
  MUX2_X1 U26485 ( .A(_02477__PTR147), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR147) );
  MUX2_X1 U26486 ( .A(_02477__PTR148), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR148) );
  MUX2_X1 U26487 ( .A(_02477__PTR149), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR149) );
  MUX2_X1 U26488 ( .A(_02477__PTR150), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR150) );
  MUX2_X1 U26489 ( .A(_02477__PTR151), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR151) );
  MUX2_X1 U26490 ( .A(_02477__PTR152), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR152) );
  MUX2_X1 U26491 ( .A(_02477__PTR153), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR153) );
  MUX2_X1 U26492 ( .A(_02477__PTR154), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR154) );
  MUX2_X1 U26493 ( .A(_02477__PTR155), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR155) );
  MUX2_X1 U26494 ( .A(_02477__PTR156), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR156) );
  MUX2_X1 U26495 ( .A(_02477__PTR157), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR157) );
  MUX2_X1 U26496 ( .A(_02477__PTR158), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR158) );
  MUX2_X1 U26497 ( .A(_02477__PTR160), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03351__PTR160) );
  MUX2_X1 U26498 ( .A(1'b0), .B(_02477__PTR320), .S(P3_P1_State2_PTR0), .Z(_03351__PTR256) );
  MUX2_X1 U26499 ( .A(1'b0), .B(_02477__PTR321), .S(P3_P1_State2_PTR0), .Z(_03351__PTR257) );
  MUX2_X1 U26500 ( .A(1'b0), .B(_02477__PTR322), .S(P3_P1_State2_PTR0), .Z(_03351__PTR258) );
  MUX2_X1 U26501 ( .A(1'b0), .B(_02477__PTR323), .S(P3_P1_State2_PTR0), .Z(_03351__PTR259) );
  MUX2_X1 U26502 ( .A(1'b0), .B(_02477__PTR324), .S(P3_P1_State2_PTR0), .Z(_03351__PTR260) );
  MUX2_X1 U26503 ( .A(1'b0), .B(_02477__PTR325), .S(P3_P1_State2_PTR0), .Z(_03351__PTR261) );
  MUX2_X1 U26504 ( .A(1'b0), .B(_02477__PTR326), .S(P3_P1_State2_PTR0), .Z(_03351__PTR262) );
  MUX2_X1 U26505 ( .A(1'b0), .B(_02477__PTR327), .S(P3_P1_State2_PTR0), .Z(_03351__PTR263) );
  MUX2_X1 U26506 ( .A(1'b0), .B(_02477__PTR328), .S(P3_P1_State2_PTR0), .Z(_03351__PTR264) );
  MUX2_X1 U26507 ( .A(1'b0), .B(_02477__PTR329), .S(P3_P1_State2_PTR0), .Z(_03351__PTR265) );
  MUX2_X1 U26508 ( .A(1'b0), .B(_02477__PTR330), .S(P3_P1_State2_PTR0), .Z(_03351__PTR266) );
  MUX2_X1 U26509 ( .A(1'b0), .B(_02477__PTR331), .S(P3_P1_State2_PTR0), .Z(_03351__PTR267) );
  MUX2_X1 U26510 ( .A(1'b0), .B(_02477__PTR332), .S(P3_P1_State2_PTR0), .Z(_03351__PTR268) );
  MUX2_X1 U26511 ( .A(1'b0), .B(_02477__PTR333), .S(P3_P1_State2_PTR0), .Z(_03351__PTR269) );
  MUX2_X1 U26512 ( .A(1'b0), .B(_02477__PTR334), .S(P3_P1_State2_PTR0), .Z(_03351__PTR270) );
  MUX2_X1 U26513 ( .A(1'b0), .B(_02477__PTR335), .S(P3_P1_State2_PTR0), .Z(_03351__PTR271) );
  MUX2_X1 U26514 ( .A(1'b0), .B(_02477__PTR336), .S(P3_P1_State2_PTR0), .Z(_03351__PTR272) );
  MUX2_X1 U26515 ( .A(1'b0), .B(_02477__PTR337), .S(P3_P1_State2_PTR0), .Z(_03351__PTR273) );
  MUX2_X1 U26516 ( .A(1'b0), .B(_02477__PTR338), .S(P3_P1_State2_PTR0), .Z(_03351__PTR274) );
  MUX2_X1 U26517 ( .A(1'b0), .B(_02477__PTR339), .S(P3_P1_State2_PTR0), .Z(_03351__PTR275) );
  MUX2_X1 U26518 ( .A(1'b0), .B(_02477__PTR340), .S(P3_P1_State2_PTR0), .Z(_03351__PTR276) );
  MUX2_X1 U26519 ( .A(1'b0), .B(_02477__PTR341), .S(P3_P1_State2_PTR0), .Z(_03351__PTR277) );
  MUX2_X1 U26520 ( .A(1'b0), .B(_02477__PTR342), .S(P3_P1_State2_PTR0), .Z(_03351__PTR278) );
  MUX2_X1 U26521 ( .A(1'b0), .B(_02477__PTR343), .S(P3_P1_State2_PTR0), .Z(_03351__PTR279) );
  MUX2_X1 U26522 ( .A(1'b0), .B(_02477__PTR344), .S(P3_P1_State2_PTR0), .Z(_03351__PTR280) );
  MUX2_X1 U26523 ( .A(1'b0), .B(_02477__PTR345), .S(P3_P1_State2_PTR0), .Z(_03351__PTR281) );
  MUX2_X1 U26524 ( .A(1'b0), .B(_02477__PTR346), .S(P3_P1_State2_PTR0), .Z(_03351__PTR282) );
  MUX2_X1 U26525 ( .A(1'b0), .B(_02477__PTR347), .S(P3_P1_State2_PTR0), .Z(_03351__PTR283) );
  MUX2_X1 U26526 ( .A(1'b0), .B(_02477__PTR348), .S(P3_P1_State2_PTR0), .Z(_03351__PTR284) );
  MUX2_X1 U26527 ( .A(1'b0), .B(_02477__PTR349), .S(P3_P1_State2_PTR0), .Z(_03351__PTR285) );
  MUX2_X1 U26528 ( .A(1'b0), .B(_02477__PTR350), .S(P3_P1_State2_PTR0), .Z(_03351__PTR286) );
  MUX2_X1 U26529 ( .A(1'b0), .B(_02477__PTR352), .S(P3_P1_State2_PTR0), .Z(_03351__PTR288) );
  MUX2_X1 U26530 ( .A(_03353__PTR0), .B(_03341__PTR0), .S(P3_P1_State2_PTR3), .Z(_02478__PTR0) );
  MUX2_X1 U26531 ( .A(_03353__PTR1), .B(_03341__PTR1), .S(P3_P1_State2_PTR3), .Z(_02478__PTR1) );
  MUX2_X1 U26532 ( .A(_03353__PTR2), .B(_03341__PTR2), .S(P3_P1_State2_PTR3), .Z(_02478__PTR2) );
  MUX2_X1 U26533 ( .A(_03353__PTR3), .B(_03341__PTR3), .S(P3_P1_State2_PTR3), .Z(_02478__PTR3) );
  MUX2_X1 U26534 ( .A(_03353__PTR4), .B(_03341__PTR4), .S(P3_P1_State2_PTR3), .Z(_02478__PTR4) );
  MUX2_X1 U26535 ( .A(_03353__PTR5), .B(_03341__PTR5), .S(P3_P1_State2_PTR3), .Z(_02478__PTR5) );
  MUX2_X1 U26536 ( .A(_03353__PTR6), .B(_03341__PTR6), .S(P3_P1_State2_PTR3), .Z(_02478__PTR6) );
  MUX2_X1 U26537 ( .A(_03353__PTR7), .B(_03341__PTR7), .S(P3_P1_State2_PTR3), .Z(_02478__PTR7) );
  MUX2_X1 U26538 ( .A(_03353__PTR8), .B(_03341__PTR8), .S(P3_P1_State2_PTR3), .Z(_02478__PTR8) );
  MUX2_X1 U26539 ( .A(_03353__PTR9), .B(_03341__PTR9), .S(P3_P1_State2_PTR3), .Z(_02478__PTR9) );
  MUX2_X1 U26540 ( .A(_03353__PTR10), .B(_03341__PTR10), .S(P3_P1_State2_PTR3), .Z(_02478__PTR10) );
  MUX2_X1 U26541 ( .A(_03353__PTR11), .B(_03341__PTR11), .S(P3_P1_State2_PTR3), .Z(_02478__PTR11) );
  MUX2_X1 U26542 ( .A(_03353__PTR12), .B(_03341__PTR12), .S(P3_P1_State2_PTR3), .Z(_02478__PTR12) );
  MUX2_X1 U26543 ( .A(_03353__PTR13), .B(_03341__PTR13), .S(P3_P1_State2_PTR3), .Z(_02478__PTR13) );
  MUX2_X1 U26544 ( .A(_03353__PTR14), .B(_03341__PTR14), .S(P3_P1_State2_PTR3), .Z(_02478__PTR14) );
  MUX2_X1 U26545 ( .A(_03353__PTR15), .B(_03341__PTR15), .S(P3_P1_State2_PTR3), .Z(_02478__PTR15) );
  MUX2_X1 U26546 ( .A(_03353__PTR16), .B(_03341__PTR16), .S(P3_P1_State2_PTR3), .Z(_02478__PTR16) );
  MUX2_X1 U26547 ( .A(_03353__PTR17), .B(_03341__PTR17), .S(P3_P1_State2_PTR3), .Z(_02478__PTR17) );
  MUX2_X1 U26548 ( .A(_03353__PTR18), .B(_03341__PTR18), .S(P3_P1_State2_PTR3), .Z(_02478__PTR18) );
  MUX2_X1 U26549 ( .A(_03353__PTR19), .B(_03341__PTR19), .S(P3_P1_State2_PTR3), .Z(_02478__PTR19) );
  MUX2_X1 U26550 ( .A(_03353__PTR20), .B(_03341__PTR20), .S(P3_P1_State2_PTR3), .Z(_02478__PTR20) );
  MUX2_X1 U26551 ( .A(_03353__PTR21), .B(_03341__PTR21), .S(P3_P1_State2_PTR3), .Z(_02478__PTR21) );
  MUX2_X1 U26552 ( .A(_03353__PTR22), .B(_03341__PTR22), .S(P3_P1_State2_PTR3), .Z(_02478__PTR22) );
  MUX2_X1 U26553 ( .A(_03353__PTR23), .B(_03341__PTR23), .S(P3_P1_State2_PTR3), .Z(_02478__PTR23) );
  MUX2_X1 U26554 ( .A(_03353__PTR24), .B(_03341__PTR24), .S(P3_P1_State2_PTR3), .Z(_02478__PTR24) );
  MUX2_X1 U26555 ( .A(_03353__PTR25), .B(_03341__PTR25), .S(P3_P1_State2_PTR3), .Z(_02478__PTR25) );
  MUX2_X1 U26556 ( .A(_03353__PTR26), .B(_03341__PTR26), .S(P3_P1_State2_PTR3), .Z(_02478__PTR26) );
  MUX2_X1 U26557 ( .A(_03353__PTR27), .B(_03341__PTR27), .S(P3_P1_State2_PTR3), .Z(_02478__PTR27) );
  MUX2_X1 U26558 ( .A(_03353__PTR28), .B(_03341__PTR28), .S(P3_P1_State2_PTR3), .Z(_02478__PTR28) );
  MUX2_X1 U26559 ( .A(_03353__PTR29), .B(_03341__PTR29), .S(P3_P1_State2_PTR3), .Z(_02478__PTR29) );
  MUX2_X1 U26560 ( .A(_03353__PTR30), .B(_03341__PTR30), .S(P3_P1_State2_PTR3), .Z(_02478__PTR30) );
  MUX2_X1 U26561 ( .A(_03353__PTR32), .B(_03341__PTR31), .S(P3_P1_State2_PTR3), .Z(_02478__PTR32) );
  MUX2_X1 U26562 ( .A(_03352__PTR0), .B(_03352__PTR256), .S(P3_P1_State2_PTR2), .Z(_03353__PTR0) );
  MUX2_X1 U26563 ( .A(_03352__PTR1), .B(_03352__PTR257), .S(P3_P1_State2_PTR2), .Z(_03353__PTR1) );
  MUX2_X1 U26564 ( .A(_03352__PTR2), .B(_03352__PTR258), .S(P3_P1_State2_PTR2), .Z(_03353__PTR2) );
  MUX2_X1 U26565 ( .A(_03352__PTR3), .B(_03352__PTR259), .S(P3_P1_State2_PTR2), .Z(_03353__PTR3) );
  MUX2_X1 U26566 ( .A(_03352__PTR4), .B(_03352__PTR260), .S(P3_P1_State2_PTR2), .Z(_03353__PTR4) );
  MUX2_X1 U26567 ( .A(_03352__PTR5), .B(_03352__PTR261), .S(P3_P1_State2_PTR2), .Z(_03353__PTR5) );
  MUX2_X1 U26568 ( .A(_03352__PTR6), .B(_03352__PTR262), .S(P3_P1_State2_PTR2), .Z(_03353__PTR6) );
  MUX2_X1 U26569 ( .A(_03352__PTR7), .B(_03352__PTR263), .S(P3_P1_State2_PTR2), .Z(_03353__PTR7) );
  MUX2_X1 U26570 ( .A(_03352__PTR8), .B(_03352__PTR264), .S(P3_P1_State2_PTR2), .Z(_03353__PTR8) );
  MUX2_X1 U26571 ( .A(_03352__PTR9), .B(_03352__PTR265), .S(P3_P1_State2_PTR2), .Z(_03353__PTR9) );
  MUX2_X1 U26572 ( .A(_03352__PTR10), .B(_03352__PTR266), .S(P3_P1_State2_PTR2), .Z(_03353__PTR10) );
  MUX2_X1 U26573 ( .A(_03352__PTR11), .B(_03352__PTR267), .S(P3_P1_State2_PTR2), .Z(_03353__PTR11) );
  MUX2_X1 U26574 ( .A(_03352__PTR12), .B(_03352__PTR268), .S(P3_P1_State2_PTR2), .Z(_03353__PTR12) );
  MUX2_X1 U26575 ( .A(_03352__PTR13), .B(_03352__PTR269), .S(P3_P1_State2_PTR2), .Z(_03353__PTR13) );
  MUX2_X1 U26576 ( .A(_03352__PTR14), .B(_03352__PTR270), .S(P3_P1_State2_PTR2), .Z(_03353__PTR14) );
  MUX2_X1 U26577 ( .A(_03352__PTR15), .B(_03352__PTR271), .S(P3_P1_State2_PTR2), .Z(_03353__PTR15) );
  MUX2_X1 U26578 ( .A(_03352__PTR16), .B(_03352__PTR272), .S(P3_P1_State2_PTR2), .Z(_03353__PTR16) );
  MUX2_X1 U26579 ( .A(_03352__PTR17), .B(_03352__PTR273), .S(P3_P1_State2_PTR2), .Z(_03353__PTR17) );
  MUX2_X1 U26580 ( .A(_03352__PTR18), .B(_03352__PTR274), .S(P3_P1_State2_PTR2), .Z(_03353__PTR18) );
  MUX2_X1 U26581 ( .A(_03352__PTR19), .B(_03352__PTR275), .S(P3_P1_State2_PTR2), .Z(_03353__PTR19) );
  MUX2_X1 U26582 ( .A(_03352__PTR20), .B(_03352__PTR276), .S(P3_P1_State2_PTR2), .Z(_03353__PTR20) );
  MUX2_X1 U26583 ( .A(_03352__PTR21), .B(_03352__PTR277), .S(P3_P1_State2_PTR2), .Z(_03353__PTR21) );
  MUX2_X1 U26584 ( .A(_03352__PTR22), .B(_03352__PTR278), .S(P3_P1_State2_PTR2), .Z(_03353__PTR22) );
  MUX2_X1 U26585 ( .A(_03352__PTR23), .B(_03352__PTR279), .S(P3_P1_State2_PTR2), .Z(_03353__PTR23) );
  MUX2_X1 U26586 ( .A(_03352__PTR24), .B(_03352__PTR280), .S(P3_P1_State2_PTR2), .Z(_03353__PTR24) );
  MUX2_X1 U26587 ( .A(_03352__PTR25), .B(_03352__PTR281), .S(P3_P1_State2_PTR2), .Z(_03353__PTR25) );
  MUX2_X1 U26588 ( .A(_03352__PTR26), .B(_03352__PTR282), .S(P3_P1_State2_PTR2), .Z(_03353__PTR26) );
  MUX2_X1 U26589 ( .A(_03352__PTR27), .B(_03352__PTR283), .S(P3_P1_State2_PTR2), .Z(_03353__PTR27) );
  MUX2_X1 U26590 ( .A(_03352__PTR28), .B(_03352__PTR284), .S(P3_P1_State2_PTR2), .Z(_03353__PTR28) );
  MUX2_X1 U26591 ( .A(_03352__PTR29), .B(_03352__PTR285), .S(P3_P1_State2_PTR2), .Z(_03353__PTR29) );
  MUX2_X1 U26592 ( .A(_03352__PTR30), .B(_03352__PTR286), .S(P3_P1_State2_PTR2), .Z(_03353__PTR30) );
  MUX2_X1 U26593 ( .A(_03352__PTR32), .B(_03352__PTR288), .S(P3_P1_State2_PTR2), .Z(_03353__PTR32) );
  MUX2_X1 U26594 ( .A(_03356__PTR0), .B(_03354__PTR64), .S(P3_P1_State2_PTR3), .Z(_02480__PTR0) );
  MUX2_X1 U26595 ( .A(_03356__PTR1), .B(_03354__PTR65), .S(P3_P1_State2_PTR3), .Z(_02480__PTR1) );
  MUX2_X1 U26596 ( .A(_03356__PTR2), .B(_03354__PTR66), .S(P3_P1_State2_PTR3), .Z(_02480__PTR2) );
  MUX2_X1 U26597 ( .A(_03356__PTR3), .B(_03354__PTR67), .S(P3_P1_State2_PTR3), .Z(_02480__PTR3) );
  MUX2_X1 U26598 ( .A(_03356__PTR4), .B(_03354__PTR68), .S(P3_P1_State2_PTR3), .Z(_02480__PTR4) );
  MUX2_X1 U26599 ( .A(_03356__PTR5), .B(_03354__PTR69), .S(P3_P1_State2_PTR3), .Z(_02480__PTR5) );
  MUX2_X1 U26600 ( .A(_03356__PTR6), .B(_03354__PTR70), .S(P3_P1_State2_PTR3), .Z(_02480__PTR6) );
  MUX2_X1 U26601 ( .A(_03356__PTR7), .B(_03354__PTR71), .S(P3_P1_State2_PTR3), .Z(_02480__PTR7) );
  MUX2_X1 U26602 ( .A(_03355__PTR0), .B(_03355__PTR32), .S(P3_P1_State2_PTR2), .Z(_03356__PTR0) );
  MUX2_X1 U26603 ( .A(_03355__PTR1), .B(_03355__PTR33), .S(P3_P1_State2_PTR2), .Z(_03356__PTR1) );
  MUX2_X1 U26604 ( .A(_03355__PTR2), .B(_03355__PTR34), .S(P3_P1_State2_PTR2), .Z(_03356__PTR2) );
  MUX2_X1 U26605 ( .A(_03355__PTR3), .B(_03355__PTR35), .S(P3_P1_State2_PTR2), .Z(_03356__PTR3) );
  MUX2_X1 U26606 ( .A(_03355__PTR4), .B(_03355__PTR36), .S(P3_P1_State2_PTR2), .Z(_03356__PTR4) );
  MUX2_X1 U26607 ( .A(_03355__PTR5), .B(_03355__PTR37), .S(P3_P1_State2_PTR2), .Z(_03356__PTR5) );
  MUX2_X1 U26608 ( .A(_03355__PTR6), .B(_03355__PTR38), .S(P3_P1_State2_PTR2), .Z(_03356__PTR6) );
  MUX2_X1 U26609 ( .A(_03355__PTR7), .B(_03355__PTR39), .S(P3_P1_State2_PTR2), .Z(_03356__PTR7) );
  MUX2_X1 U26610 ( .A(1'b0), .B(_03354__PTR16), .S(P3_P1_State2_PTR1), .Z(_03355__PTR0) );
  MUX2_X1 U26611 ( .A(1'b0), .B(_03354__PTR17), .S(P3_P1_State2_PTR1), .Z(_03355__PTR1) );
  MUX2_X1 U26612 ( .A(1'b0), .B(_03354__PTR18), .S(P3_P1_State2_PTR1), .Z(_03355__PTR2) );
  MUX2_X1 U26613 ( .A(1'b0), .B(_03354__PTR19), .S(P3_P1_State2_PTR1), .Z(_03355__PTR3) );
  MUX2_X1 U26614 ( .A(1'b0), .B(_03354__PTR20), .S(P3_P1_State2_PTR1), .Z(_03355__PTR4) );
  MUX2_X1 U26615 ( .A(1'b0), .B(_03354__PTR21), .S(P3_P1_State2_PTR1), .Z(_03355__PTR5) );
  MUX2_X1 U26616 ( .A(1'b0), .B(_03354__PTR22), .S(P3_P1_State2_PTR1), .Z(_03355__PTR6) );
  MUX2_X1 U26617 ( .A(1'b0), .B(_03354__PTR23), .S(P3_P1_State2_PTR1), .Z(_03355__PTR7) );
  MUX2_X1 U26618 ( .A(_03354__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03355__PTR32) );
  MUX2_X1 U26619 ( .A(_03354__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03355__PTR33) );
  MUX2_X1 U26620 ( .A(_03354__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03355__PTR34) );
  MUX2_X1 U26621 ( .A(_03354__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03355__PTR35) );
  MUX2_X1 U26622 ( .A(_03354__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03355__PTR36) );
  MUX2_X1 U26623 ( .A(_03354__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03355__PTR37) );
  MUX2_X1 U26624 ( .A(_03354__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03355__PTR38) );
  MUX2_X1 U26625 ( .A(_03354__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03355__PTR39) );
  MUX2_X1 U26626 ( .A(_02479__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR16) );
  MUX2_X1 U26627 ( .A(_02479__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR17) );
  MUX2_X1 U26628 ( .A(_02479__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR18) );
  MUX2_X1 U26629 ( .A(_02479__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR19) );
  MUX2_X1 U26630 ( .A(_02479__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR20) );
  MUX2_X1 U26631 ( .A(_02479__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR21) );
  MUX2_X1 U26632 ( .A(_02479__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR22) );
  MUX2_X1 U26633 ( .A(_02479__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR23) );
  MUX2_X1 U26634 ( .A(_02479__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR32) );
  MUX2_X1 U26635 ( .A(_02479__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR33) );
  MUX2_X1 U26636 ( .A(_02479__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR34) );
  MUX2_X1 U26637 ( .A(_02479__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR35) );
  MUX2_X1 U26638 ( .A(_02479__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR36) );
  MUX2_X1 U26639 ( .A(_02479__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR37) );
  MUX2_X1 U26640 ( .A(_02479__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR38) );
  MUX2_X1 U26641 ( .A(_02479__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR39) );
  MUX2_X1 U26642 ( .A(_02479__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR64) );
  MUX2_X1 U26643 ( .A(_02479__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR65) );
  MUX2_X1 U26644 ( .A(_02479__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR66) );
  MUX2_X1 U26645 ( .A(_02479__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR67) );
  MUX2_X1 U26646 ( .A(_02479__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR68) );
  MUX2_X1 U26647 ( .A(_02479__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR69) );
  MUX2_X1 U26648 ( .A(_02479__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR70) );
  MUX2_X1 U26649 ( .A(_02479__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03354__PTR71) );
  MUX2_X1 U26650 ( .A(_03359__PTR0), .B(_03357__PTR64), .S(P3_P1_State2_PTR3), .Z(_02482__PTR0) );
  MUX2_X1 U26651 ( .A(_03359__PTR1), .B(_03357__PTR65), .S(P3_P1_State2_PTR3), .Z(_02482__PTR1) );
  MUX2_X1 U26652 ( .A(_03359__PTR2), .B(_03357__PTR66), .S(P3_P1_State2_PTR3), .Z(_02482__PTR2) );
  MUX2_X1 U26653 ( .A(_03359__PTR3), .B(_03357__PTR67), .S(P3_P1_State2_PTR3), .Z(_02482__PTR3) );
  MUX2_X1 U26654 ( .A(_03359__PTR4), .B(_03357__PTR68), .S(P3_P1_State2_PTR3), .Z(_02482__PTR4) );
  MUX2_X1 U26655 ( .A(_03359__PTR5), .B(_03357__PTR69), .S(P3_P1_State2_PTR3), .Z(_02482__PTR5) );
  MUX2_X1 U26656 ( .A(_03359__PTR6), .B(_03357__PTR70), .S(P3_P1_State2_PTR3), .Z(_02482__PTR6) );
  MUX2_X1 U26657 ( .A(_03359__PTR7), .B(_03357__PTR71), .S(P3_P1_State2_PTR3), .Z(_02482__PTR7) );
  MUX2_X1 U26658 ( .A(_03358__PTR0), .B(_03358__PTR32), .S(P3_P1_State2_PTR2), .Z(_03359__PTR0) );
  MUX2_X1 U26659 ( .A(_03358__PTR1), .B(_03358__PTR33), .S(P3_P1_State2_PTR2), .Z(_03359__PTR1) );
  MUX2_X1 U26660 ( .A(_03358__PTR2), .B(_03358__PTR34), .S(P3_P1_State2_PTR2), .Z(_03359__PTR2) );
  MUX2_X1 U26661 ( .A(_03358__PTR3), .B(_03358__PTR35), .S(P3_P1_State2_PTR2), .Z(_03359__PTR3) );
  MUX2_X1 U26662 ( .A(_03358__PTR4), .B(_03358__PTR36), .S(P3_P1_State2_PTR2), .Z(_03359__PTR4) );
  MUX2_X1 U26663 ( .A(_03358__PTR5), .B(_03358__PTR37), .S(P3_P1_State2_PTR2), .Z(_03359__PTR5) );
  MUX2_X1 U26664 ( .A(_03358__PTR6), .B(_03358__PTR38), .S(P3_P1_State2_PTR2), .Z(_03359__PTR6) );
  MUX2_X1 U26665 ( .A(_03358__PTR7), .B(_03358__PTR39), .S(P3_P1_State2_PTR2), .Z(_03359__PTR7) );
  MUX2_X1 U26666 ( .A(1'b0), .B(_03357__PTR16), .S(P3_P1_State2_PTR1), .Z(_03358__PTR0) );
  MUX2_X1 U26667 ( .A(1'b0), .B(_03357__PTR17), .S(P3_P1_State2_PTR1), .Z(_03358__PTR1) );
  MUX2_X1 U26668 ( .A(1'b0), .B(_03357__PTR18), .S(P3_P1_State2_PTR1), .Z(_03358__PTR2) );
  MUX2_X1 U26669 ( .A(1'b0), .B(_03357__PTR19), .S(P3_P1_State2_PTR1), .Z(_03358__PTR3) );
  MUX2_X1 U26670 ( .A(1'b0), .B(_03357__PTR20), .S(P3_P1_State2_PTR1), .Z(_03358__PTR4) );
  MUX2_X1 U26671 ( .A(1'b0), .B(_03357__PTR21), .S(P3_P1_State2_PTR1), .Z(_03358__PTR5) );
  MUX2_X1 U26672 ( .A(1'b0), .B(_03357__PTR22), .S(P3_P1_State2_PTR1), .Z(_03358__PTR6) );
  MUX2_X1 U26673 ( .A(1'b0), .B(_03357__PTR23), .S(P3_P1_State2_PTR1), .Z(_03358__PTR7) );
  MUX2_X1 U26674 ( .A(_03357__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03358__PTR32) );
  MUX2_X1 U26675 ( .A(_03357__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03358__PTR33) );
  MUX2_X1 U26676 ( .A(_03357__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03358__PTR34) );
  MUX2_X1 U26677 ( .A(_03357__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03358__PTR35) );
  MUX2_X1 U26678 ( .A(_03357__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03358__PTR36) );
  MUX2_X1 U26679 ( .A(_03357__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03358__PTR37) );
  MUX2_X1 U26680 ( .A(_03357__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03358__PTR38) );
  MUX2_X1 U26681 ( .A(_03357__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03358__PTR39) );
  MUX2_X1 U26682 ( .A(_02481__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR16) );
  MUX2_X1 U26683 ( .A(_02481__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR17) );
  MUX2_X1 U26684 ( .A(_02481__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR18) );
  MUX2_X1 U26685 ( .A(_02481__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR19) );
  MUX2_X1 U26686 ( .A(_02481__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR20) );
  MUX2_X1 U26687 ( .A(_02481__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR21) );
  MUX2_X1 U26688 ( .A(_02481__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR22) );
  MUX2_X1 U26689 ( .A(_02481__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR23) );
  MUX2_X1 U26690 ( .A(_02481__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR32) );
  MUX2_X1 U26691 ( .A(_02481__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR33) );
  MUX2_X1 U26692 ( .A(_02481__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR34) );
  MUX2_X1 U26693 ( .A(_02481__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR35) );
  MUX2_X1 U26694 ( .A(_02481__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR36) );
  MUX2_X1 U26695 ( .A(_02481__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR37) );
  MUX2_X1 U26696 ( .A(_02481__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR38) );
  MUX2_X1 U26697 ( .A(_02481__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR39) );
  MUX2_X1 U26698 ( .A(_02481__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR64) );
  MUX2_X1 U26699 ( .A(_02481__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR65) );
  MUX2_X1 U26700 ( .A(_02481__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR66) );
  MUX2_X1 U26701 ( .A(_02481__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR67) );
  MUX2_X1 U26702 ( .A(_02481__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR68) );
  MUX2_X1 U26703 ( .A(_02481__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR69) );
  MUX2_X1 U26704 ( .A(_02481__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR70) );
  MUX2_X1 U26705 ( .A(_02481__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03357__PTR71) );
  MUX2_X1 U26706 ( .A(_03362__PTR0), .B(_03360__PTR64), .S(P3_P1_State2_PTR3), .Z(_02484__PTR0) );
  MUX2_X1 U26707 ( .A(_03362__PTR1), .B(_03360__PTR65), .S(P3_P1_State2_PTR3), .Z(_02484__PTR1) );
  MUX2_X1 U26708 ( .A(_03362__PTR2), .B(_03360__PTR66), .S(P3_P1_State2_PTR3), .Z(_02484__PTR2) );
  MUX2_X1 U26709 ( .A(_03362__PTR3), .B(_03360__PTR67), .S(P3_P1_State2_PTR3), .Z(_02484__PTR3) );
  MUX2_X1 U26710 ( .A(_03362__PTR4), .B(_03360__PTR68), .S(P3_P1_State2_PTR3), .Z(_02484__PTR4) );
  MUX2_X1 U26711 ( .A(_03362__PTR5), .B(_03360__PTR69), .S(P3_P1_State2_PTR3), .Z(_02484__PTR5) );
  MUX2_X1 U26712 ( .A(_03362__PTR6), .B(_03360__PTR70), .S(P3_P1_State2_PTR3), .Z(_02484__PTR6) );
  MUX2_X1 U26713 ( .A(_03362__PTR7), .B(_03360__PTR71), .S(P3_P1_State2_PTR3), .Z(_02484__PTR7) );
  MUX2_X1 U26714 ( .A(_03361__PTR0), .B(_03361__PTR32), .S(P3_P1_State2_PTR2), .Z(_03362__PTR0) );
  MUX2_X1 U26715 ( .A(_03361__PTR1), .B(_03361__PTR33), .S(P3_P1_State2_PTR2), .Z(_03362__PTR1) );
  MUX2_X1 U26716 ( .A(_03361__PTR2), .B(_03361__PTR34), .S(P3_P1_State2_PTR2), .Z(_03362__PTR2) );
  MUX2_X1 U26717 ( .A(_03361__PTR3), .B(_03361__PTR35), .S(P3_P1_State2_PTR2), .Z(_03362__PTR3) );
  MUX2_X1 U26718 ( .A(_03361__PTR4), .B(_03361__PTR36), .S(P3_P1_State2_PTR2), .Z(_03362__PTR4) );
  MUX2_X1 U26719 ( .A(_03361__PTR5), .B(_03361__PTR37), .S(P3_P1_State2_PTR2), .Z(_03362__PTR5) );
  MUX2_X1 U26720 ( .A(_03361__PTR6), .B(_03361__PTR38), .S(P3_P1_State2_PTR2), .Z(_03362__PTR6) );
  MUX2_X1 U26721 ( .A(_03361__PTR7), .B(_03361__PTR39), .S(P3_P1_State2_PTR2), .Z(_03362__PTR7) );
  MUX2_X1 U26722 ( .A(1'b0), .B(_03360__PTR16), .S(P3_P1_State2_PTR1), .Z(_03361__PTR0) );
  MUX2_X1 U26723 ( .A(1'b0), .B(_03360__PTR17), .S(P3_P1_State2_PTR1), .Z(_03361__PTR1) );
  MUX2_X1 U26724 ( .A(1'b0), .B(_03360__PTR18), .S(P3_P1_State2_PTR1), .Z(_03361__PTR2) );
  MUX2_X1 U26725 ( .A(1'b0), .B(_03360__PTR19), .S(P3_P1_State2_PTR1), .Z(_03361__PTR3) );
  MUX2_X1 U26726 ( .A(1'b0), .B(_03360__PTR20), .S(P3_P1_State2_PTR1), .Z(_03361__PTR4) );
  MUX2_X1 U26727 ( .A(1'b0), .B(_03360__PTR21), .S(P3_P1_State2_PTR1), .Z(_03361__PTR5) );
  MUX2_X1 U26728 ( .A(1'b0), .B(_03360__PTR22), .S(P3_P1_State2_PTR1), .Z(_03361__PTR6) );
  MUX2_X1 U26729 ( .A(1'b0), .B(_03360__PTR23), .S(P3_P1_State2_PTR1), .Z(_03361__PTR7) );
  MUX2_X1 U26730 ( .A(_03360__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03361__PTR32) );
  MUX2_X1 U26731 ( .A(_03360__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03361__PTR33) );
  MUX2_X1 U26732 ( .A(_03360__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03361__PTR34) );
  MUX2_X1 U26733 ( .A(_03360__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03361__PTR35) );
  MUX2_X1 U26734 ( .A(_03360__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03361__PTR36) );
  MUX2_X1 U26735 ( .A(_03360__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03361__PTR37) );
  MUX2_X1 U26736 ( .A(_03360__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03361__PTR38) );
  MUX2_X1 U26737 ( .A(_03360__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03361__PTR39) );
  MUX2_X1 U26738 ( .A(_02483__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR16) );
  MUX2_X1 U26739 ( .A(_02483__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR17) );
  MUX2_X1 U26740 ( .A(_02483__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR18) );
  MUX2_X1 U26741 ( .A(_02483__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR19) );
  MUX2_X1 U26742 ( .A(_02483__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR20) );
  MUX2_X1 U26743 ( .A(_02483__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR21) );
  MUX2_X1 U26744 ( .A(_02483__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR22) );
  MUX2_X1 U26745 ( .A(_02483__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR23) );
  MUX2_X1 U26746 ( .A(_02483__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR32) );
  MUX2_X1 U26747 ( .A(_02483__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR33) );
  MUX2_X1 U26748 ( .A(_02483__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR34) );
  MUX2_X1 U26749 ( .A(_02483__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR35) );
  MUX2_X1 U26750 ( .A(_02483__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR36) );
  MUX2_X1 U26751 ( .A(_02483__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR37) );
  MUX2_X1 U26752 ( .A(_02483__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR38) );
  MUX2_X1 U26753 ( .A(_02483__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR39) );
  MUX2_X1 U26754 ( .A(_02483__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR64) );
  MUX2_X1 U26755 ( .A(_02483__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR65) );
  MUX2_X1 U26756 ( .A(_02483__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR66) );
  MUX2_X1 U26757 ( .A(_02483__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR67) );
  MUX2_X1 U26758 ( .A(_02483__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR68) );
  MUX2_X1 U26759 ( .A(_02483__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR69) );
  MUX2_X1 U26760 ( .A(_02483__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR70) );
  MUX2_X1 U26761 ( .A(_02483__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03360__PTR71) );
  MUX2_X1 U26762 ( .A(_03365__PTR0), .B(_03363__PTR64), .S(P3_P1_State2_PTR3), .Z(_02486__PTR0) );
  MUX2_X1 U26763 ( .A(_03365__PTR1), .B(_03363__PTR65), .S(P3_P1_State2_PTR3), .Z(_02486__PTR1) );
  MUX2_X1 U26764 ( .A(_03365__PTR2), .B(_03363__PTR66), .S(P3_P1_State2_PTR3), .Z(_02486__PTR2) );
  MUX2_X1 U26765 ( .A(_03365__PTR3), .B(_03363__PTR67), .S(P3_P1_State2_PTR3), .Z(_02486__PTR3) );
  MUX2_X1 U26766 ( .A(_03365__PTR4), .B(_03363__PTR68), .S(P3_P1_State2_PTR3), .Z(_02486__PTR4) );
  MUX2_X1 U26767 ( .A(_03365__PTR5), .B(_03363__PTR69), .S(P3_P1_State2_PTR3), .Z(_02486__PTR5) );
  MUX2_X1 U26768 ( .A(_03365__PTR6), .B(_03363__PTR70), .S(P3_P1_State2_PTR3), .Z(_02486__PTR6) );
  MUX2_X1 U26769 ( .A(_03365__PTR7), .B(_03363__PTR71), .S(P3_P1_State2_PTR3), .Z(_02486__PTR7) );
  MUX2_X1 U26770 ( .A(_03364__PTR0), .B(_03364__PTR32), .S(P3_P1_State2_PTR2), .Z(_03365__PTR0) );
  MUX2_X1 U26771 ( .A(_03364__PTR1), .B(_03364__PTR33), .S(P3_P1_State2_PTR2), .Z(_03365__PTR1) );
  MUX2_X1 U26772 ( .A(_03364__PTR2), .B(_03364__PTR34), .S(P3_P1_State2_PTR2), .Z(_03365__PTR2) );
  MUX2_X1 U26773 ( .A(_03364__PTR3), .B(_03364__PTR35), .S(P3_P1_State2_PTR2), .Z(_03365__PTR3) );
  MUX2_X1 U26774 ( .A(_03364__PTR4), .B(_03364__PTR36), .S(P3_P1_State2_PTR2), .Z(_03365__PTR4) );
  MUX2_X1 U26775 ( .A(_03364__PTR5), .B(_03364__PTR37), .S(P3_P1_State2_PTR2), .Z(_03365__PTR5) );
  MUX2_X1 U26776 ( .A(_03364__PTR6), .B(_03364__PTR38), .S(P3_P1_State2_PTR2), .Z(_03365__PTR6) );
  MUX2_X1 U26777 ( .A(_03364__PTR7), .B(_03364__PTR39), .S(P3_P1_State2_PTR2), .Z(_03365__PTR7) );
  MUX2_X1 U26778 ( .A(1'b0), .B(_03363__PTR16), .S(P3_P1_State2_PTR1), .Z(_03364__PTR0) );
  MUX2_X1 U26779 ( .A(1'b0), .B(_03363__PTR17), .S(P3_P1_State2_PTR1), .Z(_03364__PTR1) );
  MUX2_X1 U26780 ( .A(1'b0), .B(_03363__PTR18), .S(P3_P1_State2_PTR1), .Z(_03364__PTR2) );
  MUX2_X1 U26781 ( .A(1'b0), .B(_03363__PTR19), .S(P3_P1_State2_PTR1), .Z(_03364__PTR3) );
  MUX2_X1 U26782 ( .A(1'b0), .B(_03363__PTR20), .S(P3_P1_State2_PTR1), .Z(_03364__PTR4) );
  MUX2_X1 U26783 ( .A(1'b0), .B(_03363__PTR21), .S(P3_P1_State2_PTR1), .Z(_03364__PTR5) );
  MUX2_X1 U26784 ( .A(1'b0), .B(_03363__PTR22), .S(P3_P1_State2_PTR1), .Z(_03364__PTR6) );
  MUX2_X1 U26785 ( .A(1'b0), .B(_03363__PTR23), .S(P3_P1_State2_PTR1), .Z(_03364__PTR7) );
  MUX2_X1 U26786 ( .A(_03363__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03364__PTR32) );
  MUX2_X1 U26787 ( .A(_03363__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03364__PTR33) );
  MUX2_X1 U26788 ( .A(_03363__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03364__PTR34) );
  MUX2_X1 U26789 ( .A(_03363__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03364__PTR35) );
  MUX2_X1 U26790 ( .A(_03363__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03364__PTR36) );
  MUX2_X1 U26791 ( .A(_03363__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03364__PTR37) );
  MUX2_X1 U26792 ( .A(_03363__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03364__PTR38) );
  MUX2_X1 U26793 ( .A(_03363__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03364__PTR39) );
  MUX2_X1 U26794 ( .A(_02485__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR16) );
  MUX2_X1 U26795 ( .A(_02485__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR17) );
  MUX2_X1 U26796 ( .A(_02485__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR18) );
  MUX2_X1 U26797 ( .A(_02485__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR19) );
  MUX2_X1 U26798 ( .A(_02485__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR20) );
  MUX2_X1 U26799 ( .A(_02485__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR21) );
  MUX2_X1 U26800 ( .A(_02485__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR22) );
  MUX2_X1 U26801 ( .A(_02485__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR23) );
  MUX2_X1 U26802 ( .A(_02485__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR32) );
  MUX2_X1 U26803 ( .A(_02485__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR33) );
  MUX2_X1 U26804 ( .A(_02485__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR34) );
  MUX2_X1 U26805 ( .A(_02485__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR35) );
  MUX2_X1 U26806 ( .A(_02485__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR36) );
  MUX2_X1 U26807 ( .A(_02485__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR37) );
  MUX2_X1 U26808 ( .A(_02485__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR38) );
  MUX2_X1 U26809 ( .A(_02485__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR39) );
  MUX2_X1 U26810 ( .A(_02485__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR64) );
  MUX2_X1 U26811 ( .A(_02485__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR65) );
  MUX2_X1 U26812 ( .A(_02485__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR66) );
  MUX2_X1 U26813 ( .A(_02485__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR67) );
  MUX2_X1 U26814 ( .A(_02485__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR68) );
  MUX2_X1 U26815 ( .A(_02485__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR69) );
  MUX2_X1 U26816 ( .A(_02485__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR70) );
  MUX2_X1 U26817 ( .A(_02485__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03363__PTR71) );
  MUX2_X1 U26818 ( .A(_03368__PTR0), .B(_03366__PTR64), .S(P3_P1_State2_PTR3), .Z(_02488__PTR0) );
  MUX2_X1 U26819 ( .A(_03368__PTR1), .B(_03366__PTR65), .S(P3_P1_State2_PTR3), .Z(_02488__PTR1) );
  MUX2_X1 U26820 ( .A(_03368__PTR2), .B(_03366__PTR66), .S(P3_P1_State2_PTR3), .Z(_02488__PTR2) );
  MUX2_X1 U26821 ( .A(_03368__PTR3), .B(_03366__PTR67), .S(P3_P1_State2_PTR3), .Z(_02488__PTR3) );
  MUX2_X1 U26822 ( .A(_03368__PTR4), .B(_03366__PTR68), .S(P3_P1_State2_PTR3), .Z(_02488__PTR4) );
  MUX2_X1 U26823 ( .A(_03368__PTR5), .B(_03366__PTR69), .S(P3_P1_State2_PTR3), .Z(_02488__PTR5) );
  MUX2_X1 U26824 ( .A(_03368__PTR6), .B(_03366__PTR70), .S(P3_P1_State2_PTR3), .Z(_02488__PTR6) );
  MUX2_X1 U26825 ( .A(_03368__PTR7), .B(_03366__PTR71), .S(P3_P1_State2_PTR3), .Z(_02488__PTR7) );
  MUX2_X1 U26826 ( .A(_03367__PTR0), .B(_03367__PTR32), .S(P3_P1_State2_PTR2), .Z(_03368__PTR0) );
  MUX2_X1 U26827 ( .A(_03367__PTR1), .B(_03367__PTR33), .S(P3_P1_State2_PTR2), .Z(_03368__PTR1) );
  MUX2_X1 U26828 ( .A(_03367__PTR2), .B(_03367__PTR34), .S(P3_P1_State2_PTR2), .Z(_03368__PTR2) );
  MUX2_X1 U26829 ( .A(_03367__PTR3), .B(_03367__PTR35), .S(P3_P1_State2_PTR2), .Z(_03368__PTR3) );
  MUX2_X1 U26830 ( .A(_03367__PTR4), .B(_03367__PTR36), .S(P3_P1_State2_PTR2), .Z(_03368__PTR4) );
  MUX2_X1 U26831 ( .A(_03367__PTR5), .B(_03367__PTR37), .S(P3_P1_State2_PTR2), .Z(_03368__PTR5) );
  MUX2_X1 U26832 ( .A(_03367__PTR6), .B(_03367__PTR38), .S(P3_P1_State2_PTR2), .Z(_03368__PTR6) );
  MUX2_X1 U26833 ( .A(_03367__PTR7), .B(_03367__PTR39), .S(P3_P1_State2_PTR2), .Z(_03368__PTR7) );
  MUX2_X1 U26834 ( .A(1'b0), .B(_03366__PTR16), .S(P3_P1_State2_PTR1), .Z(_03367__PTR0) );
  MUX2_X1 U26835 ( .A(1'b0), .B(_03366__PTR17), .S(P3_P1_State2_PTR1), .Z(_03367__PTR1) );
  MUX2_X1 U26836 ( .A(1'b0), .B(_03366__PTR18), .S(P3_P1_State2_PTR1), .Z(_03367__PTR2) );
  MUX2_X1 U26837 ( .A(1'b0), .B(_03366__PTR19), .S(P3_P1_State2_PTR1), .Z(_03367__PTR3) );
  MUX2_X1 U26838 ( .A(1'b0), .B(_03366__PTR20), .S(P3_P1_State2_PTR1), .Z(_03367__PTR4) );
  MUX2_X1 U26839 ( .A(1'b0), .B(_03366__PTR21), .S(P3_P1_State2_PTR1), .Z(_03367__PTR5) );
  MUX2_X1 U26840 ( .A(1'b0), .B(_03366__PTR22), .S(P3_P1_State2_PTR1), .Z(_03367__PTR6) );
  MUX2_X1 U26841 ( .A(1'b0), .B(_03366__PTR23), .S(P3_P1_State2_PTR1), .Z(_03367__PTR7) );
  MUX2_X1 U26842 ( .A(_03366__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03367__PTR32) );
  MUX2_X1 U26843 ( .A(_03366__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03367__PTR33) );
  MUX2_X1 U26844 ( .A(_03366__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03367__PTR34) );
  MUX2_X1 U26845 ( .A(_03366__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03367__PTR35) );
  MUX2_X1 U26846 ( .A(_03366__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03367__PTR36) );
  MUX2_X1 U26847 ( .A(_03366__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03367__PTR37) );
  MUX2_X1 U26848 ( .A(_03366__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03367__PTR38) );
  MUX2_X1 U26849 ( .A(_03366__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03367__PTR39) );
  MUX2_X1 U26850 ( .A(_02487__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR16) );
  MUX2_X1 U26851 ( .A(_02487__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR17) );
  MUX2_X1 U26852 ( .A(_02487__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR18) );
  MUX2_X1 U26853 ( .A(_02487__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR19) );
  MUX2_X1 U26854 ( .A(_02487__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR20) );
  MUX2_X1 U26855 ( .A(_02487__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR21) );
  MUX2_X1 U26856 ( .A(_02487__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR22) );
  MUX2_X1 U26857 ( .A(_02487__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR23) );
  MUX2_X1 U26858 ( .A(_02487__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR32) );
  MUX2_X1 U26859 ( .A(_02487__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR33) );
  MUX2_X1 U26860 ( .A(_02487__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR34) );
  MUX2_X1 U26861 ( .A(_02487__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR35) );
  MUX2_X1 U26862 ( .A(_02487__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR36) );
  MUX2_X1 U26863 ( .A(_02487__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR37) );
  MUX2_X1 U26864 ( .A(_02487__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR38) );
  MUX2_X1 U26865 ( .A(_02487__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR39) );
  MUX2_X1 U26866 ( .A(_02487__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR64) );
  MUX2_X1 U26867 ( .A(_02487__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR65) );
  MUX2_X1 U26868 ( .A(_02487__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR66) );
  MUX2_X1 U26869 ( .A(_02487__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR67) );
  MUX2_X1 U26870 ( .A(_02487__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR68) );
  MUX2_X1 U26871 ( .A(_02487__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR69) );
  MUX2_X1 U26872 ( .A(_02487__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR70) );
  MUX2_X1 U26873 ( .A(_02487__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03366__PTR71) );
  MUX2_X1 U26874 ( .A(_03371__PTR0), .B(_03369__PTR64), .S(P3_P1_State2_PTR3), .Z(_02490__PTR0) );
  MUX2_X1 U26875 ( .A(_03371__PTR1), .B(_03369__PTR65), .S(P3_P1_State2_PTR3), .Z(_02490__PTR1) );
  MUX2_X1 U26876 ( .A(_03371__PTR2), .B(_03369__PTR66), .S(P3_P1_State2_PTR3), .Z(_02490__PTR2) );
  MUX2_X1 U26877 ( .A(_03371__PTR3), .B(_03369__PTR67), .S(P3_P1_State2_PTR3), .Z(_02490__PTR3) );
  MUX2_X1 U26878 ( .A(_03371__PTR4), .B(_03369__PTR68), .S(P3_P1_State2_PTR3), .Z(_02490__PTR4) );
  MUX2_X1 U26879 ( .A(_03371__PTR5), .B(_03369__PTR69), .S(P3_P1_State2_PTR3), .Z(_02490__PTR5) );
  MUX2_X1 U26880 ( .A(_03371__PTR6), .B(_03369__PTR70), .S(P3_P1_State2_PTR3), .Z(_02490__PTR6) );
  MUX2_X1 U26881 ( .A(_03371__PTR7), .B(_03369__PTR71), .S(P3_P1_State2_PTR3), .Z(_02490__PTR7) );
  MUX2_X1 U26882 ( .A(_03370__PTR0), .B(_03370__PTR32), .S(P3_P1_State2_PTR2), .Z(_03371__PTR0) );
  MUX2_X1 U26883 ( .A(_03370__PTR1), .B(_03370__PTR33), .S(P3_P1_State2_PTR2), .Z(_03371__PTR1) );
  MUX2_X1 U26884 ( .A(_03370__PTR2), .B(_03370__PTR34), .S(P3_P1_State2_PTR2), .Z(_03371__PTR2) );
  MUX2_X1 U26885 ( .A(_03370__PTR3), .B(_03370__PTR35), .S(P3_P1_State2_PTR2), .Z(_03371__PTR3) );
  MUX2_X1 U26886 ( .A(_03370__PTR4), .B(_03370__PTR36), .S(P3_P1_State2_PTR2), .Z(_03371__PTR4) );
  MUX2_X1 U26887 ( .A(_03370__PTR5), .B(_03370__PTR37), .S(P3_P1_State2_PTR2), .Z(_03371__PTR5) );
  MUX2_X1 U26888 ( .A(_03370__PTR6), .B(_03370__PTR38), .S(P3_P1_State2_PTR2), .Z(_03371__PTR6) );
  MUX2_X1 U26889 ( .A(_03370__PTR7), .B(_03370__PTR39), .S(P3_P1_State2_PTR2), .Z(_03371__PTR7) );
  MUX2_X1 U26890 ( .A(1'b0), .B(_03369__PTR16), .S(P3_P1_State2_PTR1), .Z(_03370__PTR0) );
  MUX2_X1 U26891 ( .A(1'b0), .B(_03369__PTR17), .S(P3_P1_State2_PTR1), .Z(_03370__PTR1) );
  MUX2_X1 U26892 ( .A(1'b0), .B(_03369__PTR18), .S(P3_P1_State2_PTR1), .Z(_03370__PTR2) );
  MUX2_X1 U26893 ( .A(1'b0), .B(_03369__PTR19), .S(P3_P1_State2_PTR1), .Z(_03370__PTR3) );
  MUX2_X1 U26894 ( .A(1'b0), .B(_03369__PTR20), .S(P3_P1_State2_PTR1), .Z(_03370__PTR4) );
  MUX2_X1 U26895 ( .A(1'b0), .B(_03369__PTR21), .S(P3_P1_State2_PTR1), .Z(_03370__PTR5) );
  MUX2_X1 U26896 ( .A(1'b0), .B(_03369__PTR22), .S(P3_P1_State2_PTR1), .Z(_03370__PTR6) );
  MUX2_X1 U26897 ( .A(1'b0), .B(_03369__PTR23), .S(P3_P1_State2_PTR1), .Z(_03370__PTR7) );
  MUX2_X1 U26898 ( .A(_03369__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03370__PTR32) );
  MUX2_X1 U26899 ( .A(_03369__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03370__PTR33) );
  MUX2_X1 U26900 ( .A(_03369__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03370__PTR34) );
  MUX2_X1 U26901 ( .A(_03369__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03370__PTR35) );
  MUX2_X1 U26902 ( .A(_03369__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03370__PTR36) );
  MUX2_X1 U26903 ( .A(_03369__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03370__PTR37) );
  MUX2_X1 U26904 ( .A(_03369__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03370__PTR38) );
  MUX2_X1 U26905 ( .A(_03369__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03370__PTR39) );
  MUX2_X1 U26906 ( .A(_02489__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR16) );
  MUX2_X1 U26907 ( .A(_02489__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR17) );
  MUX2_X1 U26908 ( .A(_02489__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR18) );
  MUX2_X1 U26909 ( .A(_02489__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR19) );
  MUX2_X1 U26910 ( .A(_02489__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR20) );
  MUX2_X1 U26911 ( .A(_02489__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR21) );
  MUX2_X1 U26912 ( .A(_02489__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR22) );
  MUX2_X1 U26913 ( .A(_02489__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR23) );
  MUX2_X1 U26914 ( .A(_02489__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR32) );
  MUX2_X1 U26915 ( .A(_02489__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR33) );
  MUX2_X1 U26916 ( .A(_02489__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR34) );
  MUX2_X1 U26917 ( .A(_02489__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR35) );
  MUX2_X1 U26918 ( .A(_02489__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR36) );
  MUX2_X1 U26919 ( .A(_02489__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR37) );
  MUX2_X1 U26920 ( .A(_02489__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR38) );
  MUX2_X1 U26921 ( .A(_02489__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR39) );
  MUX2_X1 U26922 ( .A(_02489__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR64) );
  MUX2_X1 U26923 ( .A(_02489__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR65) );
  MUX2_X1 U26924 ( .A(_02489__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR66) );
  MUX2_X1 U26925 ( .A(_02489__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR67) );
  MUX2_X1 U26926 ( .A(_02489__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR68) );
  MUX2_X1 U26927 ( .A(_02489__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR69) );
  MUX2_X1 U26928 ( .A(_02489__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR70) );
  MUX2_X1 U26929 ( .A(_02489__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03369__PTR71) );
  MUX2_X1 U26930 ( .A(_03374__PTR0), .B(_03372__PTR64), .S(P3_P1_State2_PTR3), .Z(_02492__PTR0) );
  MUX2_X1 U26931 ( .A(_03374__PTR1), .B(_03372__PTR65), .S(P3_P1_State2_PTR3), .Z(_02492__PTR1) );
  MUX2_X1 U26932 ( .A(_03374__PTR2), .B(_03372__PTR66), .S(P3_P1_State2_PTR3), .Z(_02492__PTR2) );
  MUX2_X1 U26933 ( .A(_03374__PTR3), .B(_03372__PTR67), .S(P3_P1_State2_PTR3), .Z(_02492__PTR3) );
  MUX2_X1 U26934 ( .A(_03374__PTR4), .B(_03372__PTR68), .S(P3_P1_State2_PTR3), .Z(_02492__PTR4) );
  MUX2_X1 U26935 ( .A(_03374__PTR5), .B(_03372__PTR69), .S(P3_P1_State2_PTR3), .Z(_02492__PTR5) );
  MUX2_X1 U26936 ( .A(_03374__PTR6), .B(_03372__PTR70), .S(P3_P1_State2_PTR3), .Z(_02492__PTR6) );
  MUX2_X1 U26937 ( .A(_03374__PTR7), .B(_03372__PTR71), .S(P3_P1_State2_PTR3), .Z(_02492__PTR7) );
  MUX2_X1 U26938 ( .A(_03373__PTR0), .B(_03373__PTR32), .S(P3_P1_State2_PTR2), .Z(_03374__PTR0) );
  MUX2_X1 U26939 ( .A(_03373__PTR1), .B(_03373__PTR33), .S(P3_P1_State2_PTR2), .Z(_03374__PTR1) );
  MUX2_X1 U26940 ( .A(_03373__PTR2), .B(_03373__PTR34), .S(P3_P1_State2_PTR2), .Z(_03374__PTR2) );
  MUX2_X1 U26941 ( .A(_03373__PTR3), .B(_03373__PTR35), .S(P3_P1_State2_PTR2), .Z(_03374__PTR3) );
  MUX2_X1 U26942 ( .A(_03373__PTR4), .B(_03373__PTR36), .S(P3_P1_State2_PTR2), .Z(_03374__PTR4) );
  MUX2_X1 U26943 ( .A(_03373__PTR5), .B(_03373__PTR37), .S(P3_P1_State2_PTR2), .Z(_03374__PTR5) );
  MUX2_X1 U26944 ( .A(_03373__PTR6), .B(_03373__PTR38), .S(P3_P1_State2_PTR2), .Z(_03374__PTR6) );
  MUX2_X1 U26945 ( .A(_03373__PTR7), .B(_03373__PTR39), .S(P3_P1_State2_PTR2), .Z(_03374__PTR7) );
  MUX2_X1 U26946 ( .A(1'b0), .B(_03372__PTR16), .S(P3_P1_State2_PTR1), .Z(_03373__PTR0) );
  MUX2_X1 U26947 ( .A(1'b0), .B(_03372__PTR17), .S(P3_P1_State2_PTR1), .Z(_03373__PTR1) );
  MUX2_X1 U26948 ( .A(1'b0), .B(_03372__PTR18), .S(P3_P1_State2_PTR1), .Z(_03373__PTR2) );
  MUX2_X1 U26949 ( .A(1'b0), .B(_03372__PTR19), .S(P3_P1_State2_PTR1), .Z(_03373__PTR3) );
  MUX2_X1 U26950 ( .A(1'b0), .B(_03372__PTR20), .S(P3_P1_State2_PTR1), .Z(_03373__PTR4) );
  MUX2_X1 U26951 ( .A(1'b0), .B(_03372__PTR21), .S(P3_P1_State2_PTR1), .Z(_03373__PTR5) );
  MUX2_X1 U26952 ( .A(1'b0), .B(_03372__PTR22), .S(P3_P1_State2_PTR1), .Z(_03373__PTR6) );
  MUX2_X1 U26953 ( .A(1'b0), .B(_03372__PTR23), .S(P3_P1_State2_PTR1), .Z(_03373__PTR7) );
  MUX2_X1 U26954 ( .A(_03372__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03373__PTR32) );
  MUX2_X1 U26955 ( .A(_03372__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03373__PTR33) );
  MUX2_X1 U26956 ( .A(_03372__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03373__PTR34) );
  MUX2_X1 U26957 ( .A(_03372__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03373__PTR35) );
  MUX2_X1 U26958 ( .A(_03372__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03373__PTR36) );
  MUX2_X1 U26959 ( .A(_03372__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03373__PTR37) );
  MUX2_X1 U26960 ( .A(_03372__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03373__PTR38) );
  MUX2_X1 U26961 ( .A(_03372__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03373__PTR39) );
  MUX2_X1 U26962 ( .A(_02491__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR16) );
  MUX2_X1 U26963 ( .A(_02491__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR17) );
  MUX2_X1 U26964 ( .A(_02491__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR18) );
  MUX2_X1 U26965 ( .A(_02491__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR19) );
  MUX2_X1 U26966 ( .A(_02491__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR20) );
  MUX2_X1 U26967 ( .A(_02491__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR21) );
  MUX2_X1 U26968 ( .A(_02491__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR22) );
  MUX2_X1 U26969 ( .A(_02491__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR23) );
  MUX2_X1 U26970 ( .A(_02491__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR32) );
  MUX2_X1 U26971 ( .A(_02491__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR33) );
  MUX2_X1 U26972 ( .A(_02491__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR34) );
  MUX2_X1 U26973 ( .A(_02491__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR35) );
  MUX2_X1 U26974 ( .A(_02491__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR36) );
  MUX2_X1 U26975 ( .A(_02491__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR37) );
  MUX2_X1 U26976 ( .A(_02491__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR38) );
  MUX2_X1 U26977 ( .A(_02491__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR39) );
  MUX2_X1 U26978 ( .A(_02491__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR64) );
  MUX2_X1 U26979 ( .A(_02491__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR65) );
  MUX2_X1 U26980 ( .A(_02491__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR66) );
  MUX2_X1 U26981 ( .A(_02491__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR67) );
  MUX2_X1 U26982 ( .A(_02491__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR68) );
  MUX2_X1 U26983 ( .A(_02491__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR69) );
  MUX2_X1 U26984 ( .A(_02491__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR70) );
  MUX2_X1 U26985 ( .A(_02491__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03372__PTR71) );
  MUX2_X1 U26986 ( .A(_03377__PTR0), .B(_03375__PTR64), .S(P3_P1_State2_PTR3), .Z(_02494__PTR0) );
  MUX2_X1 U26987 ( .A(_03377__PTR1), .B(_03375__PTR65), .S(P3_P1_State2_PTR3), .Z(_02494__PTR1) );
  MUX2_X1 U26988 ( .A(_03377__PTR2), .B(_03375__PTR66), .S(P3_P1_State2_PTR3), .Z(_02494__PTR2) );
  MUX2_X1 U26989 ( .A(_03377__PTR3), .B(_03375__PTR67), .S(P3_P1_State2_PTR3), .Z(_02494__PTR3) );
  MUX2_X1 U26990 ( .A(_03377__PTR4), .B(_03375__PTR68), .S(P3_P1_State2_PTR3), .Z(_02494__PTR4) );
  MUX2_X1 U26991 ( .A(_03377__PTR5), .B(_03375__PTR69), .S(P3_P1_State2_PTR3), .Z(_02494__PTR5) );
  MUX2_X1 U26992 ( .A(_03377__PTR6), .B(_03375__PTR70), .S(P3_P1_State2_PTR3), .Z(_02494__PTR6) );
  MUX2_X1 U26993 ( .A(_03377__PTR7), .B(_03375__PTR71), .S(P3_P1_State2_PTR3), .Z(_02494__PTR7) );
  MUX2_X1 U26994 ( .A(_03376__PTR0), .B(_03376__PTR32), .S(P3_P1_State2_PTR2), .Z(_03377__PTR0) );
  MUX2_X1 U26995 ( .A(_03376__PTR1), .B(_03376__PTR33), .S(P3_P1_State2_PTR2), .Z(_03377__PTR1) );
  MUX2_X1 U26996 ( .A(_03376__PTR2), .B(_03376__PTR34), .S(P3_P1_State2_PTR2), .Z(_03377__PTR2) );
  MUX2_X1 U26997 ( .A(_03376__PTR3), .B(_03376__PTR35), .S(P3_P1_State2_PTR2), .Z(_03377__PTR3) );
  MUX2_X1 U26998 ( .A(_03376__PTR4), .B(_03376__PTR36), .S(P3_P1_State2_PTR2), .Z(_03377__PTR4) );
  MUX2_X1 U26999 ( .A(_03376__PTR5), .B(_03376__PTR37), .S(P3_P1_State2_PTR2), .Z(_03377__PTR5) );
  MUX2_X1 U27000 ( .A(_03376__PTR6), .B(_03376__PTR38), .S(P3_P1_State2_PTR2), .Z(_03377__PTR6) );
  MUX2_X1 U27001 ( .A(_03376__PTR7), .B(_03376__PTR39), .S(P3_P1_State2_PTR2), .Z(_03377__PTR7) );
  MUX2_X1 U27002 ( .A(1'b0), .B(_03375__PTR16), .S(P3_P1_State2_PTR1), .Z(_03376__PTR0) );
  MUX2_X1 U27003 ( .A(1'b0), .B(_03375__PTR17), .S(P3_P1_State2_PTR1), .Z(_03376__PTR1) );
  MUX2_X1 U27004 ( .A(1'b0), .B(_03375__PTR18), .S(P3_P1_State2_PTR1), .Z(_03376__PTR2) );
  MUX2_X1 U27005 ( .A(1'b0), .B(_03375__PTR19), .S(P3_P1_State2_PTR1), .Z(_03376__PTR3) );
  MUX2_X1 U27006 ( .A(1'b0), .B(_03375__PTR20), .S(P3_P1_State2_PTR1), .Z(_03376__PTR4) );
  MUX2_X1 U27007 ( .A(1'b0), .B(_03375__PTR21), .S(P3_P1_State2_PTR1), .Z(_03376__PTR5) );
  MUX2_X1 U27008 ( .A(1'b0), .B(_03375__PTR22), .S(P3_P1_State2_PTR1), .Z(_03376__PTR6) );
  MUX2_X1 U27009 ( .A(1'b0), .B(_03375__PTR23), .S(P3_P1_State2_PTR1), .Z(_03376__PTR7) );
  MUX2_X1 U27010 ( .A(_03375__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03376__PTR32) );
  MUX2_X1 U27011 ( .A(_03375__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03376__PTR33) );
  MUX2_X1 U27012 ( .A(_03375__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03376__PTR34) );
  MUX2_X1 U27013 ( .A(_03375__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03376__PTR35) );
  MUX2_X1 U27014 ( .A(_03375__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03376__PTR36) );
  MUX2_X1 U27015 ( .A(_03375__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03376__PTR37) );
  MUX2_X1 U27016 ( .A(_03375__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03376__PTR38) );
  MUX2_X1 U27017 ( .A(_03375__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03376__PTR39) );
  MUX2_X1 U27018 ( .A(_02493__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR16) );
  MUX2_X1 U27019 ( .A(_02493__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR17) );
  MUX2_X1 U27020 ( .A(_02493__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR18) );
  MUX2_X1 U27021 ( .A(_02493__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR19) );
  MUX2_X1 U27022 ( .A(_02493__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR20) );
  MUX2_X1 U27023 ( .A(_02493__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR21) );
  MUX2_X1 U27024 ( .A(_02493__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR22) );
  MUX2_X1 U27025 ( .A(_02493__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR23) );
  MUX2_X1 U27026 ( .A(_02493__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR32) );
  MUX2_X1 U27027 ( .A(_02493__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR33) );
  MUX2_X1 U27028 ( .A(_02493__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR34) );
  MUX2_X1 U27029 ( .A(_02493__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR35) );
  MUX2_X1 U27030 ( .A(_02493__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR36) );
  MUX2_X1 U27031 ( .A(_02493__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR37) );
  MUX2_X1 U27032 ( .A(_02493__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR38) );
  MUX2_X1 U27033 ( .A(_02493__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR39) );
  MUX2_X1 U27034 ( .A(_02493__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR64) );
  MUX2_X1 U27035 ( .A(_02493__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR65) );
  MUX2_X1 U27036 ( .A(_02493__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR66) );
  MUX2_X1 U27037 ( .A(_02493__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR67) );
  MUX2_X1 U27038 ( .A(_02493__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR68) );
  MUX2_X1 U27039 ( .A(_02493__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR69) );
  MUX2_X1 U27040 ( .A(_02493__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR70) );
  MUX2_X1 U27041 ( .A(_02493__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03375__PTR71) );
  MUX2_X1 U27042 ( .A(_03380__PTR0), .B(_03378__PTR64), .S(P3_P1_State2_PTR3), .Z(_02496__PTR0) );
  MUX2_X1 U27043 ( .A(_03380__PTR1), .B(_03378__PTR65), .S(P3_P1_State2_PTR3), .Z(_02496__PTR1) );
  MUX2_X1 U27044 ( .A(_03380__PTR2), .B(_03378__PTR66), .S(P3_P1_State2_PTR3), .Z(_02496__PTR2) );
  MUX2_X1 U27045 ( .A(_03380__PTR3), .B(_03378__PTR67), .S(P3_P1_State2_PTR3), .Z(_02496__PTR3) );
  MUX2_X1 U27046 ( .A(_03380__PTR4), .B(_03378__PTR68), .S(P3_P1_State2_PTR3), .Z(_02496__PTR4) );
  MUX2_X1 U27047 ( .A(_03380__PTR5), .B(_03378__PTR69), .S(P3_P1_State2_PTR3), .Z(_02496__PTR5) );
  MUX2_X1 U27048 ( .A(_03380__PTR6), .B(_03378__PTR70), .S(P3_P1_State2_PTR3), .Z(_02496__PTR6) );
  MUX2_X1 U27049 ( .A(_03380__PTR7), .B(_03378__PTR71), .S(P3_P1_State2_PTR3), .Z(_02496__PTR7) );
  MUX2_X1 U27050 ( .A(_03379__PTR0), .B(_03379__PTR32), .S(P3_P1_State2_PTR2), .Z(_03380__PTR0) );
  MUX2_X1 U27051 ( .A(_03379__PTR1), .B(_03379__PTR33), .S(P3_P1_State2_PTR2), .Z(_03380__PTR1) );
  MUX2_X1 U27052 ( .A(_03379__PTR2), .B(_03379__PTR34), .S(P3_P1_State2_PTR2), .Z(_03380__PTR2) );
  MUX2_X1 U27053 ( .A(_03379__PTR3), .B(_03379__PTR35), .S(P3_P1_State2_PTR2), .Z(_03380__PTR3) );
  MUX2_X1 U27054 ( .A(_03379__PTR4), .B(_03379__PTR36), .S(P3_P1_State2_PTR2), .Z(_03380__PTR4) );
  MUX2_X1 U27055 ( .A(_03379__PTR5), .B(_03379__PTR37), .S(P3_P1_State2_PTR2), .Z(_03380__PTR5) );
  MUX2_X1 U27056 ( .A(_03379__PTR6), .B(_03379__PTR38), .S(P3_P1_State2_PTR2), .Z(_03380__PTR6) );
  MUX2_X1 U27057 ( .A(_03379__PTR7), .B(_03379__PTR39), .S(P3_P1_State2_PTR2), .Z(_03380__PTR7) );
  MUX2_X1 U27058 ( .A(1'b0), .B(_03378__PTR16), .S(P3_P1_State2_PTR1), .Z(_03379__PTR0) );
  MUX2_X1 U27059 ( .A(1'b0), .B(_03378__PTR17), .S(P3_P1_State2_PTR1), .Z(_03379__PTR1) );
  MUX2_X1 U27060 ( .A(1'b0), .B(_03378__PTR18), .S(P3_P1_State2_PTR1), .Z(_03379__PTR2) );
  MUX2_X1 U27061 ( .A(1'b0), .B(_03378__PTR19), .S(P3_P1_State2_PTR1), .Z(_03379__PTR3) );
  MUX2_X1 U27062 ( .A(1'b0), .B(_03378__PTR20), .S(P3_P1_State2_PTR1), .Z(_03379__PTR4) );
  MUX2_X1 U27063 ( .A(1'b0), .B(_03378__PTR21), .S(P3_P1_State2_PTR1), .Z(_03379__PTR5) );
  MUX2_X1 U27064 ( .A(1'b0), .B(_03378__PTR22), .S(P3_P1_State2_PTR1), .Z(_03379__PTR6) );
  MUX2_X1 U27065 ( .A(1'b0), .B(_03378__PTR23), .S(P3_P1_State2_PTR1), .Z(_03379__PTR7) );
  MUX2_X1 U27066 ( .A(_03378__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03379__PTR32) );
  MUX2_X1 U27067 ( .A(_03378__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03379__PTR33) );
  MUX2_X1 U27068 ( .A(_03378__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03379__PTR34) );
  MUX2_X1 U27069 ( .A(_03378__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03379__PTR35) );
  MUX2_X1 U27070 ( .A(_03378__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03379__PTR36) );
  MUX2_X1 U27071 ( .A(_03378__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03379__PTR37) );
  MUX2_X1 U27072 ( .A(_03378__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03379__PTR38) );
  MUX2_X1 U27073 ( .A(_03378__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03379__PTR39) );
  MUX2_X1 U27074 ( .A(_02495__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR16) );
  MUX2_X1 U27075 ( .A(_02495__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR17) );
  MUX2_X1 U27076 ( .A(_02495__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR18) );
  MUX2_X1 U27077 ( .A(_02495__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR19) );
  MUX2_X1 U27078 ( .A(_02495__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR20) );
  MUX2_X1 U27079 ( .A(_02495__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR21) );
  MUX2_X1 U27080 ( .A(_02495__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR22) );
  MUX2_X1 U27081 ( .A(_02495__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR23) );
  MUX2_X1 U27082 ( .A(_02495__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR32) );
  MUX2_X1 U27083 ( .A(_02495__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR33) );
  MUX2_X1 U27084 ( .A(_02495__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR34) );
  MUX2_X1 U27085 ( .A(_02495__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR35) );
  MUX2_X1 U27086 ( .A(_02495__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR36) );
  MUX2_X1 U27087 ( .A(_02495__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR37) );
  MUX2_X1 U27088 ( .A(_02495__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR38) );
  MUX2_X1 U27089 ( .A(_02495__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR39) );
  MUX2_X1 U27090 ( .A(_02495__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR64) );
  MUX2_X1 U27091 ( .A(_02495__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR65) );
  MUX2_X1 U27092 ( .A(_02495__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR66) );
  MUX2_X1 U27093 ( .A(_02495__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR67) );
  MUX2_X1 U27094 ( .A(_02495__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR68) );
  MUX2_X1 U27095 ( .A(_02495__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR69) );
  MUX2_X1 U27096 ( .A(_02495__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR70) );
  MUX2_X1 U27097 ( .A(_02495__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03378__PTR71) );
  MUX2_X1 U27098 ( .A(_03383__PTR0), .B(_03381__PTR64), .S(P3_P1_State2_PTR3), .Z(_02498__PTR0) );
  MUX2_X1 U27099 ( .A(_03383__PTR1), .B(_03381__PTR65), .S(P3_P1_State2_PTR3), .Z(_02498__PTR1) );
  MUX2_X1 U27100 ( .A(_03383__PTR2), .B(_03381__PTR66), .S(P3_P1_State2_PTR3), .Z(_02498__PTR2) );
  MUX2_X1 U27101 ( .A(_03383__PTR3), .B(_03381__PTR67), .S(P3_P1_State2_PTR3), .Z(_02498__PTR3) );
  MUX2_X1 U27102 ( .A(_03383__PTR4), .B(_03381__PTR68), .S(P3_P1_State2_PTR3), .Z(_02498__PTR4) );
  MUX2_X1 U27103 ( .A(_03383__PTR5), .B(_03381__PTR69), .S(P3_P1_State2_PTR3), .Z(_02498__PTR5) );
  MUX2_X1 U27104 ( .A(_03383__PTR6), .B(_03381__PTR70), .S(P3_P1_State2_PTR3), .Z(_02498__PTR6) );
  MUX2_X1 U27105 ( .A(_03383__PTR7), .B(_03381__PTR71), .S(P3_P1_State2_PTR3), .Z(_02498__PTR7) );
  MUX2_X1 U27106 ( .A(_03382__PTR0), .B(_03382__PTR32), .S(P3_P1_State2_PTR2), .Z(_03383__PTR0) );
  MUX2_X1 U27107 ( .A(_03382__PTR1), .B(_03382__PTR33), .S(P3_P1_State2_PTR2), .Z(_03383__PTR1) );
  MUX2_X1 U27108 ( .A(_03382__PTR2), .B(_03382__PTR34), .S(P3_P1_State2_PTR2), .Z(_03383__PTR2) );
  MUX2_X1 U27109 ( .A(_03382__PTR3), .B(_03382__PTR35), .S(P3_P1_State2_PTR2), .Z(_03383__PTR3) );
  MUX2_X1 U27110 ( .A(_03382__PTR4), .B(_03382__PTR36), .S(P3_P1_State2_PTR2), .Z(_03383__PTR4) );
  MUX2_X1 U27111 ( .A(_03382__PTR5), .B(_03382__PTR37), .S(P3_P1_State2_PTR2), .Z(_03383__PTR5) );
  MUX2_X1 U27112 ( .A(_03382__PTR6), .B(_03382__PTR38), .S(P3_P1_State2_PTR2), .Z(_03383__PTR6) );
  MUX2_X1 U27113 ( .A(_03382__PTR7), .B(_03382__PTR39), .S(P3_P1_State2_PTR2), .Z(_03383__PTR7) );
  MUX2_X1 U27114 ( .A(1'b0), .B(_03381__PTR16), .S(P3_P1_State2_PTR1), .Z(_03382__PTR0) );
  MUX2_X1 U27115 ( .A(1'b0), .B(_03381__PTR17), .S(P3_P1_State2_PTR1), .Z(_03382__PTR1) );
  MUX2_X1 U27116 ( .A(1'b0), .B(_03381__PTR18), .S(P3_P1_State2_PTR1), .Z(_03382__PTR2) );
  MUX2_X1 U27117 ( .A(1'b0), .B(_03381__PTR19), .S(P3_P1_State2_PTR1), .Z(_03382__PTR3) );
  MUX2_X1 U27118 ( .A(1'b0), .B(_03381__PTR20), .S(P3_P1_State2_PTR1), .Z(_03382__PTR4) );
  MUX2_X1 U27119 ( .A(1'b0), .B(_03381__PTR21), .S(P3_P1_State2_PTR1), .Z(_03382__PTR5) );
  MUX2_X1 U27120 ( .A(1'b0), .B(_03381__PTR22), .S(P3_P1_State2_PTR1), .Z(_03382__PTR6) );
  MUX2_X1 U27121 ( .A(1'b0), .B(_03381__PTR23), .S(P3_P1_State2_PTR1), .Z(_03382__PTR7) );
  MUX2_X1 U27122 ( .A(_03381__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03382__PTR32) );
  MUX2_X1 U27123 ( .A(_03381__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03382__PTR33) );
  MUX2_X1 U27124 ( .A(_03381__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03382__PTR34) );
  MUX2_X1 U27125 ( .A(_03381__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03382__PTR35) );
  MUX2_X1 U27126 ( .A(_03381__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03382__PTR36) );
  MUX2_X1 U27127 ( .A(_03381__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03382__PTR37) );
  MUX2_X1 U27128 ( .A(_03381__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03382__PTR38) );
  MUX2_X1 U27129 ( .A(_03381__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03382__PTR39) );
  MUX2_X1 U27130 ( .A(_02497__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR16) );
  MUX2_X1 U27131 ( .A(_02497__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR17) );
  MUX2_X1 U27132 ( .A(_02497__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR18) );
  MUX2_X1 U27133 ( .A(_02497__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR19) );
  MUX2_X1 U27134 ( .A(_02497__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR20) );
  MUX2_X1 U27135 ( .A(_02497__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR21) );
  MUX2_X1 U27136 ( .A(_02497__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR22) );
  MUX2_X1 U27137 ( .A(_02497__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR23) );
  MUX2_X1 U27138 ( .A(_02497__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR32) );
  MUX2_X1 U27139 ( .A(_02497__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR33) );
  MUX2_X1 U27140 ( .A(_02497__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR34) );
  MUX2_X1 U27141 ( .A(_02497__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR35) );
  MUX2_X1 U27142 ( .A(_02497__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR36) );
  MUX2_X1 U27143 ( .A(_02497__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR37) );
  MUX2_X1 U27144 ( .A(_02497__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR38) );
  MUX2_X1 U27145 ( .A(_02497__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR39) );
  MUX2_X1 U27146 ( .A(_02497__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR64) );
  MUX2_X1 U27147 ( .A(_02497__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR65) );
  MUX2_X1 U27148 ( .A(_02497__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR66) );
  MUX2_X1 U27149 ( .A(_02497__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR67) );
  MUX2_X1 U27150 ( .A(_02497__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR68) );
  MUX2_X1 U27151 ( .A(_02497__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR69) );
  MUX2_X1 U27152 ( .A(_02497__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR70) );
  MUX2_X1 U27153 ( .A(_02497__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03381__PTR71) );
  MUX2_X1 U27154 ( .A(_03386__PTR0), .B(_03384__PTR64), .S(P3_P1_State2_PTR3), .Z(_02500__PTR0) );
  MUX2_X1 U27155 ( .A(_03386__PTR1), .B(_03384__PTR65), .S(P3_P1_State2_PTR3), .Z(_02500__PTR1) );
  MUX2_X1 U27156 ( .A(_03386__PTR2), .B(_03384__PTR66), .S(P3_P1_State2_PTR3), .Z(_02500__PTR2) );
  MUX2_X1 U27157 ( .A(_03386__PTR3), .B(_03384__PTR67), .S(P3_P1_State2_PTR3), .Z(_02500__PTR3) );
  MUX2_X1 U27158 ( .A(_03386__PTR4), .B(_03384__PTR68), .S(P3_P1_State2_PTR3), .Z(_02500__PTR4) );
  MUX2_X1 U27159 ( .A(_03386__PTR5), .B(_03384__PTR69), .S(P3_P1_State2_PTR3), .Z(_02500__PTR5) );
  MUX2_X1 U27160 ( .A(_03386__PTR6), .B(_03384__PTR70), .S(P3_P1_State2_PTR3), .Z(_02500__PTR6) );
  MUX2_X1 U27161 ( .A(_03386__PTR7), .B(_03384__PTR71), .S(P3_P1_State2_PTR3), .Z(_02500__PTR7) );
  MUX2_X1 U27162 ( .A(_03385__PTR0), .B(_03385__PTR32), .S(P3_P1_State2_PTR2), .Z(_03386__PTR0) );
  MUX2_X1 U27163 ( .A(_03385__PTR1), .B(_03385__PTR33), .S(P3_P1_State2_PTR2), .Z(_03386__PTR1) );
  MUX2_X1 U27164 ( .A(_03385__PTR2), .B(_03385__PTR34), .S(P3_P1_State2_PTR2), .Z(_03386__PTR2) );
  MUX2_X1 U27165 ( .A(_03385__PTR3), .B(_03385__PTR35), .S(P3_P1_State2_PTR2), .Z(_03386__PTR3) );
  MUX2_X1 U27166 ( .A(_03385__PTR4), .B(_03385__PTR36), .S(P3_P1_State2_PTR2), .Z(_03386__PTR4) );
  MUX2_X1 U27167 ( .A(_03385__PTR5), .B(_03385__PTR37), .S(P3_P1_State2_PTR2), .Z(_03386__PTR5) );
  MUX2_X1 U27168 ( .A(_03385__PTR6), .B(_03385__PTR38), .S(P3_P1_State2_PTR2), .Z(_03386__PTR6) );
  MUX2_X1 U27169 ( .A(_03385__PTR7), .B(_03385__PTR39), .S(P3_P1_State2_PTR2), .Z(_03386__PTR7) );
  MUX2_X1 U27170 ( .A(1'b0), .B(_03384__PTR16), .S(P3_P1_State2_PTR1), .Z(_03385__PTR0) );
  MUX2_X1 U27171 ( .A(1'b0), .B(_03384__PTR17), .S(P3_P1_State2_PTR1), .Z(_03385__PTR1) );
  MUX2_X1 U27172 ( .A(1'b0), .B(_03384__PTR18), .S(P3_P1_State2_PTR1), .Z(_03385__PTR2) );
  MUX2_X1 U27173 ( .A(1'b0), .B(_03384__PTR19), .S(P3_P1_State2_PTR1), .Z(_03385__PTR3) );
  MUX2_X1 U27174 ( .A(1'b0), .B(_03384__PTR20), .S(P3_P1_State2_PTR1), .Z(_03385__PTR4) );
  MUX2_X1 U27175 ( .A(1'b0), .B(_03384__PTR21), .S(P3_P1_State2_PTR1), .Z(_03385__PTR5) );
  MUX2_X1 U27176 ( .A(1'b0), .B(_03384__PTR22), .S(P3_P1_State2_PTR1), .Z(_03385__PTR6) );
  MUX2_X1 U27177 ( .A(1'b0), .B(_03384__PTR23), .S(P3_P1_State2_PTR1), .Z(_03385__PTR7) );
  MUX2_X1 U27178 ( .A(_03384__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03385__PTR32) );
  MUX2_X1 U27179 ( .A(_03384__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03385__PTR33) );
  MUX2_X1 U27180 ( .A(_03384__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03385__PTR34) );
  MUX2_X1 U27181 ( .A(_03384__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03385__PTR35) );
  MUX2_X1 U27182 ( .A(_03384__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03385__PTR36) );
  MUX2_X1 U27183 ( .A(_03384__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03385__PTR37) );
  MUX2_X1 U27184 ( .A(_03384__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03385__PTR38) );
  MUX2_X1 U27185 ( .A(_03384__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03385__PTR39) );
  MUX2_X1 U27186 ( .A(_02499__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR16) );
  MUX2_X1 U27187 ( .A(_02499__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR17) );
  MUX2_X1 U27188 ( .A(_02499__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR18) );
  MUX2_X1 U27189 ( .A(_02499__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR19) );
  MUX2_X1 U27190 ( .A(_02499__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR20) );
  MUX2_X1 U27191 ( .A(_02499__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR21) );
  MUX2_X1 U27192 ( .A(_02499__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR22) );
  MUX2_X1 U27193 ( .A(_02499__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR23) );
  MUX2_X1 U27194 ( .A(_02499__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR32) );
  MUX2_X1 U27195 ( .A(_02499__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR33) );
  MUX2_X1 U27196 ( .A(_02499__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR34) );
  MUX2_X1 U27197 ( .A(_02499__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR35) );
  MUX2_X1 U27198 ( .A(_02499__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR36) );
  MUX2_X1 U27199 ( .A(_02499__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR37) );
  MUX2_X1 U27200 ( .A(_02499__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR38) );
  MUX2_X1 U27201 ( .A(_02499__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR39) );
  MUX2_X1 U27202 ( .A(_02499__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR64) );
  MUX2_X1 U27203 ( .A(_02499__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR65) );
  MUX2_X1 U27204 ( .A(_02499__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR66) );
  MUX2_X1 U27205 ( .A(_02499__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR67) );
  MUX2_X1 U27206 ( .A(_02499__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR68) );
  MUX2_X1 U27207 ( .A(_02499__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR69) );
  MUX2_X1 U27208 ( .A(_02499__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR70) );
  MUX2_X1 U27209 ( .A(_02499__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03384__PTR71) );
  MUX2_X1 U27210 ( .A(_03389__PTR0), .B(_03387__PTR64), .S(P3_P1_State2_PTR3), .Z(_02502__PTR0) );
  MUX2_X1 U27211 ( .A(_03389__PTR1), .B(_03387__PTR65), .S(P3_P1_State2_PTR3), .Z(_02502__PTR1) );
  MUX2_X1 U27212 ( .A(_03389__PTR2), .B(_03387__PTR66), .S(P3_P1_State2_PTR3), .Z(_02502__PTR2) );
  MUX2_X1 U27213 ( .A(_03389__PTR3), .B(_03387__PTR67), .S(P3_P1_State2_PTR3), .Z(_02502__PTR3) );
  MUX2_X1 U27214 ( .A(_03389__PTR4), .B(_03387__PTR68), .S(P3_P1_State2_PTR3), .Z(_02502__PTR4) );
  MUX2_X1 U27215 ( .A(_03389__PTR5), .B(_03387__PTR69), .S(P3_P1_State2_PTR3), .Z(_02502__PTR5) );
  MUX2_X1 U27216 ( .A(_03389__PTR6), .B(_03387__PTR70), .S(P3_P1_State2_PTR3), .Z(_02502__PTR6) );
  MUX2_X1 U27217 ( .A(_03389__PTR7), .B(_03387__PTR71), .S(P3_P1_State2_PTR3), .Z(_02502__PTR7) );
  MUX2_X1 U27218 ( .A(_03388__PTR0), .B(_03388__PTR32), .S(P3_P1_State2_PTR2), .Z(_03389__PTR0) );
  MUX2_X1 U27219 ( .A(_03388__PTR1), .B(_03388__PTR33), .S(P3_P1_State2_PTR2), .Z(_03389__PTR1) );
  MUX2_X1 U27220 ( .A(_03388__PTR2), .B(_03388__PTR34), .S(P3_P1_State2_PTR2), .Z(_03389__PTR2) );
  MUX2_X1 U27221 ( .A(_03388__PTR3), .B(_03388__PTR35), .S(P3_P1_State2_PTR2), .Z(_03389__PTR3) );
  MUX2_X1 U27222 ( .A(_03388__PTR4), .B(_03388__PTR36), .S(P3_P1_State2_PTR2), .Z(_03389__PTR4) );
  MUX2_X1 U27223 ( .A(_03388__PTR5), .B(_03388__PTR37), .S(P3_P1_State2_PTR2), .Z(_03389__PTR5) );
  MUX2_X1 U27224 ( .A(_03388__PTR6), .B(_03388__PTR38), .S(P3_P1_State2_PTR2), .Z(_03389__PTR6) );
  MUX2_X1 U27225 ( .A(_03388__PTR7), .B(_03388__PTR39), .S(P3_P1_State2_PTR2), .Z(_03389__PTR7) );
  MUX2_X1 U27226 ( .A(1'b0), .B(_03387__PTR16), .S(P3_P1_State2_PTR1), .Z(_03388__PTR0) );
  MUX2_X1 U27227 ( .A(1'b0), .B(_03387__PTR17), .S(P3_P1_State2_PTR1), .Z(_03388__PTR1) );
  MUX2_X1 U27228 ( .A(1'b0), .B(_03387__PTR18), .S(P3_P1_State2_PTR1), .Z(_03388__PTR2) );
  MUX2_X1 U27229 ( .A(1'b0), .B(_03387__PTR19), .S(P3_P1_State2_PTR1), .Z(_03388__PTR3) );
  MUX2_X1 U27230 ( .A(1'b0), .B(_03387__PTR20), .S(P3_P1_State2_PTR1), .Z(_03388__PTR4) );
  MUX2_X1 U27231 ( .A(1'b0), .B(_03387__PTR21), .S(P3_P1_State2_PTR1), .Z(_03388__PTR5) );
  MUX2_X1 U27232 ( .A(1'b0), .B(_03387__PTR22), .S(P3_P1_State2_PTR1), .Z(_03388__PTR6) );
  MUX2_X1 U27233 ( .A(1'b0), .B(_03387__PTR23), .S(P3_P1_State2_PTR1), .Z(_03388__PTR7) );
  MUX2_X1 U27234 ( .A(_03387__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03388__PTR32) );
  MUX2_X1 U27235 ( .A(_03387__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03388__PTR33) );
  MUX2_X1 U27236 ( .A(_03387__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03388__PTR34) );
  MUX2_X1 U27237 ( .A(_03387__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03388__PTR35) );
  MUX2_X1 U27238 ( .A(_03387__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03388__PTR36) );
  MUX2_X1 U27239 ( .A(_03387__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03388__PTR37) );
  MUX2_X1 U27240 ( .A(_03387__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03388__PTR38) );
  MUX2_X1 U27241 ( .A(_03387__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03388__PTR39) );
  MUX2_X1 U27242 ( .A(_02501__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR16) );
  MUX2_X1 U27243 ( .A(_02501__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR17) );
  MUX2_X1 U27244 ( .A(_02501__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR18) );
  MUX2_X1 U27245 ( .A(_02501__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR19) );
  MUX2_X1 U27246 ( .A(_02501__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR20) );
  MUX2_X1 U27247 ( .A(_02501__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR21) );
  MUX2_X1 U27248 ( .A(_02501__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR22) );
  MUX2_X1 U27249 ( .A(_02501__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR23) );
  MUX2_X1 U27250 ( .A(_02501__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR32) );
  MUX2_X1 U27251 ( .A(_02501__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR33) );
  MUX2_X1 U27252 ( .A(_02501__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR34) );
  MUX2_X1 U27253 ( .A(_02501__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR35) );
  MUX2_X1 U27254 ( .A(_02501__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR36) );
  MUX2_X1 U27255 ( .A(_02501__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR37) );
  MUX2_X1 U27256 ( .A(_02501__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR38) );
  MUX2_X1 U27257 ( .A(_02501__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR39) );
  MUX2_X1 U27258 ( .A(_02501__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR64) );
  MUX2_X1 U27259 ( .A(_02501__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR65) );
  MUX2_X1 U27260 ( .A(_02501__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR66) );
  MUX2_X1 U27261 ( .A(_02501__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR67) );
  MUX2_X1 U27262 ( .A(_02501__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR68) );
  MUX2_X1 U27263 ( .A(_02501__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR69) );
  MUX2_X1 U27264 ( .A(_02501__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR70) );
  MUX2_X1 U27265 ( .A(_02501__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03387__PTR71) );
  MUX2_X1 U27266 ( .A(_03392__PTR0), .B(_03390__PTR64), .S(P3_P1_State2_PTR3), .Z(_02504__PTR0) );
  MUX2_X1 U27267 ( .A(_03392__PTR1), .B(_03390__PTR65), .S(P3_P1_State2_PTR3), .Z(_02504__PTR1) );
  MUX2_X1 U27268 ( .A(_03392__PTR2), .B(_03390__PTR66), .S(P3_P1_State2_PTR3), .Z(_02504__PTR2) );
  MUX2_X1 U27269 ( .A(_03392__PTR3), .B(_03390__PTR67), .S(P3_P1_State2_PTR3), .Z(_02504__PTR3) );
  MUX2_X1 U27270 ( .A(_03392__PTR4), .B(_03390__PTR68), .S(P3_P1_State2_PTR3), .Z(_02504__PTR4) );
  MUX2_X1 U27271 ( .A(_03392__PTR5), .B(_03390__PTR69), .S(P3_P1_State2_PTR3), .Z(_02504__PTR5) );
  MUX2_X1 U27272 ( .A(_03392__PTR6), .B(_03390__PTR70), .S(P3_P1_State2_PTR3), .Z(_02504__PTR6) );
  MUX2_X1 U27273 ( .A(_03392__PTR7), .B(_03390__PTR71), .S(P3_P1_State2_PTR3), .Z(_02504__PTR7) );
  MUX2_X1 U27274 ( .A(_03391__PTR0), .B(_03391__PTR32), .S(P3_P1_State2_PTR2), .Z(_03392__PTR0) );
  MUX2_X1 U27275 ( .A(_03391__PTR1), .B(_03391__PTR33), .S(P3_P1_State2_PTR2), .Z(_03392__PTR1) );
  MUX2_X1 U27276 ( .A(_03391__PTR2), .B(_03391__PTR34), .S(P3_P1_State2_PTR2), .Z(_03392__PTR2) );
  MUX2_X1 U27277 ( .A(_03391__PTR3), .B(_03391__PTR35), .S(P3_P1_State2_PTR2), .Z(_03392__PTR3) );
  MUX2_X1 U27278 ( .A(_03391__PTR4), .B(_03391__PTR36), .S(P3_P1_State2_PTR2), .Z(_03392__PTR4) );
  MUX2_X1 U27279 ( .A(_03391__PTR5), .B(_03391__PTR37), .S(P3_P1_State2_PTR2), .Z(_03392__PTR5) );
  MUX2_X1 U27280 ( .A(_03391__PTR6), .B(_03391__PTR38), .S(P3_P1_State2_PTR2), .Z(_03392__PTR6) );
  MUX2_X1 U27281 ( .A(_03391__PTR7), .B(_03391__PTR39), .S(P3_P1_State2_PTR2), .Z(_03392__PTR7) );
  MUX2_X1 U27282 ( .A(1'b0), .B(_03390__PTR16), .S(P3_P1_State2_PTR1), .Z(_03391__PTR0) );
  MUX2_X1 U27283 ( .A(1'b0), .B(_03390__PTR17), .S(P3_P1_State2_PTR1), .Z(_03391__PTR1) );
  MUX2_X1 U27284 ( .A(1'b0), .B(_03390__PTR18), .S(P3_P1_State2_PTR1), .Z(_03391__PTR2) );
  MUX2_X1 U27285 ( .A(1'b0), .B(_03390__PTR19), .S(P3_P1_State2_PTR1), .Z(_03391__PTR3) );
  MUX2_X1 U27286 ( .A(1'b0), .B(_03390__PTR20), .S(P3_P1_State2_PTR1), .Z(_03391__PTR4) );
  MUX2_X1 U27287 ( .A(1'b0), .B(_03390__PTR21), .S(P3_P1_State2_PTR1), .Z(_03391__PTR5) );
  MUX2_X1 U27288 ( .A(1'b0), .B(_03390__PTR22), .S(P3_P1_State2_PTR1), .Z(_03391__PTR6) );
  MUX2_X1 U27289 ( .A(1'b0), .B(_03390__PTR23), .S(P3_P1_State2_PTR1), .Z(_03391__PTR7) );
  MUX2_X1 U27290 ( .A(_03390__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03391__PTR32) );
  MUX2_X1 U27291 ( .A(_03390__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03391__PTR33) );
  MUX2_X1 U27292 ( .A(_03390__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03391__PTR34) );
  MUX2_X1 U27293 ( .A(_03390__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03391__PTR35) );
  MUX2_X1 U27294 ( .A(_03390__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03391__PTR36) );
  MUX2_X1 U27295 ( .A(_03390__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03391__PTR37) );
  MUX2_X1 U27296 ( .A(_03390__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03391__PTR38) );
  MUX2_X1 U27297 ( .A(_03390__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03391__PTR39) );
  MUX2_X1 U27298 ( .A(_02503__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR16) );
  MUX2_X1 U27299 ( .A(_02503__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR17) );
  MUX2_X1 U27300 ( .A(_02503__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR18) );
  MUX2_X1 U27301 ( .A(_02503__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR19) );
  MUX2_X1 U27302 ( .A(_02503__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR20) );
  MUX2_X1 U27303 ( .A(_02503__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR21) );
  MUX2_X1 U27304 ( .A(_02503__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR22) );
  MUX2_X1 U27305 ( .A(_02503__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR23) );
  MUX2_X1 U27306 ( .A(_02503__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR32) );
  MUX2_X1 U27307 ( .A(_02503__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR33) );
  MUX2_X1 U27308 ( .A(_02503__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR34) );
  MUX2_X1 U27309 ( .A(_02503__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR35) );
  MUX2_X1 U27310 ( .A(_02503__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR36) );
  MUX2_X1 U27311 ( .A(_02503__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR37) );
  MUX2_X1 U27312 ( .A(_02503__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR38) );
  MUX2_X1 U27313 ( .A(_02503__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR39) );
  MUX2_X1 U27314 ( .A(_02503__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR64) );
  MUX2_X1 U27315 ( .A(_02503__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR65) );
  MUX2_X1 U27316 ( .A(_02503__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR66) );
  MUX2_X1 U27317 ( .A(_02503__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR67) );
  MUX2_X1 U27318 ( .A(_02503__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR68) );
  MUX2_X1 U27319 ( .A(_02503__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR69) );
  MUX2_X1 U27320 ( .A(_02503__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR70) );
  MUX2_X1 U27321 ( .A(_02503__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03390__PTR71) );
  MUX2_X1 U27322 ( .A(_03395__PTR0), .B(_03393__PTR64), .S(P3_P1_State2_PTR3), .Z(_02506__PTR0) );
  MUX2_X1 U27323 ( .A(_03395__PTR1), .B(_03393__PTR65), .S(P3_P1_State2_PTR3), .Z(_02506__PTR1) );
  MUX2_X1 U27324 ( .A(_03395__PTR2), .B(_03393__PTR66), .S(P3_P1_State2_PTR3), .Z(_02506__PTR2) );
  MUX2_X1 U27325 ( .A(_03395__PTR3), .B(_03393__PTR67), .S(P3_P1_State2_PTR3), .Z(_02506__PTR3) );
  MUX2_X1 U27326 ( .A(_03395__PTR4), .B(_03393__PTR68), .S(P3_P1_State2_PTR3), .Z(_02506__PTR4) );
  MUX2_X1 U27327 ( .A(_03395__PTR5), .B(_03393__PTR69), .S(P3_P1_State2_PTR3), .Z(_02506__PTR5) );
  MUX2_X1 U27328 ( .A(_03395__PTR6), .B(_03393__PTR70), .S(P3_P1_State2_PTR3), .Z(_02506__PTR6) );
  MUX2_X1 U27329 ( .A(_03395__PTR7), .B(_03393__PTR71), .S(P3_P1_State2_PTR3), .Z(_02506__PTR7) );
  MUX2_X1 U27330 ( .A(_03394__PTR0), .B(_03394__PTR32), .S(P3_P1_State2_PTR2), .Z(_03395__PTR0) );
  MUX2_X1 U27331 ( .A(_03394__PTR1), .B(_03394__PTR33), .S(P3_P1_State2_PTR2), .Z(_03395__PTR1) );
  MUX2_X1 U27332 ( .A(_03394__PTR2), .B(_03394__PTR34), .S(P3_P1_State2_PTR2), .Z(_03395__PTR2) );
  MUX2_X1 U27333 ( .A(_03394__PTR3), .B(_03394__PTR35), .S(P3_P1_State2_PTR2), .Z(_03395__PTR3) );
  MUX2_X1 U27334 ( .A(_03394__PTR4), .B(_03394__PTR36), .S(P3_P1_State2_PTR2), .Z(_03395__PTR4) );
  MUX2_X1 U27335 ( .A(_03394__PTR5), .B(_03394__PTR37), .S(P3_P1_State2_PTR2), .Z(_03395__PTR5) );
  MUX2_X1 U27336 ( .A(_03394__PTR6), .B(_03394__PTR38), .S(P3_P1_State2_PTR2), .Z(_03395__PTR6) );
  MUX2_X1 U27337 ( .A(_03394__PTR7), .B(_03394__PTR39), .S(P3_P1_State2_PTR2), .Z(_03395__PTR7) );
  MUX2_X1 U27338 ( .A(1'b0), .B(_03393__PTR16), .S(P3_P1_State2_PTR1), .Z(_03394__PTR0) );
  MUX2_X1 U27339 ( .A(1'b0), .B(_03393__PTR17), .S(P3_P1_State2_PTR1), .Z(_03394__PTR1) );
  MUX2_X1 U27340 ( .A(1'b0), .B(_03393__PTR18), .S(P3_P1_State2_PTR1), .Z(_03394__PTR2) );
  MUX2_X1 U27341 ( .A(1'b0), .B(_03393__PTR19), .S(P3_P1_State2_PTR1), .Z(_03394__PTR3) );
  MUX2_X1 U27342 ( .A(1'b0), .B(_03393__PTR20), .S(P3_P1_State2_PTR1), .Z(_03394__PTR4) );
  MUX2_X1 U27343 ( .A(1'b0), .B(_03393__PTR21), .S(P3_P1_State2_PTR1), .Z(_03394__PTR5) );
  MUX2_X1 U27344 ( .A(1'b0), .B(_03393__PTR22), .S(P3_P1_State2_PTR1), .Z(_03394__PTR6) );
  MUX2_X1 U27345 ( .A(1'b0), .B(_03393__PTR23), .S(P3_P1_State2_PTR1), .Z(_03394__PTR7) );
  MUX2_X1 U27346 ( .A(_03393__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03394__PTR32) );
  MUX2_X1 U27347 ( .A(_03393__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03394__PTR33) );
  MUX2_X1 U27348 ( .A(_03393__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03394__PTR34) );
  MUX2_X1 U27349 ( .A(_03393__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03394__PTR35) );
  MUX2_X1 U27350 ( .A(_03393__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03394__PTR36) );
  MUX2_X1 U27351 ( .A(_03393__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03394__PTR37) );
  MUX2_X1 U27352 ( .A(_03393__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03394__PTR38) );
  MUX2_X1 U27353 ( .A(_03393__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03394__PTR39) );
  MUX2_X1 U27354 ( .A(_02505__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR16) );
  MUX2_X1 U27355 ( .A(_02505__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR17) );
  MUX2_X1 U27356 ( .A(_02505__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR18) );
  MUX2_X1 U27357 ( .A(_02505__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR19) );
  MUX2_X1 U27358 ( .A(_02505__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR20) );
  MUX2_X1 U27359 ( .A(_02505__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR21) );
  MUX2_X1 U27360 ( .A(_02505__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR22) );
  MUX2_X1 U27361 ( .A(_02505__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR23) );
  MUX2_X1 U27362 ( .A(_02505__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR32) );
  MUX2_X1 U27363 ( .A(_02505__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR33) );
  MUX2_X1 U27364 ( .A(_02505__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR34) );
  MUX2_X1 U27365 ( .A(_02505__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR35) );
  MUX2_X1 U27366 ( .A(_02505__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR36) );
  MUX2_X1 U27367 ( .A(_02505__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR37) );
  MUX2_X1 U27368 ( .A(_02505__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR38) );
  MUX2_X1 U27369 ( .A(_02505__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR39) );
  MUX2_X1 U27370 ( .A(_02505__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR64) );
  MUX2_X1 U27371 ( .A(_02505__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR65) );
  MUX2_X1 U27372 ( .A(_02505__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR66) );
  MUX2_X1 U27373 ( .A(_02505__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR67) );
  MUX2_X1 U27374 ( .A(_02505__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR68) );
  MUX2_X1 U27375 ( .A(_02505__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR69) );
  MUX2_X1 U27376 ( .A(_02505__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR70) );
  MUX2_X1 U27377 ( .A(_02505__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03393__PTR71) );
  MUX2_X1 U27378 ( .A(_03398__PTR0), .B(_03396__PTR64), .S(P3_P1_State2_PTR3), .Z(_02508__PTR0) );
  MUX2_X1 U27379 ( .A(_03398__PTR1), .B(_03396__PTR65), .S(P3_P1_State2_PTR3), .Z(_02508__PTR1) );
  MUX2_X1 U27380 ( .A(_03398__PTR2), .B(_03396__PTR66), .S(P3_P1_State2_PTR3), .Z(_02508__PTR2) );
  MUX2_X1 U27381 ( .A(_03398__PTR3), .B(_03396__PTR67), .S(P3_P1_State2_PTR3), .Z(_02508__PTR3) );
  MUX2_X1 U27382 ( .A(_03398__PTR4), .B(_03396__PTR68), .S(P3_P1_State2_PTR3), .Z(_02508__PTR4) );
  MUX2_X1 U27383 ( .A(_03398__PTR5), .B(_03396__PTR69), .S(P3_P1_State2_PTR3), .Z(_02508__PTR5) );
  MUX2_X1 U27384 ( .A(_03398__PTR6), .B(_03396__PTR70), .S(P3_P1_State2_PTR3), .Z(_02508__PTR6) );
  MUX2_X1 U27385 ( .A(_03398__PTR7), .B(_03396__PTR71), .S(P3_P1_State2_PTR3), .Z(_02508__PTR7) );
  MUX2_X1 U27386 ( .A(_03397__PTR0), .B(_03397__PTR32), .S(P3_P1_State2_PTR2), .Z(_03398__PTR0) );
  MUX2_X1 U27387 ( .A(_03397__PTR1), .B(_03397__PTR33), .S(P3_P1_State2_PTR2), .Z(_03398__PTR1) );
  MUX2_X1 U27388 ( .A(_03397__PTR2), .B(_03397__PTR34), .S(P3_P1_State2_PTR2), .Z(_03398__PTR2) );
  MUX2_X1 U27389 ( .A(_03397__PTR3), .B(_03397__PTR35), .S(P3_P1_State2_PTR2), .Z(_03398__PTR3) );
  MUX2_X1 U27390 ( .A(_03397__PTR4), .B(_03397__PTR36), .S(P3_P1_State2_PTR2), .Z(_03398__PTR4) );
  MUX2_X1 U27391 ( .A(_03397__PTR5), .B(_03397__PTR37), .S(P3_P1_State2_PTR2), .Z(_03398__PTR5) );
  MUX2_X1 U27392 ( .A(_03397__PTR6), .B(_03397__PTR38), .S(P3_P1_State2_PTR2), .Z(_03398__PTR6) );
  MUX2_X1 U27393 ( .A(_03397__PTR7), .B(_03397__PTR39), .S(P3_P1_State2_PTR2), .Z(_03398__PTR7) );
  MUX2_X1 U27394 ( .A(1'b0), .B(_03396__PTR16), .S(P3_P1_State2_PTR1), .Z(_03397__PTR0) );
  MUX2_X1 U27395 ( .A(1'b0), .B(_03396__PTR17), .S(P3_P1_State2_PTR1), .Z(_03397__PTR1) );
  MUX2_X1 U27396 ( .A(1'b0), .B(_03396__PTR18), .S(P3_P1_State2_PTR1), .Z(_03397__PTR2) );
  MUX2_X1 U27397 ( .A(1'b0), .B(_03396__PTR19), .S(P3_P1_State2_PTR1), .Z(_03397__PTR3) );
  MUX2_X1 U27398 ( .A(1'b0), .B(_03396__PTR20), .S(P3_P1_State2_PTR1), .Z(_03397__PTR4) );
  MUX2_X1 U27399 ( .A(1'b0), .B(_03396__PTR21), .S(P3_P1_State2_PTR1), .Z(_03397__PTR5) );
  MUX2_X1 U27400 ( .A(1'b0), .B(_03396__PTR22), .S(P3_P1_State2_PTR1), .Z(_03397__PTR6) );
  MUX2_X1 U27401 ( .A(1'b0), .B(_03396__PTR23), .S(P3_P1_State2_PTR1), .Z(_03397__PTR7) );
  MUX2_X1 U27402 ( .A(_03396__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03397__PTR32) );
  MUX2_X1 U27403 ( .A(_03396__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03397__PTR33) );
  MUX2_X1 U27404 ( .A(_03396__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03397__PTR34) );
  MUX2_X1 U27405 ( .A(_03396__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03397__PTR35) );
  MUX2_X1 U27406 ( .A(_03396__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03397__PTR36) );
  MUX2_X1 U27407 ( .A(_03396__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03397__PTR37) );
  MUX2_X1 U27408 ( .A(_03396__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03397__PTR38) );
  MUX2_X1 U27409 ( .A(_03396__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03397__PTR39) );
  MUX2_X1 U27410 ( .A(_02507__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR16) );
  MUX2_X1 U27411 ( .A(_02507__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR17) );
  MUX2_X1 U27412 ( .A(_02507__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR18) );
  MUX2_X1 U27413 ( .A(_02507__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR19) );
  MUX2_X1 U27414 ( .A(_02507__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR20) );
  MUX2_X1 U27415 ( .A(_02507__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR21) );
  MUX2_X1 U27416 ( .A(_02507__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR22) );
  MUX2_X1 U27417 ( .A(_02507__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR23) );
  MUX2_X1 U27418 ( .A(_02507__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR32) );
  MUX2_X1 U27419 ( .A(_02507__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR33) );
  MUX2_X1 U27420 ( .A(_02507__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR34) );
  MUX2_X1 U27421 ( .A(_02507__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR35) );
  MUX2_X1 U27422 ( .A(_02507__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR36) );
  MUX2_X1 U27423 ( .A(_02507__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR37) );
  MUX2_X1 U27424 ( .A(_02507__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR38) );
  MUX2_X1 U27425 ( .A(_02507__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR39) );
  MUX2_X1 U27426 ( .A(_02507__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR64) );
  MUX2_X1 U27427 ( .A(_02507__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR65) );
  MUX2_X1 U27428 ( .A(_02507__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR66) );
  MUX2_X1 U27429 ( .A(_02507__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR67) );
  MUX2_X1 U27430 ( .A(_02507__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR68) );
  MUX2_X1 U27431 ( .A(_02507__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR69) );
  MUX2_X1 U27432 ( .A(_02507__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR70) );
  MUX2_X1 U27433 ( .A(_02507__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03396__PTR71) );
  MUX2_X1 U27434 ( .A(_03401__PTR0), .B(_03399__PTR64), .S(P3_P1_State2_PTR3), .Z(_02510__PTR0) );
  MUX2_X1 U27435 ( .A(_03401__PTR1), .B(_03399__PTR65), .S(P3_P1_State2_PTR3), .Z(_02510__PTR1) );
  MUX2_X1 U27436 ( .A(_03401__PTR2), .B(_03399__PTR66), .S(P3_P1_State2_PTR3), .Z(_02510__PTR2) );
  MUX2_X1 U27437 ( .A(_03401__PTR3), .B(_03399__PTR67), .S(P3_P1_State2_PTR3), .Z(_02510__PTR3) );
  MUX2_X1 U27438 ( .A(_03401__PTR4), .B(_03399__PTR68), .S(P3_P1_State2_PTR3), .Z(_02510__PTR4) );
  MUX2_X1 U27439 ( .A(_03401__PTR5), .B(_03399__PTR69), .S(P3_P1_State2_PTR3), .Z(_02510__PTR5) );
  MUX2_X1 U27440 ( .A(_03401__PTR6), .B(_03399__PTR70), .S(P3_P1_State2_PTR3), .Z(_02510__PTR6) );
  MUX2_X1 U27441 ( .A(_03401__PTR7), .B(_03399__PTR71), .S(P3_P1_State2_PTR3), .Z(_02510__PTR7) );
  MUX2_X1 U27442 ( .A(_03400__PTR0), .B(_03400__PTR32), .S(P3_P1_State2_PTR2), .Z(_03401__PTR0) );
  MUX2_X1 U27443 ( .A(_03400__PTR1), .B(_03400__PTR33), .S(P3_P1_State2_PTR2), .Z(_03401__PTR1) );
  MUX2_X1 U27444 ( .A(_03400__PTR2), .B(_03400__PTR34), .S(P3_P1_State2_PTR2), .Z(_03401__PTR2) );
  MUX2_X1 U27445 ( .A(_03400__PTR3), .B(_03400__PTR35), .S(P3_P1_State2_PTR2), .Z(_03401__PTR3) );
  MUX2_X1 U27446 ( .A(_03400__PTR4), .B(_03400__PTR36), .S(P3_P1_State2_PTR2), .Z(_03401__PTR4) );
  MUX2_X1 U27447 ( .A(_03400__PTR5), .B(_03400__PTR37), .S(P3_P1_State2_PTR2), .Z(_03401__PTR5) );
  MUX2_X1 U27448 ( .A(_03400__PTR6), .B(_03400__PTR38), .S(P3_P1_State2_PTR2), .Z(_03401__PTR6) );
  MUX2_X1 U27449 ( .A(_03400__PTR7), .B(_03400__PTR39), .S(P3_P1_State2_PTR2), .Z(_03401__PTR7) );
  MUX2_X1 U27450 ( .A(1'b0), .B(_03399__PTR16), .S(P3_P1_State2_PTR1), .Z(_03400__PTR0) );
  MUX2_X1 U27451 ( .A(1'b0), .B(_03399__PTR17), .S(P3_P1_State2_PTR1), .Z(_03400__PTR1) );
  MUX2_X1 U27452 ( .A(1'b0), .B(_03399__PTR18), .S(P3_P1_State2_PTR1), .Z(_03400__PTR2) );
  MUX2_X1 U27453 ( .A(1'b0), .B(_03399__PTR19), .S(P3_P1_State2_PTR1), .Z(_03400__PTR3) );
  MUX2_X1 U27454 ( .A(1'b0), .B(_03399__PTR20), .S(P3_P1_State2_PTR1), .Z(_03400__PTR4) );
  MUX2_X1 U27455 ( .A(1'b0), .B(_03399__PTR21), .S(P3_P1_State2_PTR1), .Z(_03400__PTR5) );
  MUX2_X1 U27456 ( .A(1'b0), .B(_03399__PTR22), .S(P3_P1_State2_PTR1), .Z(_03400__PTR6) );
  MUX2_X1 U27457 ( .A(1'b0), .B(_03399__PTR23), .S(P3_P1_State2_PTR1), .Z(_03400__PTR7) );
  MUX2_X1 U27458 ( .A(_03399__PTR32), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03400__PTR32) );
  MUX2_X1 U27459 ( .A(_03399__PTR33), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03400__PTR33) );
  MUX2_X1 U27460 ( .A(_03399__PTR34), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03400__PTR34) );
  MUX2_X1 U27461 ( .A(_03399__PTR35), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03400__PTR35) );
  MUX2_X1 U27462 ( .A(_03399__PTR36), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03400__PTR36) );
  MUX2_X1 U27463 ( .A(_03399__PTR37), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03400__PTR37) );
  MUX2_X1 U27464 ( .A(_03399__PTR38), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03400__PTR38) );
  MUX2_X1 U27465 ( .A(_03399__PTR39), .B(1'b0), .S(P3_P1_State2_PTR1), .Z(_03400__PTR39) );
  MUX2_X1 U27466 ( .A(_02509__PTR16), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR16) );
  MUX2_X1 U27467 ( .A(_02509__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR17) );
  MUX2_X1 U27468 ( .A(_02509__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR18) );
  MUX2_X1 U27469 ( .A(_02509__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR19) );
  MUX2_X1 U27470 ( .A(_02509__PTR20), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR20) );
  MUX2_X1 U27471 ( .A(_02509__PTR21), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR21) );
  MUX2_X1 U27472 ( .A(_02509__PTR22), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR22) );
  MUX2_X1 U27473 ( .A(_02509__PTR23), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR23) );
  MUX2_X1 U27474 ( .A(_02509__PTR32), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR32) );
  MUX2_X1 U27475 ( .A(_02509__PTR33), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR33) );
  MUX2_X1 U27476 ( .A(_02509__PTR34), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR34) );
  MUX2_X1 U27477 ( .A(_02509__PTR35), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR35) );
  MUX2_X1 U27478 ( .A(_02509__PTR36), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR36) );
  MUX2_X1 U27479 ( .A(_02509__PTR37), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR37) );
  MUX2_X1 U27480 ( .A(_02509__PTR38), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR38) );
  MUX2_X1 U27481 ( .A(_02509__PTR39), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR39) );
  MUX2_X1 U27482 ( .A(_02509__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR64) );
  MUX2_X1 U27483 ( .A(_02509__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR65) );
  MUX2_X1 U27484 ( .A(_02509__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR66) );
  MUX2_X1 U27485 ( .A(_02509__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR67) );
  MUX2_X1 U27486 ( .A(_02509__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR68) );
  MUX2_X1 U27487 ( .A(_02509__PTR69), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR69) );
  MUX2_X1 U27488 ( .A(_02509__PTR70), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR70) );
  MUX2_X1 U27489 ( .A(_02509__PTR71), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03399__PTR71) );
  MUX2_X1 U27490 ( .A(_03404__PTR0), .B(_03402__PTR64), .S(P3_P1_State2_PTR3), .Z(_02512__PTR0) );
  MUX2_X1 U27491 ( .A(_03404__PTR1), .B(_03402__PTR65), .S(P3_P1_State2_PTR3), .Z(_02512__PTR1) );
  MUX2_X1 U27492 ( .A(_03404__PTR2), .B(_03402__PTR66), .S(P3_P1_State2_PTR3), .Z(_02512__PTR2) );
  MUX2_X1 U27493 ( .A(_03404__PTR3), .B(_03402__PTR67), .S(P3_P1_State2_PTR3), .Z(_02512__PTR3) );
  MUX2_X1 U27494 ( .A(_03404__PTR4), .B(_03402__PTR68), .S(P3_P1_State2_PTR3), .Z(_02512__PTR4) );
  MUX2_X1 U27495 ( .A(1'b0), .B(_03403__PTR32), .S(P3_P1_State2_PTR2), .Z(_03404__PTR0) );
  MUX2_X1 U27496 ( .A(_03403__PTR1), .B(_03403__PTR33), .S(P3_P1_State2_PTR2), .Z(_03404__PTR1) );
  MUX2_X1 U27497 ( .A(_03403__PTR2), .B(_03403__PTR34), .S(P3_P1_State2_PTR2), .Z(_03404__PTR2) );
  MUX2_X1 U27498 ( .A(_03403__PTR3), .B(_03403__PTR35), .S(P3_P1_State2_PTR2), .Z(_03404__PTR3) );
  MUX2_X1 U27499 ( .A(_03403__PTR4), .B(_03403__PTR36), .S(P3_P1_State2_PTR2), .Z(_03404__PTR4) );
  MUX2_X1 U27500 ( .A(1'b0), .B(_03402__PTR17), .S(P3_P1_State2_PTR1), .Z(_03403__PTR1) );
  MUX2_X1 U27501 ( .A(1'b0), .B(_03402__PTR18), .S(P3_P1_State2_PTR1), .Z(_03403__PTR2) );
  MUX2_X1 U27502 ( .A(1'b0), .B(_03402__PTR19), .S(P3_P1_State2_PTR1), .Z(_03403__PTR3) );
  MUX2_X1 U27503 ( .A(1'b0), .B(_03402__PTR36), .S(P3_P1_State2_PTR1), .Z(_03403__PTR4) );
  MUX2_X1 U27504 ( .A(1'b0), .B(_03402__PTR48), .S(P3_P1_State2_PTR1), .Z(_03403__PTR32) );
  MUX2_X1 U27505 ( .A(_03402__PTR33), .B(_03402__PTR52), .S(P3_P1_State2_PTR1), .Z(_03403__PTR33) );
  MUX2_X1 U27506 ( .A(_03402__PTR34), .B(_03402__PTR52), .S(P3_P1_State2_PTR1), .Z(_03403__PTR34) );
  MUX2_X1 U27507 ( .A(_03402__PTR35), .B(_03402__PTR52), .S(P3_P1_State2_PTR1), .Z(_03403__PTR35) );
  MUX2_X1 U27508 ( .A(_03402__PTR36), .B(_03402__PTR52), .S(P3_P1_State2_PTR1), .Z(_03403__PTR36) );
  MUX2_X1 U27509 ( .A(_02511__PTR17), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03402__PTR17) );
  MUX2_X1 U27510 ( .A(_02511__PTR18), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03402__PTR18) );
  MUX2_X1 U27511 ( .A(_02511__PTR19), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03402__PTR19) );
  MUX2_X1 U27512 ( .A(_02420__PTR1), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03402__PTR33) );
  MUX2_X1 U27513 ( .A(_02420__PTR2), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03402__PTR34) );
  MUX2_X1 U27514 ( .A(_02420__PTR3), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03402__PTR35) );
  MUX2_X1 U27515 ( .A(1'b0), .B(P3_P1_InstQueueWr_Addr_PTR4), .S(P3_P1_State2_PTR0), .Z(_03402__PTR36) );
  MUX2_X1 U27516 ( .A(1'b0), .B(_02511__PTR56), .S(P3_P1_State2_PTR0), .Z(_03402__PTR48) );
  MUX2_X1 U27517 ( .A(1'b0), .B(_02511__PTR60), .S(P3_P1_State2_PTR0), .Z(_03402__PTR52) );
  MUX2_X1 U27518 ( .A(_02511__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03402__PTR64) );
  MUX2_X1 U27519 ( .A(_02511__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03402__PTR65) );
  MUX2_X1 U27520 ( .A(_02511__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03402__PTR66) );
  MUX2_X1 U27521 ( .A(_02511__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03402__PTR67) );
  MUX2_X1 U27522 ( .A(_02511__PTR68), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03402__PTR68) );
  MUX2_X1 U27523 ( .A(_03407__PTR0), .B(_03405__PTR64), .S(P3_P1_State2_PTR3), .Z(_02514__PTR0) );
  MUX2_X1 U27524 ( .A(_03407__PTR1), .B(_03405__PTR65), .S(P3_P1_State2_PTR3), .Z(_02514__PTR1) );
  MUX2_X1 U27525 ( .A(_03407__PTR2), .B(_03405__PTR66), .S(P3_P1_State2_PTR3), .Z(_02514__PTR2) );
  MUX2_X1 U27526 ( .A(_03407__PTR3), .B(_03405__PTR67), .S(P3_P1_State2_PTR3), .Z(_02514__PTR3) );
  MUX2_X1 U27527 ( .A(_03407__PTR4), .B(_03351__PTR32), .S(P3_P1_State2_PTR3), .Z(_02514__PTR4) );
  MUX2_X1 U27528 ( .A(1'b0), .B(_03406__PTR32), .S(P3_P1_State2_PTR2), .Z(_03407__PTR0) );
  MUX2_X1 U27529 ( .A(1'b0), .B(_03406__PTR33), .S(P3_P1_State2_PTR2), .Z(_03407__PTR1) );
  MUX2_X1 U27530 ( .A(1'b0), .B(_03406__PTR34), .S(P3_P1_State2_PTR2), .Z(_03407__PTR2) );
  MUX2_X1 U27531 ( .A(1'b0), .B(_03406__PTR35), .S(P3_P1_State2_PTR2), .Z(_03407__PTR3) );
  MUX2_X1 U27532 ( .A(1'b0), .B(_03406__PTR36), .S(P3_P1_State2_PTR2), .Z(_03407__PTR4) );
  MUX2_X1 U27533 ( .A(_03405__PTR32), .B(_03405__PTR48), .S(P3_P1_State2_PTR1), .Z(_03406__PTR32) );
  MUX2_X1 U27534 ( .A(_03405__PTR33), .B(_03405__PTR49), .S(P3_P1_State2_PTR1), .Z(_03406__PTR33) );
  MUX2_X1 U27535 ( .A(_03405__PTR34), .B(_03405__PTR50), .S(P3_P1_State2_PTR1), .Z(_03406__PTR34) );
  MUX2_X1 U27536 ( .A(_03405__PTR35), .B(_03405__PTR51), .S(P3_P1_State2_PTR1), .Z(_03406__PTR35) );
  MUX2_X1 U27537 ( .A(_03405__PTR36), .B(_03405__PTR52), .S(P3_P1_State2_PTR1), .Z(_03406__PTR36) );
  MUX2_X1 U27538 ( .A(1'b0), .B(_02513__PTR40), .S(P3_P1_State2_PTR0), .Z(_03405__PTR32) );
  MUX2_X1 U27539 ( .A(1'b0), .B(_02513__PTR41), .S(P3_P1_State2_PTR0), .Z(_03405__PTR33) );
  MUX2_X1 U27540 ( .A(1'b0), .B(_02513__PTR42), .S(P3_P1_State2_PTR0), .Z(_03405__PTR34) );
  MUX2_X1 U27541 ( .A(1'b0), .B(_02513__PTR43), .S(P3_P1_State2_PTR0), .Z(_03405__PTR35) );
  MUX2_X1 U27542 ( .A(1'b0), .B(_02513__PTR44), .S(P3_P1_State2_PTR0), .Z(_03405__PTR36) );
  MUX2_X1 U27543 ( .A(1'b0), .B(_02513__PTR56), .S(P3_P1_State2_PTR0), .Z(_03405__PTR48) );
  MUX2_X1 U27544 ( .A(1'b0), .B(_02513__PTR57), .S(P3_P1_State2_PTR0), .Z(_03405__PTR49) );
  MUX2_X1 U27545 ( .A(1'b0), .B(_02513__PTR58), .S(P3_P1_State2_PTR0), .Z(_03405__PTR50) );
  MUX2_X1 U27546 ( .A(1'b0), .B(_02513__PTR59), .S(P3_P1_State2_PTR0), .Z(_03405__PTR51) );
  MUX2_X1 U27547 ( .A(1'b0), .B(_02513__PTR60), .S(P3_P1_State2_PTR0), .Z(_03405__PTR52) );
  MUX2_X1 U27548 ( .A(_02513__PTR64), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03405__PTR64) );
  MUX2_X1 U27549 ( .A(_02513__PTR65), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03405__PTR65) );
  MUX2_X1 U27550 ( .A(_02513__PTR66), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03405__PTR66) );
  MUX2_X1 U27551 ( .A(_02513__PTR67), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03405__PTR67) );
  MUX2_X1 U27552 ( .A(_03408__PTR256), .B(_03408__PTR384), .S(P3_P1_State2_PTR1), .Z(_03409__PTR256) );
  MUX2_X1 U27553 ( .A(_03408__PTR257), .B(_03408__PTR385), .S(P3_P1_State2_PTR1), .Z(_03409__PTR257) );
  MUX2_X1 U27554 ( .A(_03408__PTR258), .B(_03408__PTR386), .S(P3_P1_State2_PTR1), .Z(_03409__PTR258) );
  MUX2_X1 U27555 ( .A(_03408__PTR259), .B(_03408__PTR387), .S(P3_P1_State2_PTR1), .Z(_03409__PTR259) );
  MUX2_X1 U27556 ( .A(_03408__PTR260), .B(_03408__PTR388), .S(P3_P1_State2_PTR1), .Z(_03409__PTR260) );
  MUX2_X1 U27557 ( .A(_03408__PTR261), .B(_03408__PTR389), .S(P3_P1_State2_PTR1), .Z(_03409__PTR261) );
  MUX2_X1 U27558 ( .A(_03408__PTR262), .B(_03408__PTR390), .S(P3_P1_State2_PTR1), .Z(_03409__PTR262) );
  MUX2_X1 U27559 ( .A(_03408__PTR263), .B(_03408__PTR391), .S(P3_P1_State2_PTR1), .Z(_03409__PTR263) );
  MUX2_X1 U27560 ( .A(_03408__PTR264), .B(_03408__PTR392), .S(P3_P1_State2_PTR1), .Z(_03409__PTR264) );
  MUX2_X1 U27561 ( .A(_03408__PTR265), .B(_03408__PTR393), .S(P3_P1_State2_PTR1), .Z(_03409__PTR265) );
  MUX2_X1 U27562 ( .A(_03408__PTR266), .B(_03408__PTR394), .S(P3_P1_State2_PTR1), .Z(_03409__PTR266) );
  MUX2_X1 U27563 ( .A(_03408__PTR267), .B(_03408__PTR395), .S(P3_P1_State2_PTR1), .Z(_03409__PTR267) );
  MUX2_X1 U27564 ( .A(_03408__PTR268), .B(_03408__PTR396), .S(P3_P1_State2_PTR1), .Z(_03409__PTR268) );
  MUX2_X1 U27565 ( .A(_03408__PTR269), .B(_03408__PTR397), .S(P3_P1_State2_PTR1), .Z(_03409__PTR269) );
  MUX2_X1 U27566 ( .A(_03408__PTR270), .B(_03408__PTR398), .S(P3_P1_State2_PTR1), .Z(_03409__PTR270) );
  MUX2_X1 U27567 ( .A(_03408__PTR271), .B(_03408__PTR399), .S(P3_P1_State2_PTR1), .Z(_03409__PTR271) );
  MUX2_X1 U27568 ( .A(_03408__PTR272), .B(_03408__PTR400), .S(P3_P1_State2_PTR1), .Z(_03409__PTR272) );
  MUX2_X1 U27569 ( .A(_03408__PTR273), .B(_03408__PTR401), .S(P3_P1_State2_PTR1), .Z(_03409__PTR273) );
  MUX2_X1 U27570 ( .A(_03408__PTR274), .B(_03408__PTR402), .S(P3_P1_State2_PTR1), .Z(_03409__PTR274) );
  MUX2_X1 U27571 ( .A(_03408__PTR275), .B(_03408__PTR403), .S(P3_P1_State2_PTR1), .Z(_03409__PTR275) );
  MUX2_X1 U27572 ( .A(_03408__PTR276), .B(_03408__PTR404), .S(P3_P1_State2_PTR1), .Z(_03409__PTR276) );
  MUX2_X1 U27573 ( .A(_03408__PTR277), .B(_03408__PTR405), .S(P3_P1_State2_PTR1), .Z(_03409__PTR277) );
  MUX2_X1 U27574 ( .A(_03408__PTR278), .B(_03408__PTR406), .S(P3_P1_State2_PTR1), .Z(_03409__PTR278) );
  MUX2_X1 U27575 ( .A(_03408__PTR279), .B(_03408__PTR407), .S(P3_P1_State2_PTR1), .Z(_03409__PTR279) );
  MUX2_X1 U27576 ( .A(_03408__PTR280), .B(_03408__PTR408), .S(P3_P1_State2_PTR1), .Z(_03409__PTR280) );
  MUX2_X1 U27577 ( .A(_03408__PTR281), .B(_03408__PTR409), .S(P3_P1_State2_PTR1), .Z(_03409__PTR281) );
  MUX2_X1 U27578 ( .A(_03408__PTR282), .B(_03408__PTR410), .S(P3_P1_State2_PTR1), .Z(_03409__PTR282) );
  MUX2_X1 U27579 ( .A(_03408__PTR283), .B(_03408__PTR411), .S(P3_P1_State2_PTR1), .Z(_03409__PTR283) );
  MUX2_X1 U27580 ( .A(_03408__PTR284), .B(_03408__PTR412), .S(P3_P1_State2_PTR1), .Z(_03409__PTR284) );
  MUX2_X1 U27581 ( .A(_03408__PTR285), .B(_03408__PTR413), .S(P3_P1_State2_PTR1), .Z(_03409__PTR285) );
  MUX2_X1 U27582 ( .A(_03408__PTR286), .B(_03408__PTR414), .S(P3_P1_State2_PTR1), .Z(_03409__PTR286) );
  MUX2_X1 U27583 ( .A(_03408__PTR288), .B(_03351__PTR32), .S(P3_P1_State2_PTR1), .Z(_03409__PTR288) );
  MUX2_X1 U27584 ( .A(1'b0), .B(_02519__PTR320), .S(P3_P1_State2_PTR0), .Z(_03408__PTR256) );
  MUX2_X1 U27585 ( .A(1'b0), .B(_02519__PTR321), .S(P3_P1_State2_PTR0), .Z(_03408__PTR257) );
  MUX2_X1 U27586 ( .A(1'b0), .B(_02519__PTR322), .S(P3_P1_State2_PTR0), .Z(_03408__PTR258) );
  MUX2_X1 U27587 ( .A(1'b0), .B(_02519__PTR323), .S(P3_P1_State2_PTR0), .Z(_03408__PTR259) );
  MUX2_X1 U27588 ( .A(1'b0), .B(_02519__PTR324), .S(P3_P1_State2_PTR0), .Z(_03408__PTR260) );
  MUX2_X1 U27589 ( .A(1'b0), .B(_02519__PTR325), .S(P3_P1_State2_PTR0), .Z(_03408__PTR261) );
  MUX2_X1 U27590 ( .A(1'b0), .B(_02519__PTR326), .S(P3_P1_State2_PTR0), .Z(_03408__PTR262) );
  MUX2_X1 U27591 ( .A(1'b0), .B(_02519__PTR327), .S(P3_P1_State2_PTR0), .Z(_03408__PTR263) );
  MUX2_X1 U27592 ( .A(1'b0), .B(_02519__PTR328), .S(P3_P1_State2_PTR0), .Z(_03408__PTR264) );
  MUX2_X1 U27593 ( .A(1'b0), .B(_02519__PTR329), .S(P3_P1_State2_PTR0), .Z(_03408__PTR265) );
  MUX2_X1 U27594 ( .A(1'b0), .B(_02519__PTR330), .S(P3_P1_State2_PTR0), .Z(_03408__PTR266) );
  MUX2_X1 U27595 ( .A(1'b0), .B(_02519__PTR331), .S(P3_P1_State2_PTR0), .Z(_03408__PTR267) );
  MUX2_X1 U27596 ( .A(1'b0), .B(_02519__PTR332), .S(P3_P1_State2_PTR0), .Z(_03408__PTR268) );
  MUX2_X1 U27597 ( .A(1'b0), .B(_02519__PTR333), .S(P3_P1_State2_PTR0), .Z(_03408__PTR269) );
  MUX2_X1 U27598 ( .A(1'b0), .B(_02519__PTR334), .S(P3_P1_State2_PTR0), .Z(_03408__PTR270) );
  MUX2_X1 U27599 ( .A(1'b0), .B(_02519__PTR335), .S(P3_P1_State2_PTR0), .Z(_03408__PTR271) );
  MUX2_X1 U27600 ( .A(1'b0), .B(_02519__PTR336), .S(P3_P1_State2_PTR0), .Z(_03408__PTR272) );
  MUX2_X1 U27601 ( .A(1'b0), .B(_02519__PTR337), .S(P3_P1_State2_PTR0), .Z(_03408__PTR273) );
  MUX2_X1 U27602 ( .A(1'b0), .B(_02519__PTR338), .S(P3_P1_State2_PTR0), .Z(_03408__PTR274) );
  MUX2_X1 U27603 ( .A(1'b0), .B(_02519__PTR339), .S(P3_P1_State2_PTR0), .Z(_03408__PTR275) );
  MUX2_X1 U27604 ( .A(1'b0), .B(_02519__PTR340), .S(P3_P1_State2_PTR0), .Z(_03408__PTR276) );
  MUX2_X1 U27605 ( .A(1'b0), .B(_02519__PTR341), .S(P3_P1_State2_PTR0), .Z(_03408__PTR277) );
  MUX2_X1 U27606 ( .A(1'b0), .B(_02519__PTR342), .S(P3_P1_State2_PTR0), .Z(_03408__PTR278) );
  MUX2_X1 U27607 ( .A(1'b0), .B(_02519__PTR343), .S(P3_P1_State2_PTR0), .Z(_03408__PTR279) );
  MUX2_X1 U27608 ( .A(1'b0), .B(_02519__PTR344), .S(P3_P1_State2_PTR0), .Z(_03408__PTR280) );
  MUX2_X1 U27609 ( .A(1'b0), .B(_02519__PTR345), .S(P3_P1_State2_PTR0), .Z(_03408__PTR281) );
  MUX2_X1 U27610 ( .A(1'b0), .B(_02519__PTR346), .S(P3_P1_State2_PTR0), .Z(_03408__PTR282) );
  MUX2_X1 U27611 ( .A(1'b0), .B(_02519__PTR347), .S(P3_P1_State2_PTR0), .Z(_03408__PTR283) );
  MUX2_X1 U27612 ( .A(1'b0), .B(_02519__PTR348), .S(P3_P1_State2_PTR0), .Z(_03408__PTR284) );
  MUX2_X1 U27613 ( .A(1'b0), .B(_02519__PTR349), .S(P3_P1_State2_PTR0), .Z(_03408__PTR285) );
  MUX2_X1 U27614 ( .A(1'b0), .B(_02519__PTR350), .S(P3_P1_State2_PTR0), .Z(_03408__PTR286) );
  MUX2_X1 U27615 ( .A(1'b0), .B(_02519__PTR352), .S(P3_P1_State2_PTR0), .Z(_03408__PTR288) );
  MUX2_X1 U27616 ( .A(P3_P1_lWord_PTR0), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR384) );
  MUX2_X1 U27617 ( .A(P3_P1_lWord_PTR1), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR385) );
  MUX2_X1 U27618 ( .A(P3_P1_lWord_PTR2), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR386) );
  MUX2_X1 U27619 ( .A(P3_P1_lWord_PTR3), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR387) );
  MUX2_X1 U27620 ( .A(P3_P1_lWord_PTR4), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR388) );
  MUX2_X1 U27621 ( .A(P3_P1_lWord_PTR5), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR389) );
  MUX2_X1 U27622 ( .A(P3_P1_lWord_PTR6), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR390) );
  MUX2_X1 U27623 ( .A(P3_P1_lWord_PTR7), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR391) );
  MUX2_X1 U27624 ( .A(P3_P1_lWord_PTR8), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR392) );
  MUX2_X1 U27625 ( .A(P3_P1_lWord_PTR9), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR393) );
  MUX2_X1 U27626 ( .A(P3_P1_lWord_PTR10), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR394) );
  MUX2_X1 U27627 ( .A(P3_P1_lWord_PTR11), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR395) );
  MUX2_X1 U27628 ( .A(P3_P1_lWord_PTR12), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR396) );
  MUX2_X1 U27629 ( .A(P3_P1_lWord_PTR13), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR397) );
  MUX2_X1 U27630 ( .A(P3_P1_lWord_PTR14), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR398) );
  MUX2_X1 U27631 ( .A(P3_P1_lWord_PTR15), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR399) );
  MUX2_X1 U27632 ( .A(P3_P1_uWord_PTR0), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR400) );
  MUX2_X1 U27633 ( .A(P3_P1_uWord_PTR1), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR401) );
  MUX2_X1 U27634 ( .A(P3_P1_uWord_PTR2), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR402) );
  MUX2_X1 U27635 ( .A(P3_P1_uWord_PTR3), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR403) );
  MUX2_X1 U27636 ( .A(P3_P1_uWord_PTR4), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR404) );
  MUX2_X1 U27637 ( .A(P3_P1_uWord_PTR5), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR405) );
  MUX2_X1 U27638 ( .A(P3_P1_uWord_PTR6), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR406) );
  MUX2_X1 U27639 ( .A(P3_P1_uWord_PTR7), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR407) );
  MUX2_X1 U27640 ( .A(P3_P1_uWord_PTR8), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR408) );
  MUX2_X1 U27641 ( .A(P3_P1_uWord_PTR9), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR409) );
  MUX2_X1 U27642 ( .A(P3_P1_uWord_PTR10), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR410) );
  MUX2_X1 U27643 ( .A(P3_P1_uWord_PTR11), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR411) );
  MUX2_X1 U27644 ( .A(P3_P1_uWord_PTR12), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR412) );
  MUX2_X1 U27645 ( .A(P3_P1_uWord_PTR13), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR413) );
  MUX2_X1 U27646 ( .A(P3_P1_uWord_PTR14), .B(1'b0), .S(P3_P1_State2_PTR0), .Z(_03408__PTR414) );
  BUF_X1 U27647 ( .A(_01855__PTR1), .Z(_00466__PTR1) );
  BUF_X1 U27648 ( .A(_00471__PTR1), .Z(_00472__PTR0) );
  BUF_X1 U27649 ( .A(_01870__PTR1), .Z(_00519__PTR1) );
  BUF_X1 U27650 ( .A(_00469__PTR1), .Z(_00584__PTR1) );
  BUF_X1 U27651 ( .A(_02719__PTR3), .Z(_00618__PTR1) );
  BUF_X1 U27652 ( .A(_00618__PTR2), .Z(_00620__PTR2) );
  BUF_X1 U27653 ( .A(_02412__PTR4), .Z(_00624__PTR0) );
  BUF_X1 U27654 ( .A(_02412__PTR5), .Z(_00625__PTR0) );
  BUF_X1 U27655 ( .A(_02412__PTR6), .Z(_00626__PTR0) );
  BUF_X1 U27656 ( .A(_02148__PTR1), .Z(_00790__PTR1) );
  BUF_X1 U27657 ( .A(_00803__PTR1), .Z(_00804__PTR0) );
  BUF_X1 U27658 ( .A(_02163__PTR1), .Z(_00843__PTR1) );
  BUF_X1 U27659 ( .A(_00793__PTR1), .Z(_00908__PTR1) );
  BUF_X1 U27660 ( .A(_02964__PTR3), .Z(_00942__PTR1) );
  BUF_X1 U27661 ( .A(_00942__PTR2), .Z(_00944__PTR2) );
  BUF_X1 U27662 ( .A(_02701__PTR4), .Z(_00948__PTR0) );
  BUF_X1 U27663 ( .A(_02701__PTR5), .Z(_00949__PTR0) );
  BUF_X1 U27664 ( .A(_02701__PTR6), .Z(_00950__PTR0) );
  BUF_X1 U27665 ( .A(_02437__PTR1), .Z(_01114__PTR1) );
  BUF_X1 U27666 ( .A(_01127__PTR1), .Z(_01128__PTR0) );
  BUF_X1 U27667 ( .A(_02452__PTR1), .Z(_01167__PTR1) );
  BUF_X1 U27668 ( .A(_01117__PTR1), .Z(_01232__PTR1) );
  BUF_X1 U27669 ( .A(_03209__PTR3), .Z(_01266__PTR1) );
  BUF_X1 U27670 ( .A(_01266__PTR2), .Z(_01268__PTR2) );
  BUF_X1 U27671 ( .A(_01277__PTR0), .Z(_01281__PTR0) );
  BUF_X1 U27672 ( .A(_01281__PTR1), .Z(_01285__PTR1) );
  BUF_X1 U27673 ( .A(_01283__PTR1), .Z(_01289__PTR1) );
  BUF_X1 U27674 ( .A(_01288__PTR1), .Z(_01291__PTR1) );
  BUF_X1 U27675 ( .A(_01283__PTR1), .Z(_01292__PTR1) );
  BUF_X1 U27676 ( .A(_01288__PTR1), .Z(_01294__PTR1) );
  BUF_X1 U27677 ( .A(_01283__PTR1), .Z(_01295__PTR1) );
  BUF_X1 U27678 ( .A(_01288__PTR1), .Z(_01297__PTR1) );
  BUF_X1 U27679 ( .A(_01283__PTR1), .Z(_01298__PTR1) );
  BUF_X1 U27680 ( .A(_01288__PTR1), .Z(_01300__PTR1) );
  BUF_X1 U27681 ( .A(_01283__PTR1), .Z(_01301__PTR1) );
  BUF_X1 U27682 ( .A(_01288__PTR1), .Z(_01303__PTR1) );
  BUF_X1 U27683 ( .A(_01283__PTR1), .Z(_01304__PTR1) );
  BUF_X1 U27684 ( .A(_01288__PTR1), .Z(_01306__PTR1) );
  BUF_X1 U27685 ( .A(_01283__PTR1), .Z(_01307__PTR1) );
  BUF_X1 U27686 ( .A(_01288__PTR1), .Z(_01309__PTR1) );
  BUF_X1 U27687 ( .A(_01283__PTR1), .Z(_01310__PTR1) );
  BUF_X1 U27688 ( .A(_01288__PTR1), .Z(_01312__PTR1) );
  BUF_X1 U27689 ( .A(_01283__PTR1), .Z(_01313__PTR1) );
  BUF_X1 U27690 ( .A(_01288__PTR1), .Z(_01315__PTR1) );
  BUF_X1 U27691 ( .A(_01283__PTR1), .Z(_01316__PTR1) );
  BUF_X1 U27692 ( .A(_01288__PTR1), .Z(_01318__PTR1) );
  BUF_X1 U27693 ( .A(_01283__PTR1), .Z(_01319__PTR1) );
  BUF_X1 U27694 ( .A(_01288__PTR1), .Z(_01321__PTR1) );
  BUF_X1 U27695 ( .A(_01283__PTR1), .Z(_01322__PTR1) );
  BUF_X1 U27696 ( .A(_01288__PTR1), .Z(_01324__PTR1) );
  BUF_X1 U27697 ( .A(_01283__PTR1), .Z(_01325__PTR1) );
  BUF_X1 U27698 ( .A(_01288__PTR1), .Z(_01327__PTR1) );
  BUF_X1 U27699 ( .A(_01283__PTR1), .Z(_01328__PTR1) );
  BUF_X1 U27700 ( .A(_01288__PTR1), .Z(_01330__PTR1) );
  BUF_X1 U27701 ( .A(_01283__PTR1), .Z(_01331__PTR1) );
  BUF_X1 U27702 ( .A(_01288__PTR1), .Z(_01333__PTR1) );
  BUF_X1 U27703 ( .A(_01339__PTR1), .Z(_01341__PTR1) );
  BUF_X1 U27704 ( .A(_01349__PTR0), .Z(_01353__PTR0) );
  BUF_X1 U27705 ( .A(_01353__PTR1), .Z(_01357__PTR1) );
  BUF_X1 U27706 ( .A(_01355__PTR1), .Z(_01361__PTR1) );
  BUF_X1 U27707 ( .A(_01360__PTR1), .Z(_01363__PTR1) );
  BUF_X1 U27708 ( .A(_01355__PTR1), .Z(_01364__PTR1) );
  BUF_X1 U27709 ( .A(_01360__PTR1), .Z(_01366__PTR1) );
  BUF_X1 U27710 ( .A(_01355__PTR1), .Z(_01367__PTR1) );
  BUF_X1 U27711 ( .A(_01360__PTR1), .Z(_01369__PTR1) );
  BUF_X1 U27712 ( .A(_01355__PTR1), .Z(_01370__PTR1) );
  BUF_X1 U27713 ( .A(_01360__PTR1), .Z(_01372__PTR1) );
  BUF_X1 U27714 ( .A(_01355__PTR1), .Z(_01373__PTR1) );
  BUF_X1 U27715 ( .A(_01360__PTR1), .Z(_01375__PTR1) );
  BUF_X1 U27716 ( .A(_01355__PTR1), .Z(_01376__PTR1) );
  BUF_X1 U27717 ( .A(_01360__PTR1), .Z(_01378__PTR1) );
  BUF_X1 U27718 ( .A(_01355__PTR1), .Z(_01379__PTR1) );
  BUF_X1 U27719 ( .A(_01360__PTR1), .Z(_01381__PTR1) );
  BUF_X1 U27720 ( .A(_01355__PTR1), .Z(_01382__PTR1) );
  BUF_X1 U27721 ( .A(_01360__PTR1), .Z(_01384__PTR1) );
  BUF_X1 U27722 ( .A(_01355__PTR1), .Z(_01385__PTR1) );
  BUF_X1 U27723 ( .A(_01360__PTR1), .Z(_01387__PTR1) );
  BUF_X1 U27724 ( .A(_01355__PTR1), .Z(_01388__PTR1) );
  BUF_X1 U27725 ( .A(_01360__PTR1), .Z(_01390__PTR1) );
  BUF_X1 U27726 ( .A(_01355__PTR1), .Z(_01391__PTR1) );
  BUF_X1 U27727 ( .A(_01360__PTR1), .Z(_01393__PTR1) );
  BUF_X1 U27728 ( .A(_01355__PTR1), .Z(_01394__PTR1) );
  BUF_X1 U27729 ( .A(_01360__PTR1), .Z(_01396__PTR1) );
  BUF_X1 U27730 ( .A(_01355__PTR1), .Z(_01397__PTR1) );
  BUF_X1 U27731 ( .A(_01360__PTR1), .Z(_01399__PTR1) );
  BUF_X1 U27732 ( .A(_01355__PTR1), .Z(_01400__PTR1) );
  BUF_X1 U27733 ( .A(_01360__PTR1), .Z(_01402__PTR1) );
  BUF_X1 U27734 ( .A(_01355__PTR1), .Z(_01403__PTR1) );
  BUF_X1 U27735 ( .A(_01360__PTR1), .Z(_01405__PTR1) );
  BUF_X1 U27736 ( .A(_01411__PTR1), .Z(_01413__PTR1) );
  BUF_X1 U27737 ( .A(_01421__PTR0), .Z(_01425__PTR0) );
  BUF_X1 U27738 ( .A(_01425__PTR1), .Z(_01429__PTR1) );
  BUF_X1 U27739 ( .A(_01427__PTR1), .Z(_01433__PTR1) );
  BUF_X1 U27740 ( .A(_01432__PTR1), .Z(_01435__PTR1) );
  BUF_X1 U27741 ( .A(_01427__PTR1), .Z(_01436__PTR1) );
  BUF_X1 U27742 ( .A(_01432__PTR1), .Z(_01438__PTR1) );
  BUF_X1 U27743 ( .A(_01427__PTR1), .Z(_01439__PTR1) );
  BUF_X1 U27744 ( .A(_01432__PTR1), .Z(_01441__PTR1) );
  BUF_X1 U27745 ( .A(_01427__PTR1), .Z(_01442__PTR1) );
  BUF_X1 U27746 ( .A(_01432__PTR1), .Z(_01444__PTR1) );
  BUF_X1 U27747 ( .A(_01427__PTR1), .Z(_01445__PTR1) );
  BUF_X1 U27748 ( .A(_01432__PTR1), .Z(_01447__PTR1) );
  BUF_X1 U27749 ( .A(_01427__PTR1), .Z(_01448__PTR1) );
  BUF_X1 U27750 ( .A(_01432__PTR1), .Z(_01450__PTR1) );
  BUF_X1 U27751 ( .A(_01427__PTR1), .Z(_01451__PTR1) );
  BUF_X1 U27752 ( .A(_01432__PTR1), .Z(_01453__PTR1) );
  BUF_X1 U27753 ( .A(_01427__PTR1), .Z(_01454__PTR1) );
  BUF_X1 U27754 ( .A(_01432__PTR1), .Z(_01456__PTR1) );
  BUF_X1 U27755 ( .A(_01427__PTR1), .Z(_01457__PTR1) );
  BUF_X1 U27756 ( .A(_01432__PTR1), .Z(_01459__PTR1) );
  BUF_X1 U27757 ( .A(_01427__PTR1), .Z(_01460__PTR1) );
  BUF_X1 U27758 ( .A(_01432__PTR1), .Z(_01462__PTR1) );
  BUF_X1 U27759 ( .A(_01427__PTR1), .Z(_01463__PTR1) );
  BUF_X1 U27760 ( .A(_01432__PTR1), .Z(_01465__PTR1) );
  BUF_X1 U27761 ( .A(_01427__PTR1), .Z(_01466__PTR1) );
  BUF_X1 U27762 ( .A(_01432__PTR1), .Z(_01468__PTR1) );
  BUF_X1 U27763 ( .A(_01427__PTR1), .Z(_01469__PTR1) );
  BUF_X1 U27764 ( .A(_01432__PTR1), .Z(_01471__PTR1) );
  BUF_X1 U27765 ( .A(_01427__PTR1), .Z(_01472__PTR1) );
  BUF_X1 U27766 ( .A(_01432__PTR1), .Z(_01474__PTR1) );
  BUF_X1 U27767 ( .A(_01427__PTR1), .Z(_01475__PTR1) );
  BUF_X1 U27768 ( .A(_01432__PTR1), .Z(_01477__PTR1) );
  BUF_X1 U27769 ( .A(_01483__PTR1), .Z(_01485__PTR1) );
  BUF_X1 U27770 ( .A(_01424__PTR1), .Z(_01491__PTR1) );
  BUF_X1 U27771 ( .A(_01421__PTR0), .Z(_01492__PTR0) );
  BUF_X1 U27772 ( .A(_01423__PTR1), .Z(_01493__PTR1) );
  BUF_X1 U27773 ( .A(_01352__PTR1), .Z(_01500__PTR1) );
  BUF_X1 U27774 ( .A(_01349__PTR0), .Z(_01501__PTR0) );
  BUF_X1 U27775 ( .A(_01351__PTR1), .Z(_01502__PTR1) );
  BUF_X1 U27776 ( .A(_01507__PTR0), .Z(_01511__PTR0) );
  BUF_X1 U27777 ( .A(_01280__PTR1), .Z(_01522__PTR1) );
  BUF_X1 U27778 ( .A(_01508__PTR0), .Z(_01523__PTR0) );
  BUF_X1 U27779 ( .A(_01507__PTR0), .Z(_01526__PTR0) );
  BUF_X1 U27780 ( .A(_01277__PTR0), .Z(_01527__PTR0) );
  BUF_X1 U27781 ( .A(_01279__PTR1), .Z(_01528__PTR1) );
  BUF_X1 U27782 ( .A(_01511__PTR3), .Z(_01531__PTR3) );
  BUF_X1 U27783 ( .A(_01526__PTR3), .Z(_01538__PTR3) );
  BUF_X1 U27784 ( .A(_01508__PTR0), .Z(_01542__PTR0) );
  BUF_X1 U27785 ( .A(_01548__PTR0), .Z(_01552__PTR0) );
  BUF_X1 U27786 ( .A(_01549__PTR0), .Z(_01557__PTR0) );
  BUF_X1 U27787 ( .A(_01548__PTR0), .Z(_01560__PTR0) );
  BUF_X1 U27788 ( .A(_01552__PTR3), .Z(_01563__PTR3) );
  BUF_X1 U27789 ( .A(_01560__PTR3), .Z(_01567__PTR3) );
  BUF_X1 U27790 ( .A(_01549__PTR0), .Z(_01571__PTR0) );
  BUF_X1 U27791 ( .A(_01577__PTR1), .Z(_01581__PTR1) );
  BUF_X1 U27792 ( .A(_01587__PTR1), .Z(_01589__PTR1) );
  BUF_X1 U27793 ( .A(_01589__PTR0), .Z(_01591__PTR0) );
  BUF_X1 U27794 ( .A(_01589__PTR0), .Z(_01593__PTR0) );
  BUF_X1 U27795 ( .A(_01586__PTR2), .Z(_01594__PTR2) );
  BUF_X1 U27796 ( .A(_01595__PTR1), .Z(_01596__PTR1) );
  BUF_X1 U27797 ( .A(_01600__PTR1), .Z(_01601__PTR1) );
  BUF_X1 U27798 ( .A(_01601__PTR0), .Z(_01603__PTR0) );
  BUF_X1 U27799 ( .A(_01603__PTR1), .Z(_01604__PTR1) );
  BUF_X1 U27800 ( .A(_01598__PTR1), .Z(_01605__PTR1) );
  BUF_X1 U27801 ( .A(_01598__PTR0), .Z(_01606__PTR0) );
  BUF_X1 U27802 ( .A(_01589__PTR0), .Z(_01607__PTR0) );
  BUF_X1 U27803 ( .A(_01544__PTR0), .Z(_01616__PTR0) );
  BUF_X1 U27804 ( .A(_01618__PTR0), .Z(_01622__PTR0) );
  BUF_X1 U27805 ( .A(_01632__PTR1), .Z(_01636__PTR1) );
  BUF_X1 U27806 ( .A(_01642__PTR1), .Z(_01644__PTR1) );
  BUF_X1 U27807 ( .A(_01644__PTR0), .Z(_01646__PTR0) );
  BUF_X1 U27808 ( .A(_01644__PTR0), .Z(_01648__PTR0) );
  BUF_X1 U27809 ( .A(_01641__PTR2), .Z(_01649__PTR2) );
  BUF_X1 U27810 ( .A(_01650__PTR1), .Z(_01651__PTR1) );
  BUF_X1 U27811 ( .A(_01655__PTR1), .Z(_01656__PTR1) );
  BUF_X1 U27812 ( .A(_01656__PTR0), .Z(_01658__PTR0) );
  BUF_X1 U27813 ( .A(_01658__PTR1), .Z(_01659__PTR1) );
  BUF_X1 U27814 ( .A(_01653__PTR1), .Z(_01660__PTR1) );
  BUF_X1 U27815 ( .A(_01653__PTR0), .Z(_01661__PTR0) );
  BUF_X1 U27816 ( .A(_01644__PTR0), .Z(_01662__PTR0) );
  BUF_X1 U27817 ( .A(_01675__PTR1), .Z(_01679__PTR1) );
  BUF_X1 U27818 ( .A(_01617__PTR0), .Z(_01681__PTR0) );
  BUF_X1 U27819 ( .A(_01617__PTR3), .Z(_01684__PTR3) );
  BUF_X1 U27820 ( .A(_01692__PTR1), .Z(_01694__PTR1) );
  BUF_X1 U27821 ( .A(_01694__PTR0), .Z(_01696__PTR0) );
  BUF_X1 U27822 ( .A(_01694__PTR0), .Z(_01698__PTR0) );
  BUF_X1 U27823 ( .A(_01691__PTR2), .Z(_01699__PTR2) );
  BUF_X1 U27824 ( .A(_01700__PTR1), .Z(_01701__PTR1) );
  BUF_X1 U27825 ( .A(_01705__PTR1), .Z(_01706__PTR1) );
  BUF_X1 U27826 ( .A(_01706__PTR0), .Z(_01708__PTR0) );
  BUF_X1 U27827 ( .A(_01708__PTR1), .Z(_01709__PTR1) );
  BUF_X1 U27828 ( .A(_01703__PTR1), .Z(_01710__PTR1) );
  BUF_X1 U27829 ( .A(_01703__PTR0), .Z(_01711__PTR0) );
  BUF_X1 U27830 ( .A(_01694__PTR0), .Z(_01712__PTR0) );
  BUF_X1 U27831 ( .A(_01681__PTR3), .Z(_01725__PTR3) );
  BUF_X1 U27832 ( .A(_01618__PTR0), .Z(_01729__PTR0) );
  BUF_X1 U27833 ( .A(_02123__PTR6), .Z(_01731__PTR0) );
  BUF_X1 U27834 ( .A(_02123__PTR5), .Z(_01732__PTR0) );
  BUF_X1 U27835 ( .A(_02123__PTR4), .Z(_01733__PTR0) );
  BUF_X1 U27836 ( .A(_01577__PTR1), .Z(_01753__PTR1) );
  BUF_X1 U27837 ( .A(_01632__PTR1), .Z(_01758__PTR1) );
  BUF_X1 U27838 ( .A(_01675__PTR1), .Z(_01763__PTR1) );
  BUF_X1 U27839 ( .A(P1_P1_InstQueueWr_Addr_PTR0), .Z(_01838__PTR0) );
  BUF_X1 U27840 ( .A(_01836__PTR0), .Z(_01840__PTR0) );
  BUF_X1 U27841 ( .A(P1_RequestPending), .Z(_01861__PTR3) );
  BUF_X1 U27842 ( .A(_01855__PTR1), .Z(_01863__PTR1) );
  BUF_X1 U27843 ( .A(P1_ReadRequest), .Z(_01865__PTR2) );
  BUF_X1 U27844 ( .A(P1_MemoryFetch), .Z(_01868__PTR2) );
  BUF_X1 U27845 ( .A(_01863__PTR3), .Z(_01870__PTR2) );
  BUF_X1 U27846 ( .A(P1_CodeFetch), .Z(_01872__PTR1) );
  BUF_X1 U27847 ( .A(_01863__PTR3), .Z(_01874__PTR1) );
  BUF_X1 U27848 ( .A(_01897__PTR32), .Z(_01897__PTR31) );
  BUF_X1 U27849 ( .A(P1_P1_PhyAddrPointer_PTR0), .Z(_01996__PTR0) );
  BUF_X1 U27850 ( .A(P1_EBX_PTR0), .Z(_02009__PTR0) );
  BUF_X1 U27851 ( .A(P1_P1_InstAddrPointer_PTR0), .Z(_02019__PTR0) );
  BUF_X1 U27852 ( .A(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02020__PTR0) );
  BUF_X1 U27853 ( .A(_02010__PTR0), .Z(_02026__PTR0) );
  BUF_X1 U27854 ( .A(_02015__PTR0), .Z(_02029__PTR0) );
  BUF_X1 U27855 ( .A(P1_P1_InstAddrPointer_PTR0), .Z(_02037__PTR0) );
  BUF_X1 U27856 ( .A(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02038__PTR0) );
  BUF_X1 U27857 ( .A(_02083__PTR1), .Z(_02083__PTR0) );
  BUF_X1 U27858 ( .A(_01863__PTR2), .Z(_02120__PTR1) );
  BUF_X1 U27859 ( .A(P2_P1_InstQueueWr_Addr_PTR0), .Z(_02131__PTR0) );
  BUF_X1 U27860 ( .A(_02129__PTR0), .Z(_02133__PTR0) );
  BUF_X1 U27861 ( .A(P2_RequestPending), .Z(_02154__PTR3) );
  BUF_X1 U27862 ( .A(_02148__PTR1), .Z(_02156__PTR1) );
  BUF_X1 U27863 ( .A(P2_ReadRequest), .Z(_02158__PTR2) );
  BUF_X1 U27864 ( .A(P2_MemoryFetch), .Z(_02161__PTR2) );
  BUF_X1 U27865 ( .A(_02156__PTR3), .Z(_02163__PTR2) );
  BUF_X1 U27866 ( .A(P2_CodeFetch), .Z(_02165__PTR1) );
  BUF_X1 U27867 ( .A(_02156__PTR3), .Z(_02167__PTR1) );
  BUF_X1 U27868 ( .A(_02189__PTR32), .Z(_02189__PTR31) );
  BUF_X1 U27869 ( .A(P2_P1_PhyAddrPointer_PTR0), .Z(_02288__PTR0) );
  BUF_X1 U27870 ( .A(P2_EBX_PTR0), .Z(_02299__PTR0) );
  BUF_X1 U27871 ( .A(P2_P1_InstAddrPointer_PTR0), .Z(_02309__PTR0) );
  BUF_X1 U27872 ( .A(P2_P1_InstQueueRd_Addr_PTR0), .Z(_02310__PTR0) );
  BUF_X1 U27873 ( .A(_02300__PTR0), .Z(_02316__PTR0) );
  BUF_X1 U27874 ( .A(_02305__PTR0), .Z(_02319__PTR0) );
  BUF_X1 U27875 ( .A(P2_P1_InstAddrPointer_PTR0), .Z(_02327__PTR0) );
  BUF_X1 U27876 ( .A(P2_P1_InstQueueRd_Addr_PTR0), .Z(_02328__PTR0) );
  BUF_X1 U27877 ( .A(_02372__PTR1), .Z(_02372__PTR0) );
  BUF_X1 U27878 ( .A(_02156__PTR2), .Z(_02409__PTR1) );
  BUF_X1 U27879 ( .A(P3_P1_InstQueueWr_Addr_PTR0), .Z(_02420__PTR0) );
  BUF_X1 U27880 ( .A(_02418__PTR0), .Z(_02422__PTR0) );
  BUF_X1 U27881 ( .A(P3_RequestPending), .Z(_02443__PTR3) );
  BUF_X1 U27882 ( .A(_02437__PTR1), .Z(_02445__PTR1) );
  BUF_X1 U27883 ( .A(P3_ReadRequest), .Z(_02447__PTR2) );
  BUF_X1 U27884 ( .A(P3_MemoryFetch), .Z(_02450__PTR2) );
  BUF_X1 U27885 ( .A(_02445__PTR3), .Z(_02452__PTR2) );
  BUF_X1 U27886 ( .A(P3_CodeFetch), .Z(_02454__PTR1) );
  BUF_X1 U27887 ( .A(_02445__PTR3), .Z(_02456__PTR1) );
  BUF_X1 U27888 ( .A(_02478__PTR32), .Z(_02478__PTR31) );
  BUF_X1 U27889 ( .A(P3_P1_PhyAddrPointer_PTR0), .Z(_02577__PTR0) );
  BUF_X1 U27890 ( .A(P3_EBX_PTR0), .Z(_02588__PTR0) );
  BUF_X1 U27891 ( .A(P3_P1_InstAddrPointer_PTR0), .Z(_02598__PTR0) );
  BUF_X1 U27892 ( .A(P3_P1_InstQueueRd_Addr_PTR0), .Z(_02599__PTR0) );
  BUF_X1 U27893 ( .A(_02589__PTR0), .Z(_02605__PTR0) );
  BUF_X1 U27894 ( .A(_02594__PTR0), .Z(_02608__PTR0) );
  BUF_X1 U27895 ( .A(P3_P1_InstAddrPointer_PTR0), .Z(_02616__PTR0) );
  BUF_X1 U27896 ( .A(P3_P1_InstQueueRd_Addr_PTR0), .Z(_02617__PTR0) );
  BUF_X1 U27897 ( .A(_02661__PTR1), .Z(_02661__PTR0) );
  BUF_X1 U27898 ( .A(_02445__PTR2), .Z(_02698__PTR1) );
  BUF_X1 U27899 ( .A(_02718__PTR0), .Z(_02729__PTR0) );
  BUF_X1 U27900 ( .A(_01836__PTR0), .Z(_02735__PTR0) );
  BUF_X1 U27901 ( .A(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02750__PTR0) );
  BUF_X1 U27902 ( .A(P1_P1_InstQueueWr_Addr_PTR0), .Z(_02779__PTR0) );
  BUF_X1 U27903 ( .A(_01836__PTR0), .Z(_02780__PTR0) );
  BUF_X1 U27904 ( .A(_02783__PTR0), .Z(_02784__PTR0) );
  BUF_X1 U27905 ( .A(P1_P1_InstQueueWr_Addr_PTR0), .Z(_02785__PTR0) );
  BUF_X1 U27906 ( .A(_02788__PTR0), .Z(_02789__PTR0) );
  BUF_X1 U27907 ( .A(_01836__PTR0), .Z(_02790__PTR0) );
  BUF_X1 U27908 ( .A(P1_P1_InstQueueWr_Addr_PTR0), .Z(_02791__PTR0) );
  BUF_X1 U27909 ( .A(P1_P1_PhyAddrPointer_PTR2), .Z(_02794__PTR0) );
  BUF_X1 U27910 ( .A(_02795__PTR0), .Z(_02796__PTR0) );
  BUF_X1 U27911 ( .A(P1_P1_PhyAddrPointer_PTR1), .Z(_02797__PTR0) );
  BUF_X1 U27912 ( .A(P1_P1_InstAddrPointer_PTR0), .Z(_02798__PTR0) );
  BUF_X1 U27913 ( .A(P1_P1_InstAddrPointer_PTR1), .Z(_02801__PTR0) );
  BUF_X1 U27914 ( .A(_02803__PTR0), .Z(_02804__PTR0) );
  BUF_X1 U27915 ( .A(_02809__PTR0), .Z(_02810__PTR0) );
  BUF_X1 U27916 ( .A(P1_P1_InstQueueRd_Addr_PTR2), .Z(_02812__PTR0) );
  BUF_X1 U27917 ( .A(P1_P1_InstQueueRd_Addr_PTR0), .Z(_02813__PTR0) );
  BUF_X1 U27918 ( .A(P1_P1_InstQueueRd_Addr_PTR1), .Z(_02817__PTR0) );
  BUF_X1 U27919 ( .A(P1_rEIP_PTR1), .Z(_02821__PTR0) );
  BUF_X1 U27920 ( .A(_01882__PTR7), .Z(_02822__PTR0) );
  BUF_X1 U27921 ( .A(_02825__PTR0), .Z(_02826__PTR0) );
  BUF_X1 U27922 ( .A(P1_EAX_PTR0), .Z(_02827__PTR0) );
  BUF_X1 U27923 ( .A(P1_EBX_PTR0), .Z(_02828__PTR0) );
  BUF_X1 U27924 ( .A(P1_P1_InstAddrPointer_PTR0), .Z(_02829__PTR0) );
  BUF_X1 U27925 ( .A(_02715__PTR0), .Z(_02945__PTR0) );
  BUF_X1 U27926 ( .A(P1_P1_PhyAddrPointer_PTR0), .Z(_02946__PTR0) );
  BUF_X1 U27927 ( .A(_02100__PTR32), .Z(_02947__PTR0) );
  BUF_X1 U27928 ( .A(P1_EBX_PTR0), .Z(_02948__PTR0) );
  BUF_X1 U27929 ( .A(P1_P1_InstAddrPointer_PTR0), .Z(_02949__PTR0) );
  BUF_X1 U27930 ( .A(_02963__PTR0), .Z(_02974__PTR0) );
  BUF_X1 U27931 ( .A(_02129__PTR0), .Z(_02980__PTR0) );
  BUF_X1 U27932 ( .A(P2_P1_InstQueueRd_Addr_PTR0), .Z(_02995__PTR0) );
  BUF_X1 U27933 ( .A(P2_P1_InstQueueWr_Addr_PTR0), .Z(_03024__PTR0) );
  BUF_X1 U27934 ( .A(_02129__PTR0), .Z(_03025__PTR0) );
  BUF_X1 U27935 ( .A(_03028__PTR0), .Z(_03029__PTR0) );
  BUF_X1 U27936 ( .A(P2_P1_InstQueueWr_Addr_PTR0), .Z(_03030__PTR0) );
  BUF_X1 U27937 ( .A(_03033__PTR0), .Z(_03034__PTR0) );
  BUF_X1 U27938 ( .A(_02129__PTR0), .Z(_03035__PTR0) );
  BUF_X1 U27939 ( .A(P2_P1_InstQueueWr_Addr_PTR0), .Z(_03036__PTR0) );
  BUF_X1 U27940 ( .A(P2_P1_PhyAddrPointer_PTR2), .Z(_03039__PTR0) );
  BUF_X1 U27941 ( .A(_03040__PTR0), .Z(_03041__PTR0) );
  BUF_X1 U27942 ( .A(P2_P1_PhyAddrPointer_PTR1), .Z(_03042__PTR0) );
  BUF_X1 U27943 ( .A(P2_P1_InstAddrPointer_PTR0), .Z(_03043__PTR0) );
  BUF_X1 U27944 ( .A(P2_P1_InstAddrPointer_PTR1), .Z(_03046__PTR0) );
  BUF_X1 U27945 ( .A(_03048__PTR0), .Z(_03049__PTR0) );
  BUF_X1 U27946 ( .A(_03054__PTR0), .Z(_03055__PTR0) );
  BUF_X1 U27947 ( .A(P2_P1_InstQueueRd_Addr_PTR2), .Z(_03057__PTR0) );
  BUF_X1 U27948 ( .A(P2_P1_InstQueueRd_Addr_PTR0), .Z(_03058__PTR0) );
  BUF_X1 U27949 ( .A(P2_P1_InstQueueRd_Addr_PTR1), .Z(_03062__PTR0) );
  BUF_X1 U27950 ( .A(P2_rEIP_PTR1), .Z(_03066__PTR0) );
  BUF_X1 U27951 ( .A(_02174__PTR7), .Z(_03067__PTR0) );
  BUF_X1 U27952 ( .A(_03070__PTR0), .Z(_03071__PTR0) );
  BUF_X1 U27953 ( .A(P2_EAX_PTR0), .Z(_03072__PTR0) );
  BUF_X1 U27954 ( .A(P2_EBX_PTR0), .Z(_03073__PTR0) );
  BUF_X1 U27955 ( .A(P2_P1_InstAddrPointer_PTR0), .Z(_03074__PTR0) );
  BUF_X1 U27956 ( .A(_02960__PTR0), .Z(_03190__PTR0) );
  BUF_X1 U27957 ( .A(P2_P1_PhyAddrPointer_PTR0), .Z(_03191__PTR0) );
  BUF_X1 U27958 ( .A(_02389__PTR32), .Z(_03192__PTR0) );
  BUF_X1 U27959 ( .A(P2_EBX_PTR0), .Z(_03193__PTR0) );
  BUF_X1 U27960 ( .A(P2_P1_InstAddrPointer_PTR0), .Z(_03194__PTR0) );
  BUF_X1 U27961 ( .A(_03208__PTR0), .Z(_03219__PTR0) );
  BUF_X1 U27962 ( .A(_02418__PTR0), .Z(_03225__PTR0) );
  BUF_X1 U27963 ( .A(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03240__PTR0) );
  BUF_X1 U27964 ( .A(P3_P1_InstQueueWr_Addr_PTR0), .Z(_03269__PTR0) );
  BUF_X1 U27965 ( .A(_02418__PTR0), .Z(_03270__PTR0) );
  BUF_X1 U27966 ( .A(_03273__PTR0), .Z(_03274__PTR0) );
  BUF_X1 U27967 ( .A(P3_P1_InstQueueWr_Addr_PTR0), .Z(_03275__PTR0) );
  BUF_X1 U27968 ( .A(_03278__PTR0), .Z(_03279__PTR0) );
  BUF_X1 U27969 ( .A(_02418__PTR0), .Z(_03280__PTR0) );
  BUF_X1 U27970 ( .A(P3_P1_InstQueueWr_Addr_PTR0), .Z(_03281__PTR0) );
  BUF_X1 U27971 ( .A(P3_P1_PhyAddrPointer_PTR2), .Z(_03284__PTR0) );
  BUF_X1 U27972 ( .A(_03285__PTR0), .Z(_03286__PTR0) );
  BUF_X1 U27973 ( .A(P3_P1_PhyAddrPointer_PTR1), .Z(_03287__PTR0) );
  BUF_X1 U27974 ( .A(P3_P1_InstAddrPointer_PTR0), .Z(_03288__PTR0) );
  BUF_X1 U27975 ( .A(P3_P1_InstAddrPointer_PTR1), .Z(_03291__PTR0) );
  BUF_X1 U27976 ( .A(_03293__PTR0), .Z(_03294__PTR0) );
  BUF_X1 U27977 ( .A(_03299__PTR0), .Z(_03300__PTR0) );
  BUF_X1 U27978 ( .A(P3_P1_InstQueueRd_Addr_PTR2), .Z(_03302__PTR0) );
  BUF_X1 U27979 ( .A(P3_P1_InstQueueRd_Addr_PTR0), .Z(_03303__PTR0) );
  BUF_X1 U27980 ( .A(P3_P1_InstQueueRd_Addr_PTR1), .Z(_03307__PTR0) );
  BUF_X1 U27981 ( .A(P3_rEIP_PTR1), .Z(_03311__PTR0) );
  BUF_X1 U27982 ( .A(_02463__PTR7), .Z(_03312__PTR0) );
  BUF_X1 U27983 ( .A(_03315__PTR0), .Z(_03316__PTR0) );
  BUF_X1 U27984 ( .A(P3_EAX_PTR0), .Z(_03317__PTR0) );
  BUF_X1 U27985 ( .A(P3_EBX_PTR0), .Z(_03318__PTR0) );
  BUF_X1 U27986 ( .A(P3_P1_InstAddrPointer_PTR0), .Z(_03319__PTR0) );
  BUF_X1 U27987 ( .A(_03205__PTR0), .Z(_03435__PTR0) );
  BUF_X1 U27988 ( .A(P3_P1_PhyAddrPointer_PTR0), .Z(_03436__PTR0) );
  BUF_X1 U27989 ( .A(_02678__PTR32), .Z(_03437__PTR0) );
  BUF_X1 U27990 ( .A(P3_EBX_PTR0), .Z(_03438__PTR0) );
  BUF_X1 U27991 ( .A(P3_P1_InstAddrPointer_PTR0), .Z(_03439__PTR0) );
  BUF_X1 U27992 ( .A(_05712__PTR0), .Z(_05713__PTR0) );
  BUF_X1 U27993 ( .A(_05717__PTR0), .Z(_05718__PTR0) );
  BUF_X1 U27994 ( .A(bs16), .Z(P1_BS16_n) );
  BUF_X1 U27995 ( .A(clock), .Z(P1_CLOCK) );
  BUF_X1 U27996 ( .A(P1_StateBS16), .Z(P1_DataWidth_PTR1) );
  BUF_X1 U27997 ( .A(hold), .Z(P1_HOLD) );
  BUF_X1 U27998 ( .A(na), .Z(P1_NA_n) );
  BUF_X1 U27999 ( .A(reset), .Z(P1_RESET) );
  BUF_X1 U28000 ( .A(bs16), .Z(P2_BS16_n) );
  BUF_X1 U28001 ( .A(clock), .Z(P2_CLOCK) );
  BUF_X1 U28002 ( .A(P2_StateBS16), .Z(P2_DataWidth_PTR1) );
  BUF_X1 U28003 ( .A(hold), .Z(P2_HOLD) );
  BUF_X1 U28004 ( .A(na), .Z(P2_NA_n) );
  BUF_X1 U28005 ( .A(reset), .Z(P2_RESET) );
  BUF_X1 U28006 ( .A(bs16), .Z(P3_BS16_n) );
  BUF_X1 U28007 ( .A(clock), .Z(P3_CLOCK) );
  BUF_X1 U28008 ( .A(P3_StateBS16), .Z(P3_DataWidth_PTR1) );
  BUF_X1 U28009 ( .A(hold), .Z(P3_HOLD) );
  BUF_X1 U28010 ( .A(na), .Z(P3_NA_n) );
  BUF_X1 U28011 ( .A(reset), .Z(P3_RESET) );
  BUF_X1 U28012 ( .A(P1_ADS_n), .Z(ads1) );
  BUF_X1 U28013 ( .A(P2_ADS_n), .Z(ads2) );
  BUF_X1 U28014 ( .A(P3_ADS_n), .Z(ads3) );
  BUF_X1 U28015 ( .A(P1_ADS_n), .Z(ast1) );
  BUF_X1 U28016 ( .A(P3_ADS_n), .Z(ast2) );
  BUF_X1 U28017 ( .A(P3_D_C_n), .Z(dc) );
  BUF_X1 U28018 ( .A(P1_D_C_n), .Z(dc1) );
  BUF_X1 U28019 ( .A(P2_D_C_n), .Z(dc2) );
  BUF_X1 U28020 ( .A(P3_D_C_n), .Z(dc3) );
  BUF_X1 U28021 ( .A(P1_Datai_PTR31), .Z(di1_PTR31) );
  BUF_X1 U28022 ( .A(P2_Datai_PTR31), .Z(di2_PTR31) );
  BUF_X1 U28023 ( .A(P3_M_IO_n), .Z(mio) );
  BUF_X1 U28024 ( .A(P1_M_IO_n), .Z(mio1) );
  BUF_X1 U28025 ( .A(P2_M_IO_n), .Z(mio2) );
  BUF_X1 U28026 ( .A(P3_M_IO_n), .Z(mio3) );
  BUF_X1 U28027 ( .A(P1_READY_n), .Z(rdy1) );
  BUF_X1 U28028 ( .A(P2_READY_n), .Z(rdy2) );
  BUF_X1 U28029 ( .A(P3_READY_n), .Z(rdy3) );
  BUF_X1 U28030 ( .A(P3_W_R_n), .Z(wr) );
  BUF_X1 U28031 ( .A(P1_W_R_n), .Z(wr1) );
  BUF_X1 U28032 ( .A(P2_W_R_n), .Z(wr2) );
  BUF_X1 U28033 ( .A(P3_W_R_n), .Z(wr3) );
  INV_X1 U28034 ( .A(reset), .ZN(reset_n_DEFINE));
endmodule